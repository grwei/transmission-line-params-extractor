* begin ansoft header
* node 1 Diff1
* node 2 Comm1
* node 3 Diff2
* node 4 Comm2
* node 5 Diff3
* node 6 Comm3
* node 7 Diff4
* node 8 Comm4
* node 9 Diff5
* node 10 Comm5
* node 11 Diff6
* node 12 Comm6
* node 13 Diff7
* node 14 Comm7
* node 15 Diff8
* node 16 Comm8
* node 17 Diff9
* node 18 Comm9
* node 19 Diff10
* node 20 Comm10
* node 21 Diff11
* node 22 Comm11
* node 23 Diff12
* node 24 Comm12
* node 25 Diff13
* node 26 Comm13
* node 27 Diff14
* node 28 Comm14
* node 29 Diff15
* node 30 Comm15
* node 31 Diff16
* node 32 Comm16
* 
* created by ElectronicsDesktop
* end ansoft header

.subckt m16lines_HFSS_lfws 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 
rc1_2to1 2 33 1e-05
cs1_2to1 33 1 0.43408179455715p
rp_2to1 2 1 41390.659886936
rc1_2to3 2 34 1e-05
cs1_2to3 34 3 10.664435386465p
rp_2to3 2 3 990.68894188762
rc1_2to4 2 35 1e-05
cs1_2to4 35 4 97.124998694598p
rp_2to4 2 4 75.364565719858
rc1_2to5 2 36 1e-05
cs1_2to5 36 5 452.43317342452p
rp_2to5 2 5 13.485862322185
rc1_2to6 2 37 1e-05
cs1_2to6 37 6 2124.187782732p
rp_2to6 2 6 1.6352715677474
rc1_2to7 2 38 1e-05
cs1_2to7 38 7 3464.2569938979p
rp_2to7 2 7 0.018817616523916
rl1_2to8 2 39 0.0029134010723771
ls1_2to8 39 8 0.003416255975422n
rl1_2to9 2 40 0.0015505610375966
ls1_2to9 40 9 0.0067397400527922n
rc1_2to10 2 41 1e-05
cs1_2to10 41 10 3.4407525557479p
rp_2to10 2 10 3784.8250409959
rc1_2to11 2 42 1e-05
cs1_2to11 42 11 45.390473163145p
rp_2to11 2 11 181.09912618268
rc1_2to12 2 43 1e-05
cs1_2to12 43 12 256.29687646216p
rp_2to12 2 12 24.541666344787
rc1_2to13 2 44 1e-05
cs1_2to13 44 13 1086.5873837108p
rp_2to13 2 13 4.3050098311267
rc1_2to14 2 45 1e-05
cs1_2to14 45 14 2294.6043994303p
rp_2to14 2 14 0.027870601751483
rl1_2to15 2 46 0.0038372206099278
ls1_2to15 46 15 0.00042239001477525n
rl1_2to16 2 47 0.0020257860301404
ls1_2to16 47 16 0.0059306747472775n
rc1_2to17 2 48 1e-05
cs1_2to17 48 17 21779.721499163p
rp_2to17 2 17 0.0019213881768801
rc1_2to18 2 49 1e-05
cs1_2to18 49 18 0.42952508420833p
rp_2to18 2 18 42402.051243127
rc1_2to19 2 50 1e-05
cs1_2to19 50 19 10.381139925389p
rp_2to19 2 19 1040.3209430754
rc1_2to20 2 51 1e-05
cs1_2to20 51 20 91.856461729948p
rp_2to20 2 20 83.505989219319
rc1_2to21 2 52 1e-05
cs1_2to21 52 21 415.67813099365p
rp_2to21 2 21 15.996579916625
rc1_2to22 2 53 1e-05
cs1_2to22 53 22 1804.3830000351p
rp_2to22 2 22 2.3484932306927
rc1_2to23 2 54 1e-05
cs1_2to23 54 23 3459.4895676585p
rp_2to23 2 23 0.018799421041757
rl1_2to24 2 55 0.002894323622245
ls1_2to24 55 24 0.0030224235354907n
rl1_2to25 2 56 0.0015469773533464
ls1_2to25 56 25 0.006582320456149n
rc1_2to26 2 57 1e-05
cs1_2to26 57 26 3.3786469495314p
rp_2to26 2 26 3920.1214457864
rc1_2to27 2 58 1e-05
cs1_2to27 58 27 43.44438642174p
rp_2to27 2 27 196.38065659284
rc1_2to28 2 59 1e-05
cs1_2to28 59 28 238.49706808318p
rp_2to28 2 28 28.073794463092
rc1_2to29 2 60 1e-05
cs1_2to29 60 29 969.2632134196p
rp_2to29 2 29 5.4394858976793
rc1_2to30 2 61 1e-05
cs1_2to30 61 30 8460.9620162697p
rp_2to30 2 30 0.096381725921629
rc1_2to31 2 62 1e-05
cs1_2to31 62 31 6465.3351859619p
rp_2to31 2 31 0.010406958733205
rl1_2to32 2 63 0.0020176151338025
ls1_2to32 63 32 0.0057003390872672n
rc1_3to1 3 64 1e-05
cs1_3to1 64 1 0.40778087971151p
rp_3to1 3 1 42594.380204055
rc1_3to4 3 65 1e-05
cs1_3to4 65 4 9.6828022767863p
rp_3to4 3 4 1052.481928341
rc1_3to5 3 66 1e-05
cs1_3to5 66 5 84.801408962731p
rp_3to5 3 5 83.631652564291
rc1_3to6 3 67 1e-05
cs1_3to6 67 6 391.61877573791p
rp_3to6 3 6 14.766656975539
rc1_3to7 3 68 1e-05
cs1_3to7 68 7 1964.8877295861p
rp_3to7 3 7 1.5383573059525
rc1_3to8 3 69 1e-05
cs1_3to8 69 8 2910.1312264085p
rp_3to8 3 8 0.022922445961842
rl1_3to9 3 70 0.0036210421544318
ls1_3to9 70 9 0.0049966038453599n
rc1_3to10 3 71 1e-05
cs1_3to10 71 10 1.6409308297333p
rp_3to10 3 10 8471.7986324814
rc1_3to11 3 72 1e-05
cs1_3to11 72 11 3.1650325914742p
rp_3to11 3 11 3963.8241725317
rc1_3to12 3 73 1e-05
cs1_3to12 73 12 40.158826940051p
rp_3to12 3 12 198.44560453678
rc1_3to13 3 74 1e-05
cs1_3to13 74 13 221.43749510833p
rp_3to13 3 13 27.897735745969
rc1_3to14 3 75 1e-05
cs1_3to14 75 14 959.98182314133p
rp_3to14 3 14 4.5639230876466
rc1_3to15 3 76 1e-05
cs1_3to15 76 15 1926.8380600001p
rp_3to15 3 15 0.033933518807305
rl1_3to16 3 77 0.0047295911482651
ls1_3to16 77 16 0.0015853897299152n
rl1_3to17 3 78 1.8678864323761
ls1_3to17 78 17 0.38882010173217n
rc1_3to18 3 79 1e-05
cs1_3to18 79 18 10.355078693972p
rp_3to18 3 18 1045.3032465023
rc1_3to19 3 80 1e-05
cs1_3to19 80 19 0.40337336386337p
rp_3to19 3 19 43630.818166172
rc1_3to20 3 81 1e-05
cs1_3to20 81 20 9.4144580418227p
rp_3to20 3 20 1106.8103972871
rc1_3to21 3 82 1e-05
cs1_3to21 82 21 80.058174843223p
rp_3to21 3 21 92.893946752706
rc1_3to22 3 83 1e-05
cs1_3to22 83 22 358.57709243447p
rp_3to22 3 22 17.595333382078
rc1_3to23 3 84 1e-05
cs1_3to23 84 23 1628.3558488915p
rp_3to23 3 23 2.3533000133124
rc1_3to24 3 85 1e-05
cs1_3to24 85 24 2906.0208071473p
rp_3to24 3 24 0.02289811686601
rl1_3to25 3 86 0.0035974726085369
ls1_3to25 86 25 0.0044899571981151n
rc1_3to26 3 87 1e-05
cs1_3to26 87 26 1.6152484895649p
rp_3to26 3 26 8714.2605326182
rc1_3to27 3 88 1e-05
cs1_3to27 88 27 3.1054679970442p
rp_3to27 3 27 4109.2972518166
rc1_3to28 3 89 1e-05
cs1_3to28 89 28 38.377375881225p
rp_3to28 3 28 215.68562948465
rc1_3to29 3 90 1e-05
cs1_3to29 90 29 205.56137715745p
rp_3to29 3 29 32.169120241265
rc1_3to30 3 91 1e-05
cs1_3to30 91 30 848.67789729082p
rp_3to30 3 30 5.8933554726936
rc1_3to31 3 92 1e-05
cs1_3to31 92 31 1924.2437762607p
rp_3to31 3 31 0.033898410077245
rl1_3to32 3 93 0.0046934398412629
ls1_3to32 93 32 0.00086695368304338n
rc1_4to1 4 94 1e-05
cs1_4to1 94 1 0.40737981687342p
rp_4to1 4 1 42620.032527463
rc1_4to5 4 95 1e-05
cs1_4to5 95 5 9.6722271933707p
rp_4to5 4 5 1053.265296082
rc1_4to6 4 96 1e-05
cs1_4to6 96 6 84.684204851442p
rp_4to6 4 6 83.559300685433
rc1_4to7 4 97 1e-05
cs1_4to7 97 7 391.26623583898p
rp_4to7 4 7 14.711842269825
rc1_4to8 4 98 1e-05
cs1_4to8 98 8 1964.1517328659p
rp_4to8 4 8 1.5294683058948
rc1_4to9 4 99 1e-05
cs1_4to9 99 9 2846.2655856939p
rp_4to9 4 9 0.023413754616059
rc1_4to10 4 100 1e-05
cs1_4to10 100 10 25.621622295383p
rp_4to10 4 10 334.91702114436
rc1_4to11 4 101 1e-05
cs1_4to11 101 11 1.6371883684841p
rp_4to11 4 11 8456.6640404641
rc1_4to12 4 102 1e-05
cs1_4to12 102 12 3.163016040155p
rp_4to12 4 12 3965.6731864235
rc1_4to13 4 103 1e-05
cs1_4to13 103 13 40.121901266587p
rp_4to13 4 13 198.28482637616
rc1_4to14 4 104 1e-05
cs1_4to14 104 14 221.10407383716p
rp_4to14 4 14 27.992883756412
rc1_4to15 4 105 1e-05
cs1_4to15 105 15 957.75324733892p
rp_4to15 4 15 4.5599601075123
rc1_4to16 4 106 1e-05
cs1_4to16 106 16 1911.9979753731p
rp_4to16 4 16 0.034237880967906
rl1_4to17 4 107 1.1623473826621
ls1_4to17 107 17 0.057465998179336n
rc1_4to18 4 108 1e-05
cs1_4to18 108 18 91.139607263141p
rp_4to18 4 18 84.742638940046
rc1_4to19 4 109 1e-05
cs1_4to19 109 19 9.41418854785p
rp_4to19 4 19 1106.8682341974
rc1_4to20 4 110 1e-05
cs1_4to20 110 20 0.40297442198914p
rp_4to20 4 20 43657.683556508
rc1_4to21 4 111 1e-05
cs1_4to21 111 21 9.4039247915955p
rp_4to21 4 21 1107.9688049362
rc1_4to22 4 112 1e-05
cs1_4to22 112 22 79.943910783496p
rp_4to22 4 22 92.866503665118
rc1_4to23 4 113 1e-05
cs1_4to23 113 23 358.13293344022p
rp_4to23 4 23 17.553172448538
rc1_4to24 4 114 1e-05
cs1_4to24 114 24 1628.8991613819p
rp_4to24 4 24 2.3374439788267
rc1_4to25 4 115 1e-05
cs1_4to25 115 25 2842.3177180685p
rp_4to25 4 25 0.023392796886955
rc1_4to26 4 116 1e-05
cs1_4to26 116 26 24.622131045002p
rp_4to26 4 26 359.22812535239
rc1_4to27 4 117 1e-05
cs1_4to27 117 27 1.6115081584508p
rp_4to27 4 27 8698.0308911601
rc1_4to28 4 118 1e-05
cs1_4to28 118 28 3.103481511012p
rp_4to28 4 28 4111.3927611256
rc1_4to29 4 119 1e-05
cs1_4to29 119 29 38.339662442765p
rp_4to29 4 29 215.56987261815
rc1_4to30 4 120 1e-05
cs1_4to30 120 30 205.24161203617p
rp_4to30 4 30 32.171054661037
rc1_4to31 4 121 1e-05
cs1_4to31 121 31 846.93249965584p
rp_4to31 4 31 5.8863294589644
rc1_4to32 4 122 1e-05
cs1_4to32 122 32 1909.4329924479p
rp_4to32 4 32 0.034206054997471
rc1_5to1 5 123 1e-05
cs1_5to1 123 1 0.40735319539791p
rp_5to1 5 1 42624.825050511
rc1_5to6 5 124 1e-05
cs1_5to6 124 6 9.6825304567708p
rp_5to6 5 6 1051.9503926414
rc1_5to7 5 125 1e-05
cs1_5to7 125 7 84.689425377131p
rp_5to7 5 7 83.592151086761
rc1_5to8 5 126 1e-05
cs1_5to8 126 8 390.40779123232p
rp_5to8 5 8 14.7825860326
rc1_5to9 5 127 1e-05
cs1_5to9 127 9 1872.4038281212p
rp_5to9 5 9 1.68293670631
rc1_5to10 5 128 1e-05
cs1_5to10 128 10 162.96232555316p
rp_5to10 5 10 39.730137982769
rc1_5to11 5 129 1e-05
cs1_5to11 129 11 25.470527874519p
rp_5to11 5 11 335.34814386765
rc1_5to12 5 130 1e-05
cs1_5to12 130 12 1.6372662005446p
rp_5to12 5 12 8462.3781631081
rc1_5to13 5 131 1e-05
cs1_5to13 131 13 3.1662735699149p
rp_5to13 5 13 3961.3346366609
rc1_5to14 5 132 1e-05
cs1_5to14 132 14 40.104037675354p
rp_5to14 5 14 198.43810171648
rc1_5to15 5 133 1e-05
cs1_5to15 133 15 220.73832664504p
rp_5to15 5 15 27.991994960699
rc1_5to16 5 134 1e-05
cs1_5to16 134 16 948.14038480639p
rp_5to16 5 16 4.6534939239561
rl1_5to17 5 135 -0.0090603570564981
ls1_5to17 135 17 -0.0020936348737897n
rc1_5to18 5 136 1e-05
cs1_5to18 136 18 409.99683102598p
rp_5to18 5 18 16.454091261392
rc1_5to19 5 137 1e-05
cs1_5to19 137 19 80.053218636336p
rp_5to19 5 19 92.899474690701
rc1_5to20 5 138 1e-05
cs1_5to20 138 20 9.4039731229805p
rp_5to20 5 20 1107.9659488605
rc1_5to21 5 139 1e-05
cs1_5to21 139 21 0.40294870518602p
rp_5to21 5 21 43658.200238807
rc1_5to22 5 140 1e-05
cs1_5to22 140 22 9.413929865223p
rp_5to22 5 22 1106.6725988123
rc1_5to23 5 141 1e-05
cs1_5to23 141 23 79.946119424018p
rp_5to23 5 23 92.890172979948
rc1_5to24 5 142 1e-05
cs1_5to24 142 24 357.52196550318p
rp_5to24 5 24 17.639707074703
rc1_5to25 5 143 1e-05
cs1_5to25 143 25 1564.8084720635p
rp_5to25 5 25 2.5168491481335
rc1_5to26 5 144 1e-05
cs1_5to26 144 26 151.99686894282p
rp_5to26 5 26 45.129417868203
rc1_5to27 5 145 1e-05
cs1_5to27 145 27 24.478742346628p
rp_5to27 5 27 359.68412203006
rc1_5to28 5 146 1e-05
cs1_5to28 146 28 1.6115697132391p
rp_5to28 5 28 8704.9823564178
rc1_5to29 5 147 1e-05
cs1_5to29 147 29 3.1066454316985p
rp_5to29 5 29 4107.2966438835
rc1_5to30 5 148 1e-05
cs1_5to30 148 30 38.323362588465p
rp_5to30 5 30 215.64858557301
rc1_5to31 5 149 1e-05
cs1_5to31 149 31 204.94808309294p
rp_5to31 5 31 32.132239016041
rc1_5to32 5 150 1e-05
cs1_5to32 150 32 839.22874176109p
rp_5to32 5 32 5.9879816702615
rc1_6to1 6 151 1e-05
cs1_6to1 151 1 0.40812417666464p
rp_6to1 6 1 42517.141067228
rc1_6to7 6 152 1e-05
cs1_6to7 152 7 9.6713472280431p
rp_6to7 6 7 1052.691316204
rc1_6to8 6 153 1e-05
cs1_6to8 153 8 84.59928018204p
rp_6to8 6 8 83.794173217592
rc1_6to9 6 154 1e-05
cs1_6to9 154 9 381.59759625461p
rp_6to9 6 9 14.680866534261
rc1_6to10 6 155 1e-05
cs1_6to10 155 10 699.11167186741p
rp_6to10 6 10 7.1720461161316
rc1_6to11 6 156 1e-05
cs1_6to11 156 11 161.53511453863p
rp_6to11 6 11 39.834962577992
rc1_6to12 6 157 1e-05
cs1_6to12 157 12 25.489973511655p
rp_6to12 6 12 334.93242042543
rc1_6to13 6 158 1e-05
cs1_6to13 158 13 1.6367999299665p
rp_6to13 6 13 8468.0155121434
rc1_6to14 6 159 1e-05
cs1_6to14 159 14 3.1590346726456p
rp_6to14 6 14 3971.8653067511
rc1_6to15 6 160 1e-05
cs1_6to15 160 15 40.053317047658p
rp_6to15 6 15 198.69245714875
rc1_6to16 6 161 1e-05
cs1_6to16 161 16 219.6621384765p
rp_6to16 6 16 27.815882197113
rc1_6to17 6 162 1e-05
cs1_6to17 162 17 1287090.4924425p
rp_6to17 6 17 100000
rc1_6to18 6 163 1e-05
cs1_6to18 163 18 1747.955098383p
rp_6to18 6 18 2.5254630044835
rc1_6to19 6 164 1e-05
cs1_6to19 164 19 358.35976974562p
rp_6to19 6 19 17.623659451896
rc1_6to20 6 165 1e-05
cs1_6to20 165 20 79.937249122073p
rp_6to20 6 20 92.890884789924
rc1_6to21 6 166 1e-05
cs1_6to21 166 21 9.4137715166221p
rp_6to21 6 21 1106.7717577474
rc1_6to22 6 167 1e-05
cs1_6to22 167 22 0.40370847763494p
rp_6to22 6 22 43550.843643301
rc1_6to23 6 168 1e-05
cs1_6to23 168 23 9.4027537724334p
rp_6to23 6 23 1107.2218046208
rc1_6to24 6 169 1e-05
cs1_6to24 169 24 79.857347467079p
rp_6to24 6 24 93.117445158847
rc1_6to25 6 170 1e-05
cs1_6to25 170 25 349.64177510883p
rp_6to25 6 25 17.399320378025
rc1_6to26 6 171 1e-05
cs1_6to26 171 26 626.7113747648p
rp_6to26 6 26 8.9576097856605
rc1_6to27 6 172 1e-05
cs1_6to27 172 27 150.67257201431p
rp_6to27 6 27 45.264692187646
rc1_6to28 6 173 1e-05
cs1_6to28 173 28 24.495961025259p
rp_6to28 6 28 359.3568574003
rc1_6to29 6 174 1e-05
cs1_6to29 174 29 1.6111235679665p
rp_6to29 6 29 8711.5651449333
rc1_6to30 6 175 1e-05
cs1_6to30 175 30 3.099576000031p
rp_6to30 6 30 4116.393128378
rc1_6to31 6 176 1e-05
cs1_6to31 176 31 38.273801527484p
rp_6to31 6 31 216.01211278475
rc1_6to32 6 177 1e-05
cs1_6to32 177 32 203.89032555113p
rp_6to32 6 32 31.977468879319
rc1_7to1 7 178 1e-05
cs1_7to1 178 1 0.40735020458797p
rp_7to1 7 1 42626.709391353
rc1_7to8 7 179 1e-05
cs1_7to8 179 8 9.6809212577354p
rp_7to8 7 8 1052.0629766652
rc1_7to9 7 180 1e-05
cs1_7to9 180 9 83.259731550702p
rp_7to9 7 9 85.300344659774
rc1_7to10 7 181 1e-05
cs1_7to10 181 10 6011.5575116811p
rp_7to10 7 10 0.11334389345366
rc1_7to11 7 182 1e-05
cs1_7to11 182 11 696.26871455145p
rp_7to11 7 11 7.0974764835869
rc1_7to12 7 183 1e-05
cs1_7to12 183 12 161.53202806141p
rp_7to12 7 12 39.823190173475
rc1_7to13 7 184 1e-05
cs1_7to13 184 13 25.449808185213p
rp_7to13 7 13 335.64664063688
rc1_7to14 7 185 1e-05
cs1_7to14 185 14 1.6396509834084p
rp_7to14 7 14 8441.5253767633
rc1_7to15 7 186 1e-05
cs1_7to15 186 15 3.1604276122535p
rp_7to15 7 15 3970.132934284
rc1_7to16 7 187 1e-05
cs1_7to16 187 16 40.015885540341p
rp_7to16 7 16 198.78634912832
rc1_7to17 7 188 1e-05
cs1_7to17 188 17 3252595.4003063p
rp_7to17 7 17 100000
rc1_7to18 7 189 1e-05
cs1_7to18 189 18 3458.2581519831p
rp_7to18 7 18 0.018853048450245
rc1_7to19 7 190 1e-05
cs1_7to19 190 19 1627.3211778794p
rp_7to19 7 19 2.3587146932138
rc1_7to20 7 191 1e-05
cs1_7to20 191 20 358.13908101186p
rp_7to20 7 20 17.557558430722
rc1_7to21 7 192 1e-05
cs1_7to21 192 21 79.942335738561p
rp_7to21 7 21 92.902541224599
rc1_7to22 7 193 1e-05
cs1_7to22 193 22 9.4028498967086p
rp_7to22 7 22 1107.2032780498
rc1_7to23 7 194 1e-05
cs1_7to23 194 23 0.40294535967671p
rp_7to23 7 23 43660.399763543
rc1_7to24 7 195 1e-05
cs1_7to24 195 24 9.4122201391753p
rp_7to24 7 24 1106.7317562903
rc1_7to25 7 196 1e-05
cs1_7to25 196 25 78.605584552903p
rp_7to25 7 25 94.688469037102
rc1_7to26 7 197 1e-05
cs1_7to26 197 26 4088.5312738207p
rp_7to26 7 26 0.45242017621156
rc1_7to27 7 198 1e-05
cs1_7to27 198 27 624.23045590231p
rp_7to27 7 27 8.8609713336366
rc1_7to28 7 199 1e-05
cs1_7to28 199 28 150.68097607031p
rp_7to28 7 28 45.242613521392
rc1_7to29 7 200 1e-05
cs1_7to29 200 29 24.458078114692p
rp_7to29 7 29 360.03556787729
rc1_7to30 7 201 1e-05
cs1_7to30 201 30 1.6138772662731p
rp_7to30 7 30 8685.3953938528
rc1_7to31 7 202 1e-05
cs1_7to31 202 31 3.1009804734731p
rp_7to31 7 31 4115.4499751324
rc1_7to32 7 203 1e-05
cs1_7to32 203 32 38.235559221215p
rp_7to32 7 32 216.0766188857
rc1_8to1 8 204 1e-05
cs1_8to1 204 1 0.40728437752553p
rp_8to1 8 1 42635.21033486
rc1_8to9 8 205 1e-05
cs1_8to9 205 9 9.5754746697567p
rp_8to9 8 9 1062.2730920591
rc1_8to10 8 206 1e-05
cs1_8to10 206 10 4436.9236046467p
rp_8to10 8 10 0.015383244797449
rc1_8to11 8 207 1e-05
cs1_8to11 207 11 5915.2668968357p
rp_8to11 8 11 0.090361572337287
rc1_8to12 8 208 1e-05
cs1_8to12 208 12 694.23293402233p
rp_8to12 8 12 7.1343818712593
rc1_8to13 8 209 1e-05
cs1_8to13 209 13 161.17330901904p
rp_8to13 8 13 39.972319127337
rc1_8to14 8 210 1e-05
cs1_8to14 210 14 25.50413779011p
rp_8to14 8 14 334.64555316423
rc1_8to15 8 211 1e-05
cs1_8to15 211 15 1.6391999903976p
rp_8to15 8 15 8447.9273554885
rc1_8to16 8 212 1e-05
cs1_8to16 212 16 3.1615973951071p
rp_8to16 8 16 3963.8818442309
rl1_8to17 8 213 -0.0022361131784248
ls1_8to17 213 17 -0.00019038384954982n
rl1_8to18 8 214 0.0028691223377737
ls1_8to18 214 18 0.0028730357906478n
rc1_8to19 8 215 1e-05
cs1_8to19 215 19 2905.938769372p
rp_8to19 8 19 0.023015910628761
rc1_8to20 8 216 1e-05
cs1_8to20 216 20 1628.3717786704p
rp_8to20 8 20 2.3395223026997
rc1_8to21 8 217 1e-05
cs1_8to21 217 21 357.42375004506p
rp_8to21 8 21 17.641691365936
rc1_8to22 8 218 1e-05
cs1_8to22 218 22 79.862846506008p
rp_8to22 8 22 93.098103366292
rc1_8to23 8 219 1e-05
cs1_8to23 219 23 9.4121998745626p
rp_8to23 8 23 1106.7268131209
rc1_8to24 8 220 1e-05
cs1_8to24 220 24 0.40287973615723p
rp_8to24 8 24 43669.382562517
rc1_8to25 8 221 1e-05
cs1_8to25 221 25 9.3087388573641p
rp_8to25 8 25 1116.9711243712
rc1_8to26 8 222 1e-05
cs1_8to26 222 26 4430.3490216608p
rp_8to26 8 26 0.015369362329458
rc1_8to27 8 223 1e-05
cs1_8to27 223 27 4249.8801224687p
rp_8to27 8 27 0.39576869735111
rc1_8to28 8 224 1e-05
cs1_8to28 224 28 622.80536040969p
rp_8to28 8 28 8.8928076244755
rc1_8to29 8 225 1e-05
cs1_8to29 225 29 150.37107364835p
rp_8to29 8 29 45.377902262115
rc1_8to30 8 226 1e-05
cs1_8to30 226 30 24.50904491708p
rp_8to30 8 30 359.07745612187
rc1_8to31 8 227 1e-05
cs1_8to31 227 31 1.6134516492575p
rp_8to31 8 31 8691.2656550616
rc1_8to32 8 228 1e-05
cs1_8to32 228 32 3.1019128758795p
rp_8to32 8 32 4108.8590248666
rc1_9to1 9 229 1e-05
cs1_9to1 229 1 0.40543133453018p
rp_9to1 9 1 42702.205408303
rl1_9to10 9 230 0.0027374117503969
ls1_9to10 230 10 0.0069874981651625n
rc1_9to11 9 231 1e-05
cs1_9to11 231 11 4293.7032389729p
rp_9to11 9 11 0.015921480929876
rc1_9to12 9 232 1e-05
cs1_9to12 232 12 5789.9634772412p
rp_9to12 9 12 0.12511196208849
rc1_9to13 9 233 1e-05
cs1_9to13 233 13 674.58917006878p
rp_9to13 9 13 7.5210186184948
rc1_9to14 9 234 1e-05
cs1_9to14 234 14 158.4669099211p
rp_9to14 9 14 40.954718111196
rc1_9to15 9 235 1e-05
cs1_9to15 235 15 25.161199038468p
rp_9to15 9 15 339.44118726559
rc1_9to16 9 236 1e-05
cs1_9to16 236 16 1.6245357831107p
rp_9to16 9 16 8507.6775631663
rc1_9to17 9 237 1e-05
cs1_9to17 237 17 21035091.901457p
rp_9to17 9 17 100000
rl1_9to18 9 238 0.0015390568218798
ls1_9to18 238 18 0.0064883040950072n
rl1_9to19 9 239 0.0035901415367951
ls1_9to19 239 19 0.0044896813216199n
rc1_9to20 9 240 1e-05
cs1_9to20 240 20 2842.2318333032p
rp_9to20 9 20 0.023501269839189
rc1_9to21 9 241 1e-05
cs1_9to21 241 21 1563.4820452018p
rp_9to21 9 21 2.5228171783861
rc1_9to22 9 242 1e-05
cs1_9to22 242 22 349.77859523215p
rp_9to22 9 22 17.374947451082
rc1_9to23 9 243 1e-05
cs1_9to23 243 23 78.605953043862p
rp_9to23 9 23 94.675543001042
rc1_9to24 9 244 1e-05
cs1_9to24 244 24 9.3087663570312p
rp_9to24 9 24 1116.9861478216
rc1_9to25 9 245 1e-05
cs1_9to25 245 25 0.40102401326546p
rp_9to25 9 25 43735.736996064
rl1_9to26 9 246 0.0027213042067914
ls1_9to26 246 26 0.0066266734528071n
rc1_9to27 9 247 1e-05
cs1_9to27 247 27 4287.39736746p
rp_9to27 9 27 0.015907965474159
rc1_9to28 9 248 1e-05
cs1_9to28 248 28 3944.9903462456p
rp_9to28 9 28 0.47247266330035
rc1_9to29 9 249 1e-05
cs1_9to29 249 29 606.31317157522p
rp_9to29 9 29 9.3999088444888
rc1_9to30 9 250 1e-05
cs1_9to30 250 30 147.87947344773p
rp_9to30 9 30 46.459359301257
rc1_9to31 9 251 1e-05
cs1_9to31 251 31 24.178631487412p
rp_9to31 9 31 363.97255882806
rc1_9to32 9 252 1e-05
cs1_9to32 252 32 1.59892250665p
rp_9to32 9 32 8749.6180853568
rc1_10to1 10 253 1e-05
cs1_10to1 253 1 0.40836221920745p
rp_10to1 10 1 42608.217947673
rc1_10to11 10 254 1e-05
cs1_10to11 254 11 9.7146592543504p
rp_10to11 10 11 1052.7685820302
rc1_10to12 10 255 1e-05
cs1_10to12 255 12 85.394590047521p
rp_10to12 10 12 83.485645266074
rc1_10to13 10 256 1e-05
cs1_10to13 256 13 394.12767639182p
rp_10to13 10 13 14.800829409172
rc1_10to14 10 257 1e-05
cs1_10to14 257 14 1953.4906562728p
rp_10to14 10 14 1.5856770745522
rc1_10to15 10 258 1e-05
cs1_10to15 258 15 2941.4492638335p
rp_10to15 10 15 0.022600588631973
rl1_10to16 10 259 0.0035314574030448
ls1_10to16 259 16 0.0048850474133477n
rl1_10to17 10 260 -0.064608550669489
ls1_10to17 260 17 -0.0039681993913563n
rc1_10to18 10 261 1e-05
cs1_10to18 261 18 3.3749005332901p
rp_10to18 10 18 3929.0587311958
rc1_10to19 10 262 1e-05
cs1_10to19 262 19 1.6152991335403p
rp_10to19 10 19 8713.7629714936
rc1_10to20 10 263 1e-05
cs1_10to20 263 20 24.628505965415p
rp_10to20 10 20 359.06397412619
rc1_10to21 10 264 1e-05
cs1_10to21 264 21 152.0787944166p
rp_10to21 10 21 45.087565558726
rc1_10to22 10 265 1e-05
cs1_10to22 265 22 627.80534691705p
rp_10to22 10 22 8.9205732030245
rc1_10to23 10 266 1e-05
cs1_10to23 266 23 4106.2082607834p
rp_10to23 10 23 0.44589860381214
rc1_10to24 10 267 1e-05
cs1_10to24 267 24 4430.5786716447p
rp_10to24 10 24 0.015342215708446
rl1_10to25 10 268 0.0027115031560485
ls1_10to25 268 25 0.0066258008820171n
rc1_10to26 10 269 1e-05
cs1_10to26 269 26 0.40395514049077p
rp_10to26 10 26 43647.71231187
rc1_10to27 10 270 1e-05
cs1_10to27 270 27 9.446411139505p
rp_10to27 10 27 1107.092725619
rc1_10to28 10 271 1e-05
cs1_10to28 271 28 80.634372955866p
rp_10to28 10 28 92.705172054695
rc1_10to29 10 272 1e-05
cs1_10to29 272 29 361.0189388466p
rp_10to29 10 29 17.607429899369
rc1_10to30 10 273 1e-05
cs1_10to30 273 30 1625.5842957369p
rp_10to30 10 30 2.3998804486491
rc1_10to31 10 274 1e-05
cs1_10to31 274 31 2937.2568673695p
rp_10to31 10 31 0.02257787384228
rl1_10to32 10 275 0.0035107370356884
ls1_10to32 275 32 0.0043750096418616n
rc1_11to1 11 276 1e-05
cs1_11to1 276 1 0.40725800365321p
rp_11to1 11 1 42637.79131721
rc1_11to12 11 277 1e-05
cs1_11to12 277 12 9.6763129366613p
rp_11to12 11 12 1052.8414313637
rc1_11to13 11 278 1e-05
cs1_11to13 278 13 84.702264070127p
rp_11to13 11 13 83.573051339283
rc1_11to14 11 279 1e-05
cs1_11to14 279 14 391.4258292324p
rp_11to14 11 14 14.723982233894
rc1_11to15 11 280 1e-05
cs1_11to15 280 15 1966.77593299p
rp_11to15 11 15 1.5259927469838
rc1_11to16 11 281 1e-05
cs1_11to16 281 16 2887.9947435947p
rp_11to16 11 16 0.02311067727286
rc1_11to17 11 282 1e-05
cs1_11to17 282 17 116223.46392435p
rp_11to17 11 17 100000
rc1_11to18 11 283 1e-05
cs1_11to18 283 18 43.206273252336p
rp_11to18 11 18 198.46984264128
rc1_11to19 11 284 1e-05
cs1_11to19 284 19 3.1054417783124p
rp_11to19 11 19 4109.3619194126
rc1_11to20 11 285 1e-05
cs1_11to20 285 20 1.6115111740797p
rp_11to20 11 20 8698.0177791484
rc1_11to21 11 286 1e-05
cs1_11to21 286 21 24.478976286718p
rp_11to21 11 21 359.67327064976
rc1_11to22 11 287 1e-05
cs1_11to22 287 22 150.71599569741p
rp_11to22 11 22 45.232392123951
rc1_11to23 11 288 1e-05
cs1_11to23 288 23 624.54090919458p
rp_11to23 11 23 8.8460378516815
rc1_11to24 11 289 1e-05
cs1_11to24 289 24 4273.627225798p
rp_11to24 11 24 0.38995861300629
rc1_11to25 11 290 1e-05
cs1_11to25 290 25 4287.701821941p
rp_11to25 11 25 0.015843194423573
rc1_11to26 11 291 1e-05
cs1_11to26 291 26 9.4451784411767p
rp_11to26 11 26 1107.3452759381
rc1_11to27 11 292 1e-05
cs1_11to27 292 27 0.40285472874182p
rp_11to27 11 27 43674.051131622
rc1_11to28 11 293 1e-05
cs1_11to28 293 28 9.4080660961902p
rp_11to28 11 28 1107.3322054029
rc1_11to29 11 294 1e-05
cs1_11to29 294 29 79.963554847588p
rp_11to29 11 29 92.832828653407
rc1_11to30 11 295 1e-05
cs1_11to30 295 30 358.36311585269p
rp_11to30 11 30 17.547060963911
rc1_11to31 11 296 1e-05
cs1_11to31 296 31 1631.5598693468p
rp_11to31 11 31 2.3305521309348
rc1_11to32 11 297 1e-05
cs1_11to32 297 32 2883.9833808305p
rp_11to32 11 32 0.02308926150279
rc1_12to1 12 298 1e-05
cs1_12to1 298 1 0.4076582163172p
rp_12to1 12 1 42573.362176589
rc1_12to13 12 299 1e-05
cs1_12to13 299 13 9.6854911814231p
rp_12to13 12 13 1051.0785035312
rc1_12to14 12 300 1e-05
cs1_12to14 300 14 84.683750249262p
rp_12to14 12 14 83.5721893615
rc1_12to15 12 301 1e-05
cs1_12to15 301 15 390.52185773757p
rp_12to15 12 15 14.794859173487
rc1_12to16 12 302 1e-05
cs1_12to16 302 16 1937.2200316145p
rp_12to16 12 16 1.5757057598282
rl1_12to17 12 303 -0.12667023049375
ls1_12to17 303 17 -0.026189380609664n
rc1_12to18 12 304 1e-05
cs1_12to18 304 18 235.80160946037p
rp_12to18 12 18 28.71031295864
rc1_12to19 12 305 1e-05
cs1_12to19 305 19 38.373877976095p
rp_12to19 12 19 215.7256542323
rc1_12to20 12 306 1e-05
cs1_12to20 306 20 3.1034756225977p
rp_12to20 12 20 4111.470101532
rc1_12to21 12 307 1e-05
cs1_12to21 307 21 1.6115667228164p
rp_12to21 12 21 8705.0807271772
rc1_12to22 12 308 1e-05
cs1_12to22 308 22 24.496269491696p
rp_12to22 12 22 359.33657602445
rc1_12to23 12 309 1e-05
cs1_12to23 309 23 150.66837416716p
rp_12to23 12 23 45.242867271423
rc1_12to24 12 310 1e-05
cs1_12to24 310 24 622.67559504621p
rp_12to24 12 24 8.9019047867794
rc1_12to25 12 311 1e-05
cs1_12to25 311 25 3933.4718491049p
rp_12to25 12 25 0.47602776743452
rc1_12to26 12 312 1e-05
cs1_12to26 312 26 80.592796721066p
rp_12to26 12 26 92.805095083805
rc1_12to27 12 313 1e-05
cs1_12to27 313 27 9.4079255763819p
rp_12to27 12 27 1107.3823052086
rc1_12to28 12 314 1e-05
cs1_12to28 314 28 0.40324892581467p
rp_12to28 12 28 43604.907911916
rc1_12to29 12 315 1e-05
cs1_12to29 315 29 9.4165484862614p
rp_12to29 12 29 1105.6727746903
rc1_12to30 12 316 1e-05
cs1_12to30 316 30 79.935858827336p
rp_12to30 12 30 92.866004673239
rc1_12to31 12 317 1e-05
cs1_12to31 317 31 357.48179430583p
rp_12to31 12 31 17.638253679898
rc1_12to32 12 318 1e-05
cs1_12to32 318 32 1607.1915685992p
rp_12to32 12 32 2.4016513280701
rc1_13to1 13 319 1e-05
cs1_13to1 319 1 0.40758530957895p
rp_13to1 13 1 42591.560605255
rc1_13to14 13 320 1e-05
cs1_13to14 320 14 9.6588726578309p
rp_13to14 13 14 1055.2831694123
rc1_13to15 13 321 1e-05
cs1_13to15 321 15 84.494088373308p
rp_13to15 13 15 83.894550888974
rc1_13to16 13 322 1e-05
cs1_13to16 322 16 387.55514035847p
rp_13to16 13 16 15.139701548754
rl1_13to17 13 323 -0.0050755048644889
ls1_13to17 323 17 -0.00089265417011337n
rc1_13to18 13 324 1e-05
cs1_13to18 324 18 949.78501016526p
rp_13to18 13 18 5.6729966006498
rc1_13to19 13 325 1e-05
cs1_13to19 325 19 205.5260998816p
rp_13to19 13 19 32.174448058787
rc1_13to20 13 326 1e-05
cs1_13to20 326 20 38.339714175903p
rp_13to20 13 20 215.57188397902
rc1_13to21 13 327 1e-05
cs1_13to21 327 21 3.1066399316009p
rp_13to21 13 21 4107.31407054
rc1_13to22 13 328 1e-05
cs1_13to22 328 22 1.6111262665111p
rp_13to22 13 22 8711.4837870262
rc1_13to23 13 329 1e-05
cs1_13to23 329 23 24.458042089919p
rp_13to23 13 23 360.01489554173
rc1_13to24 13 330 1e-05
cs1_13to24 330 24 150.37481185373p
rp_13to24 13 24 45.377374478881
rc1_13to25 13 331 1e-05
cs1_13to25 331 25 606.2857327761p
rp_13to25 13 25 9.4020590029256
rc1_13to26 13 332 1e-05
cs1_13to26 332 26 360.70870597973p
rp_13to26 13 26 17.631673124798
rc1_13to27 13 333 1e-05
cs1_13to27 333 27 79.95793632763p
rp_13to27 13 27 92.839264750399
rc1_13to28 13 334 1e-05
cs1_13to28 334 28 9.4166099448217p
rp_13to28 13 28 1105.6153909576
rc1_13to29 13 335 1e-05
cs1_13to29 335 29 0.40317778715906p
rp_13to29 13 29 43623.688720983
rc1_13to30 13 336 1e-05
cs1_13to30 336 30 9.3911288496808p
rp_13to30 13 30 1109.8085399395
rc1_13to31 13 337 1e-05
cs1_13to31 337 31 79.768401902229p
rp_13to31 13 31 93.183631516479
rc1_13to32 13 338 1e-05
cs1_13to32 338 32 354.90343123786p
rp_13to32 13 32 18.017037588905
rc1_14to1 14 339 1e-05
cs1_14to1 339 1 0.40781143760205p
rp_14to1 14 1 42551.589763148
rc1_14to15 14 340 1e-05
cs1_14to15 340 15 9.6790512647667p
rp_14to15 14 15 1052.1337749148
rc1_14to16 14 341 1e-05
cs1_14to16 341 16 84.4378369414p
rp_14to16 14 16 84.021652235399
rc1_14to17 14 342 1e-05
cs1_14to17 342 17 2299563.5222415p
rp_14to17 14 17 100000
rc1_14to18 14 343 1e-05
cs1_14to18 343 18 7720.5767864198p
rp_14to18 14 18 0.14367964845667
rc1_14to19 14 344 1e-05
cs1_14to19 344 19 848.36771453559p
rp_14to19 14 19 5.8997495277763
rc1_14to20 14 345 1e-05
cs1_14to20 345 20 205.2433033809p
rp_14to20 14 20 32.182078498703
rc1_14to21 14 346 1e-05
cs1_14to21 346 21 38.32250016789p
rp_14to21 14 21 215.67037284636
rc1_14to22 14 347 1e-05
cs1_14to22 347 22 3.099587122184p
rp_14to22 14 22 4116.3665228754
rc1_14to23 14 348 1e-05
cs1_14to23 348 23 1.6138778300794p
rp_14to23 14 23 8685.3757632025
rc1_14to24 14 349 1e-05
cs1_14to24 349 24 24.509210707016p
rp_14to24 14 24 359.08951073074
rc1_14to25 14 350 1e-05
cs1_14to25 350 25 147.87887440095p
rp_14to25 14 25 46.468382407502
rc1_14to26 14 351 1e-05
cs1_14to26 351 26 1622.5519127827p
rp_14to26 14 26 2.4129460935922
rc1_14to27 14 352 1e-05
cs1_14to27 352 27 358.25854774366p
rp_14to27 14 27 17.569758956844
rc1_14to28 14 353 1e-05
cs1_14to28 353 28 79.939549421091p
rp_14to28 14 28 92.873846934543
rc1_14to29 14 354 1e-05
cs1_14to29 354 29 9.3911396953626p
rp_14to29 14 29 1109.8330980551
rc1_14to30 14 355 1e-05
cs1_14to30 355 30 0.40339825880484p
rp_14to30 14 30 43587.515859644
rc1_14to31 14 356 1e-05
cs1_14to31 356 31 9.4103650781846p
rp_14to31 14 31 1106.8640733723
rc1_14to32 14 357 1e-05
cs1_14to32 357 32 79.703533876496p
rp_14to32 14 32 93.373202708674
rc1_15to1 15 358 1e-05
cs1_15to1 358 1 0.40711148558218p
rp_15to1 15 1 42664.123883659
rc1_15to16 15 359 1e-05
cs1_15to16 359 16 9.6735239169251p
rp_15to16 15 16 1051.6940759693
rl1_15to17 15 360 -0.001615127167627
ls1_15to17 360 17 -0.00017454493916822n
rc1_15to18 15 361 1e-05
cs1_15to18 361 18 6463.2229813688p
rp_15to18 15 18 0.010497826075554
rc1_15to19 15 362 1e-05
cs1_15to19 362 19 1924.3484339331p
rp_15to19 15 19 0.033868704979773
rc1_15to20 15 363 1e-05
cs1_15to20 363 20 847.31092612729p
rp_15to20 15 20 5.8780575569734
rc1_15to21 15 364 1e-05
cs1_15to21 364 21 204.94398310286p
rp_15to21 15 21 32.129357720825
rc1_15to22 15 365 1e-05
cs1_15to22 365 22 38.276059563361p
rp_15to22 15 22 215.96246587591
rc1_15to23 15 366 1e-05
cs1_15to23 366 23 3.1009836494058p
rp_15to23 15 23 4115.3748005403
rc1_15to24 15 367 1e-05
cs1_15to24 367 24 1.6134532676084p
rp_15to24 15 24 8691.2162767943
rc1_15to25 15 368 1e-05
cs1_15to25 368 25 24.17888175481p
rp_15to25 15 25 363.94007487624
rc1_15to26 15 369 1e-05
cs1_15to26 369 26 2937.3235611567p
rp_15to26 15 26 0.022674310764423
rc1_15to27 15 370 1e-05
cs1_15to27 370 27 1630.6837206942p
rp_15to27 15 27 2.32992519102
rc1_15to28 15 371 1e-05
cs1_15to28 371 28 357.61248434333p
rp_15to28 15 28 17.622539475932
rc1_15to29 15 372 1e-05
cs1_15to29 372 29 79.77165801941p
rp_15to29 15 29 93.169559421502
rc1_15to30 15 373 1e-05
cs1_15to30 373 30 9.4103920225861p
rp_15to30 15 30 1106.7938032187
rc1_15to31 15 374 1e-05
cs1_15to31 374 31 0.40271109502024p
rp_15to31 15 31 43696.54269428
rc1_15to32 15 375 1e-05
cs1_15to32 375 32 9.4043514606956p
rp_15to32 15 32 1106.3016600741
rc1_16to1 16 376 1e-05
cs1_16to1 376 1 0.40735437317061p
rp_16to1 16 1 42576.897690305
rc1_16to17 16 377 1e-05
cs1_16to17 377 17 16363942.529701p
rp_16to17 16 17 100000
rl1_16to18 16 378 0.0020227811538381
ls1_16to18 378 18 0.0056109353791881n
rl1_16to19 16 379 0.0047021677739806
ls1_16to19 379 19 0.00088851758175202n
rc1_16to20 16 380 1e-05
cs1_16to20 380 20 1909.4922961207p
rp_16to20 16 20 0.034289592891252
rc1_16to21 16 381 1e-05
cs1_16to21 381 21 839.37737445411p
rp_16to21 16 21 5.9830685952541
rc1_16to22 16 382 1e-05
cs1_16to22 382 22 203.96747427031p
rp_16to22 16 22 31.949020118536
rc1_16to23 16 383 1e-05
cs1_16to23 383 23 38.236747963492p
rp_16to23 16 23 216.03517723592
rc1_16to24 16 384 1e-05
cs1_16to24 384 24 3.101924198617p
rp_16to24 16 24 4108.818655811
rc1_16to25 16 385 1e-05
cs1_16to25 385 25 1.5989246300972p
rp_16to25 16 25 8749.5203547477
rl1_16to26 16 386 0.0035190051940038
ls1_16to26 386 26 0.0043962810976615n
rc1_16to27 16 387 1e-05
cs1_16to27 387 27 2883.9493557808p
rp_16to27 16 27 0.02317076022628
rc1_16to28 16 388 1e-05
cs1_16to28 388 28 1610.8251504658p
rp_16to28 16 28 2.3857230372652
rc1_16to29 16 389 1e-05
cs1_16to29 389 29 355.00346148003p
rp_16to29 16 29 18.010377304048
rc1_16to30 16 390 1e-05
cs1_16to30 390 30 79.708433913528p
rp_16to30 16 30 93.343286895877
rc1_16to31 16 391 1e-05
cs1_16to31 391 31 9.4043857866133p
rp_16to31 16 31 1106.3383913506
rc1_16to32 16 392 1e-05
cs1_16to32 392 32 0.40293959897948p
rp_16to32 16 32 43611.937609344
rl1_17to1 17 393 3877.4008078524
ls1_17to1 393 1 238.69691606866n
rs2_17to1 17 394 0.045497522217195
ls2_17to1 394 1 2.1214599800265n
rl1_17to18 17 395 0.01091658679262
ls1_17to18 395 18 0.64624315446553n
rl1_17to19 17 396 0.0005507001953059
ls1_17to19 396 19 0.080754994625889n
rl1_17to20 17 397 24.225751110154
ls1_17to20 397 20 5.3695069507164n
rs2_17to20 17 398 0.00023788066164449
ls2_17to20 398 20 0.020995754291586n
rl1_17to21 17 399 0.00032600178632035
ls1_17to21 399 21 0.0072483470791022n
rl1_17to22 17 400 0.00013841660074146
ls1_17to22 400 22 0.0028052963685809n
rl1_17to23 17 401 7.6135052843624e-05
ls1_17to23 401 23 0.0011491701892959n
rl1_17to24 17 402 4.9638671866278e-05
ls1_17to24 402 24 0.00046739954514983n
rl1_17to25 17 403 2.4071607765927e-05
ls1_17to25 403 25 0.00017744341498623n
rl1_17to26 17 404 0.0017614358641308
ls1_17to26 404 26 0.16203980599713n
rl1_17to27 17 405 1959.7673778891
ls1_17to27 405 27 174.20865917343n
rs2_17to27 17 406 0.00036453121475418
ls2_17to27 406 27 0.033630075135049n
rl1_17to28 17 407 0.00029271028140215
ls1_17to28 407 28 0.010683290726585n
rl1_17to29 17 408 0.00021635970065319
ls1_17to29 408 29 0.0040544482675638n
rl1_17to30 17 409 9.7302866976085e-05
ls1_17to30 409 30 0.0016354519762951n
rl1_17to31 17 410 7.1501898038073e-05
ls1_17to31 410 31 0.00068847095515629n
rl1_17to32 17 411 4.2692676949942e-05
ls1_17to32 411 32 0.00027629091776461n
rc1_18to1 18 412 1e-05
cs1_18to1 412 1 0.43502714728595p
rp_18to1 18 1 41246.693390004
rc1_18to19 18 413 1e-05
cs1_18to19 413 19 10.733002264686p
rp_18to19 18 19 980.3864334489
rc1_18to20 18 414 1e-05
cs1_18to20 414 20 98.716135861426p
rp_18to20 18 20 73.132165378393
rc1_18to21 18 415 1e-05
cs1_18to21 415 21 467.013775116p
rp_18to21 18 21 12.573667309455
rc1_18to22 18 416 1e-05
cs1_18to22 416 22 2304.1387511576p
rp_18to22 18 22 1.3345306724197
rc1_18to23 18 417 1e-05
cs1_18to23 417 23 3467.5163806732p
rp_18to23 18 23 0.018831929654522
rl1_18to24 18 418 0.0029773787573099
ls1_18to24 418 24 0.0037236742163561n
rl1_18to25 18 419 0.0015939365311556
ls1_18to25 419 25 0.0069049271049764n
rc1_18to26 18 420 1e-05
cs1_18to26 420 26 3.4551343973896p
rp_18to26 18 26 3759.7043221012
rc1_18to27 18 421 1e-05
cs1_18to27 421 27 45.924994747989p
rp_18to27 18 27 177.29326593291
rc1_18to28 18 422 1e-05
cs1_18to28 422 28 262.5555472089p
rp_18to28 18 28 23.398175331679
rc1_18to29 18 423 1e-05
cs1_18to29 423 29 1142.6954417932p
rp_18to29 18 29 3.8271561947727
rc1_18to30 18 424 1e-05
cs1_18to30 424 30 2296.4216487116p
rp_18to30 18 30 0.027887190426542
rl1_18to31 18 425 0.0039170080647683
ls1_18to31 425 31 0.00083698995205366n
rl1_18to32 18 426 0.0020864190216311
ls1_18to32 426 32 0.0061488476932654n
rc1_19to1 19 427 1e-05
cs1_19to1 427 1 0.40779697082642p
rp_19to1 19 1 42591.313342486
rc1_19to20 19 428 1e-05
cs1_19to20 428 20 9.6865567054527p
rp_19to20 19 20 1051.3102584357
rc1_19to21 19 429 1e-05
cs1_19to21 429 21 85.007575295755p
rp_19to21 19 21 83.057493045031
rc1_19to22 19 430 1e-05
cs1_19to22 430 22 394.77860306033p
rp_19to22 19 22 14.438134622264
rc1_19to23 19 431 1e-05
cs1_19to23 431 23 2033.5148872956p
rp_19to23 19 23 1.3942910166114
rc1_19to24 19 432 1e-05
cs1_19to24 432 24 2911.6097829018p
rp_19to24 19 24 0.022933050285289
rl1_19to25 19 433 0.0036846326148087
ls1_19to25 433 25 0.0052387992478942n
rc1_19to26 19 434 1e-05
cs1_19to26 434 26 1.6413265629722p
rp_19to26 19 26 8467.6068003722
rc1_19to27 19 435 1e-05
cs1_19to27 435 27 3.1655258565379p
rp_19to27 19 27 3962.8523771462
rc1_19to28 19 436 1e-05
cs1_19to28 436 28 40.209549806847p
rp_19to28 19 28 197.73350149134
rc1_19to29 19 437 1e-05
cs1_19to29 437 29 222.57867235545p
rp_19to29 19 29 27.57029778911
rc1_19to30 19 438 1e-05
cs1_19to30 438 30 977.05676422861p
rp_19to30 19 30 4.3460275854328
rc1_19to31 19 439 1e-05
cs1_19to31 439 31 1927.6244241457p
rp_19to31 19 31 0.033947160497986
rl1_19to32 19 440 0.0048086986790943
ls1_19to32 440 32 0.0018778281473456n
rc1_20to1 20 441 1e-05
cs1_20to1 441 1 0.40738711038703p
rp_20to1 20 1 42619.048374495
rc1_20to21 20 442 1e-05
cs1_20to21 442 21 9.6750168426386p
rp_20to21 20 21 1052.2173765043
rc1_20to22 20 443 1e-05
cs1_20to22 443 22 84.862244371151p
rp_20to22 20 22 83.074628312966
rc1_20to23 20 444 1e-05
cs1_20to23 444 23 394.40140358155p
rp_20to23 20 23 14.397899386426
rc1_20to24 20 445 1e-05
cs1_20to24 445 24 2039.7049162987p
rp_20to24 20 24 1.3742421921072
rc1_20to25 20 446 1e-05
cs1_20to25 446 25 2847.7697635202p
rp_20to25 20 25 0.023424027579948
rc1_20to26 20 447 1e-05
cs1_20to26 447 26 25.657339130017p
rp_20to26 20 26 333.82303359587
rc1_20to27 20 448 1e-05
cs1_20to27 448 27 1.6372760853802p
rp_20to27 20 27 8454.699773072
rc1_20to28 20 449 1e-05
cs1_20to28 449 28 3.163332313405p
rp_20to28 20 28 3964.6212297497
rc1_20to29 20 450 1e-05
cs1_20to29 450 29 40.165953285014p
rp_20to29 20 29 197.60291390737
rc1_20to30 20 451 1e-05
cs1_20to30 451 30 222.22949988895p
rp_20to30 20 30 27.472819166735
rc1_20to31 20 452 1e-05
cs1_20to31 452 31 976.14493928319p
rp_20to31 20 31 4.3239997201953
rc1_20to32 20 453 1e-05
cs1_20to32 453 32 1912.7860449618p
rp_20to32 20 32 0.034251810150047
rc1_21to1 21 454 1e-05
cs1_21to1 454 1 0.40735997264775p
rp_21to1 21 1 42622.246476837
rc1_21to22 21 455 1e-05
cs1_21to22 455 22 9.6852010772747p
rp_21to22 21 22 1051.060596596
rc1_21to23 21 456 1e-05
cs1_21to23 456 23 84.868722593171p
rp_21to23 21 23 83.082329864828
rc1_21to24 21 457 1e-05
cs1_21to24 457 24 393.67183067197p
rp_21to24 21 24 14.474175168433
rc1_21to25 21 458 1e-05
cs1_21to25 458 25 1942.5832310992p
rp_21to25 21 25 1.5155773087741
rc1_21to26 21 459 1e-05
cs1_21to26 459 26 163.81518864697p
rp_21to26 21 26 39.208385003886
rc1_21to27 21 460 1e-05
cs1_21to27 460 27 25.48942006961p
rp_21to27 21 27 334.56786782632
rc1_21to28 21 461 1e-05
cs1_21to28 461 28 1.6373406232182p
rp_21to28 21 28 8460.8080470689
rc1_21to29 21 462 1e-05
cs1_21to29 462 29 3.166589037934p
rp_21to29 21 29 3961.1401238675
rc1_21to30 21 463 1e-05
cs1_21to30 463 30 40.147455355102p
rp_21to30 21 30 197.67869876793
rc1_21to31 21 464 1e-05
cs1_21to31 464 31 221.90480051454p
rp_21to31 21 31 27.437988637809
rc1_21to32 21 465 1e-05
cs1_21to32 465 32 966.04354155071p
rp_21to32 21 32 4.4100394926603
rc1_22to1 22 466 1e-05
cs1_22to1 466 1 0.40813177804738p
rp_22to1 22 1 42515.767123682
rc1_22to23 22 467 1e-05
cs1_22to23 467 23 9.6738526874499p
rp_22to23 22 23 1051.7233734281
rc1_22to24 22 468 1e-05
cs1_22to24 468 24 84.775465640067p
rp_22to24 22 24 83.285463793166
rc1_22to25 22 469 1e-05
cs1_22to25 469 25 384.6729703856p
rp_22to25 22 25 14.442567567966
rc1_22to26 22 470 1e-05
cs1_22to26 470 26 709.39267355289p
rp_22to26 22 26 6.8951897517596
rc1_22to27 22 471 1e-05
cs1_22to27 471 27 162.13846701101p
rp_22to27 22 27 39.415818525898
rc1_22to28 22 472 1e-05
cs1_22to28 472 28 25.506861650278p
rp_22to28 22 28 334.2438504843
rc1_22to29 22 473 1e-05
cs1_22to29 473 29 1.6368743363645p
rp_22to29 22 29 8466.7395121274
rc1_22to30 22 474 1e-05
cs1_22to30 474 30 3.1593211838317p
rp_22to30 22 30 3970.0818680689
rc1_22to31 22 475 1e-05
cs1_22to31 475 31 40.096126480652p
rp_22to31 22 31 198.09873194829
rc1_22to32 22 476 1e-05
cs1_22to32 476 32 220.73948927831p
rp_22to32 22 32 27.449448094158
rc1_23to1 23 477 1e-05
cs1_23to1 477 1 0.40735686975929p
rp_23to1 23 1 42624.802530499
rc1_23to24 23 478 1e-05
cs1_23to24 478 24 9.6836128645392p
rp_23to24 23 24 1051.0609400593
rc1_23to25 23 479 1e-05
cs1_23to25 479 25 83.437270293159p
rp_23to25 23 25 84.768817185629
rc1_23to26 23 480 1e-05
cs1_23to26 480 26 5735.0819755638p
rp_23to26 23 26 0.079093991646932
rc1_23to27 23 481 1e-05
cs1_23to27 481 27 705.50590400895p
rp_23to27 23 27 6.8352436032481
rc1_23to28 23 482 1e-05
cs1_23to28 482 28 162.11268512461p
rp_23to28 23 28 39.413121446739
rc1_23to29 23 483 1e-05
cs1_23to29 483 29 25.466840623531p
rp_23to29 23 29 334.90943251362
rc1_23to30 23 484 1e-05
cs1_23to30 484 30 1.6397283080709p
rp_23to30 23 30 8440.0838759818
rc1_23to31 23 485 1e-05
cs1_23to31 485 31 3.160727104739p
rp_23to31 23 31 3969.2108926329
rc1_23to32 23 486 1e-05
cs1_23to32 486 32 40.059386548494p
rp_23to32 23 32 198.06236622649
rc1_24to1 24 487 1e-05
cs1_24to1 487 1 0.40729104688662p
rp_24to1 24 1 42633.259469884
rc1_24to25 24 488 1e-05
cs1_24to25 488 25 9.5782195442973p
rp_24to25 24 25 1061.2229551489
rc1_24to26 24 489 1e-05
cs1_24to26 489 26 4439.9681166968p
rp_24to26 24 26 0.015393290698778
rc1_24to27 24 490 1e-05
cs1_24to27 490 27 1545.3890259821p
rp_24to27 24 27 0.042263819003194
rc1_24to28 24 491 1e-05
cs1_24to28 491 28 703.4443171284p
rp_24to28 24 28 6.8764229676901
rc1_24to29 24 492 1e-05
cs1_24to29 492 29 161.78497681038p
rp_24to29 24 29 39.526888946405
rc1_24to30 24 493 1e-05
cs1_24to30 493 30 25.522101873373p
rp_24to30 24 30 333.92385048049
rc1_24to31 24 494 1e-05
cs1_24to31 494 31 1.6392857445533p
rp_24to31 24 31 8446.2044888207
rc1_24to32 24 495 1e-05
cs1_24to32 495 32 3.1619124126523p
rp_24to32 24 32 3962.0851698771
rc1_25to1 25 496 1e-05
cs1_25to1 496 1 0.40543835822388p
rp_25to1 25 1 42700.336366257
rl1_25to26 25 497 0.0027929181020933
ls1_25to26 497 26 0.0071850025527n
rc1_25to27 25 498 1e-05
cs1_25to27 498 27 4296.6604360358p
rp_25to27 25 27 0.015930639811838
rc1_25to28 25 499 1e-05
cs1_25to28 499 28 5658.0538132149p
rp_25to28 25 28 0.086432274832281
rc1_25to29 25 500 1e-05
cs1_25to29 500 29 683.45944783702p
rp_25to29 25 29 7.3239965429597
rc1_25to30 25 501 1e-05
cs1_25to30 501 30 159.07213009293p
rp_25to30 25 30 40.511173695573
rc1_25to31 25 502 1e-05
cs1_25to31 502 31 25.17976632776p
rp_25to31 25 31 338.64184227904
rc1_25to32 25 503 1e-05
cs1_25to32 503 32 1.6246160344991p
rp_25to32 25 32 8505.6868945903
rc1_26to1 26 504 1e-05
cs1_26to1 504 1 0.40841192589195p
rp_26to1 26 1 42600.887196369
rc1_26to27 26 505 1e-05
cs1_26to27 505 27 9.7216068210888p
rp_26to27 26 27 1051.0922358759
rc1_26to28 26 506 1e-05
cs1_26to28 506 28 85.668668918212p
rp_26to28 26 28 82.816083003251
rc1_26to29 26 507 1e-05
cs1_26to29 507 29 397.98321910081p
rp_26to29 26 29 14.389089274563
rc1_26to30 26 508 1e-05
cs1_26to30 508 30 2028.1192031926p
rp_26to30 26 30 1.4282796950693
rc1_26to31 26 509 1e-05
cs1_26to31 509 31 2943.0885600124p
rp_26to31 26 31 0.022612937597407
rl1_26to32 26 510 0.0036036936706991
ls1_26to32 510 32 0.0051291035036634n
rc1_27to1 27 511 1e-05
cs1_27to1 511 1 0.40726567416878p
rp_27to1 27 1 42635.301386126
rc1_27to28 27 512 1e-05
cs1_27to28 512 28 9.6791674801902p
rp_27to28 27 28 1051.8128567367
rc1_27to29 27 513 1e-05
cs1_27to29 513 29 84.88739797213p
rp_27to29 27 29 83.024087947094
rc1_27to30 27 514 1e-05
cs1_27to30 514 30 394.6280303724p
rp_27to30 27 30 14.393374901583
rc1_27to31 27 515 1e-05
cs1_27to31 515 31 2044.6781365878p
rp_27to31 27 31 1.3647694945073
rc1_27to32 27 516 1e-05
cs1_27to32 516 32 2889.5727444515p
rp_27to32 27 32 0.023123603934605
rc1_28to1 28 517 1e-05
cs1_28to1 517 1 0.40766513179276p
rp_28to1 28 1 42571.77048133
rc1_28to29 28 518 1e-05
cs1_28to29 518 29 9.6881334772063p
rp_28to29 28 29 1050.1024320635
rc1_28to30 28 519 1e-05
cs1_28to30 519 30 84.858509881753p
rp_28to30 28 30 83.082975154106
rc1_28to31 28 520 1e-05
cs1_28to31 520 31 393.73813181256p
rp_28to31 28 31 14.446482202281
rc1_28to32 28 521 1e-05
cs1_28to32 521 32 2008.1684704474p
rp_28to32 28 32 1.4189991465209
rc1_29to1 29 522 1e-05
cs1_29to1 522 1 0.40759262208907p
rp_29to1 29 1 42589.314575103
rc1_29to30 29 523 1e-05
cs1_29to30 523 30 9.6614556814286p
rp_29to30 29 30 1054.2758925151
rc1_29to31 29 524 1e-05
cs1_29to31 524 31 84.67770328488p
rp_29to31 29 31 83.344748493082
rc1_29to32 29 525 1e-05
cs1_29to32 525 32 390.75980907997p
rp_29to32 29 32 14.720830094001
rc1_30to1 30 526 1e-05
cs1_30to1 526 1 0.40781870145709p
rp_30to1 30 1 42549.517057362
rc1_30to31 30 527 1e-05
cs1_30to31 527 31 9.6817740323717p
rp_30to31 30 31 1051.1393254118
rc1_30to32 30 528 1e-05
cs1_30to32 528 32 84.622077770275p
rp_30to32 30 32 83.474864644289
rc1_31to1 31 529 1e-05
cs1_31to1 529 1 0.40711773392063p
rp_31to1 31 1 42661.36608065
rc1_31to32 31 530 1e-05
cs1_31to32 530 32 9.6763931273005p
rp_31to32 31 32 1050.6017977891
rc1_32to1 32 531 1e-05
cs1_32to1 531 1 0.40736135216154p
rp_32to1 32 1 42574.843218934
rc1_1to0 1 532 1e-05
cs1_1to0 532 0 0.1587076898489p
rp_1to0 1 0 102252.42191635
rc1_2to0 2 533 1e-05
cs1_2to0 533 0 0.13737444693441p
rp_2to0 2 0 111297.1512637
rc1_3to0 3 534 1e-05
cs1_3to0 534 0 0.13526971508984p
rp_3to0 3 0 113090.34553058
rc1_4to0 4 535 1e-05
cs1_4to0 535 0 0.13489931077123p
rp_4to0 4 0 110207.58012295
rc1_5to0 5 536 1e-05
cs1_5to0 536 0 0.13474917091716p
rp_5to0 5 0 108843.90599685
rc1_6to0 6 537 1e-05
cs1_6to0 537 0 0.13506522380771p
rp_6to0 6 0 113741.47487156
rc1_7to0 7 538 1e-05
cs1_7to0 538 0 0.13493199386525p
rp_7to0 7 0 114124.51297854
rc1_8to0 8 539 1e-05
cs1_8to0 539 0 0.13577710323177p
rp_8to0 8 0 113195.02088027
rc1_9to0 9 540 1e-05
cs1_9to0 540 0 0.15856962580861p
rp_9to0 9 0 103268.03707777
rc1_10to0 10 541 1e-05
cs1_10to0 541 0 0.13579518564933p
rp_10to0 10 0 110333.63209519
rc1_11to0 11 542 1e-05
cs1_11to0 542 0 0.13486711847735p
rp_11to0 11 0 111071.88913359
rc1_12to0 12 543 1e-05
cs1_12to0 543 0 0.13492777716963p
rp_12to0 12 0 115256.91826147
rc1_13to0 13 544 1e-05
cs1_13to0 544 0 0.13477083114449p
rp_13to0 13 0 114446.97661831
rc1_14to0 14 545 1e-05
cs1_14to0 545 0 0.1350451295156p
rp_14to0 14 0 107574.71996649
rc1_15to0 15 546 1e-05
cs1_15to0 546 0 0.1351419884185p
rp_15to0 15 0 109182.54737611
rc1_16to0 16 547 1e-05
cs1_16to0 547 0 0.13746681152166p
rp_16to0 16 0 109454.60409097
rc1_17to0 17 548 1e-05
cs1_17to0 548 0 0.15771872579925p
rp_17to0 17 0 102819.35585508
rc1_18to0 18 549 1e-05
cs1_18to0 549 0 0.13662660693869p
rp_18to0 18 0 114205.71863582
rc1_19to0 19 550 1e-05
cs1_19to0 550 0 0.13441916968016p
rp_19to0 19 0 112584.06676425
rc1_20to0 20 551 1e-05
cs1_20to0 551 0 0.1338569359882p
rp_20to0 20 0 115658.9828005
rc1_21to0 21 552 1e-05
cs1_21to0 552 0 0.13378496843226p
rp_21to0 21 0 117343.48430682
rc1_22to0 22 553 1e-05
cs1_22to0 553 0 0.1339611381753p
rp_22to0 22 0 111577.89504655
rc1_23to0 23 554 1e-05
cs1_23to0 554 0 0.1340699183362p
rp_23to0 23 0 111714.22377891
rc1_24to0 24 555 1e-05
cs1_24to0 555 0 0.13487801038486p
rp_24to0 24 0 112677.93952924
rc1_25to0 25 556 1e-05
cs1_25to0 556 0 0.15759976408982p
rp_25to0 25 0 102036.99423683
rc1_26to0 26 557 1e-05
cs1_26to0 557 0 0.13488310192435p
rp_26to0 26 0 115549.79170562
rc1_27to0 27 558 1e-05
cs1_27to0 558 0 0.13403181129014p
rp_27to0 27 0 114832.51978209
rc1_28to0 28 559 1e-05
cs1_28to0 559 0 0.13391777346909p
rp_28to0 28 0 110311.62432555
rc1_29to0 29 560 1e-05
cs1_29to0 560 0 0.13384371421577p
rp_29to0 29 0 111359.38024123
rc1_30to0 30 561 1e-05
cs1_30to0 561 0 0.13402245450904p
rp_30to0 30 0 118314.40177251
rc1_31to0 31 562 1e-05
cs1_31to0 562 0 0.13426908900929p
rp_31to0 31 0 117094.05413846
rc1_32to0 32 563 1e-05
cs1_32to0 563 0 0.13670763052309p
rp_32to0 32 0 115898.03735148
.ends m16lines_HFSS_lfws

