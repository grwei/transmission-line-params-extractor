* BEGIN ANSOFT HEADER
* node 1    trace_p_0_T1
* node 2    trace_n_0_T1
* node 3    trace_p_1_T1
* node 4    trace_n_1_T1
* node 5    trace_p_0_T2
* node 6    trace_n_0_T2
* node 7    trace_p_1_T2
* node 8    trace_n_1_T2
*   Format: HSPICE
*   Topckt: m4linesveryHighFreq_HFSS_100mil_fws
*     Date: Sat Jun 06 18:38:45 2020
*    Notes: Frequency range: 1e+08 to 2.996e+11 Hz, 600 points
*         : Maximum number of poles: 10000
*         : S-Matrix fitting error tolerance: 0.001
*         : Causality check tolerance: auto
*         : Passivity enforcement: on (by iterated fitting)
*         : Causality enforcement: off
*         : Fitting method: FastFit
*         : Matrix fitting: By entire matrix (required by FastFit)
*         : Ensure Z-parameter accuracy: on
*         : Relative error control: off
*         : Common ground option: on
*         : Final fitting error: 0.259208
*         : Final model order: 448
* END ANSOFT HEADER

.subckt m4linesveryHighFreq_HFSS_100mil_fws 1 2 3 4 5 6 7 8
Vam1 1 n2 dc 0
Rport1 n2 0 50 noise=0
Vam2 2 n4 dc 0
Rport2 n4 0 50 noise=0
Vam3 3 n6 dc 0
Rport3 n6 0 50 noise=0
Vam4 4 n8 dc 0
Rport4 n8 0 50 noise=0
Vam5 5 n10 dc 0
Rport5 n10 0 50 noise=0
Vam6 6 n12 dc 0
Rport6 n12 0 50 noise=0
Vam7 7 n14 dc 0
Rport7 n14 0 50 noise=0
Vam8 8 n16 dc 0
Rport8 n16 0 50 noise=0

Fi1 0 ni1 Vam1 50
Gi1 0 ni1 1 0 1
Rt1 ni1 0 1 noise=0
Fi2 0 ni2 Vam2 50
Gi2 0 ni2 2 0 1
Rt2 ni2 0 1 noise=0
Fi3 0 ni3 Vam3 50
Gi3 0 ni3 3 0 1
Rt3 ni3 0 1 noise=0
Fi4 0 ni4 Vam4 50
Gi4 0 ni4 4 0 1
Rt4 ni4 0 1 noise=0
Fi5 0 ni5 Vam5 50
Gi5 0 ni5 5 0 1
Rt5 ni5 0 1 noise=0
Fi6 0 ni6 Vam6 50
Gi6 0 ni6 6 0 1
Rt6 ni6 0 1 noise=0
Fi7 0 ni7 Vam7 50
Gi7 0 ni7 7 0 1
Rt7 ni7 0 1 noise=0
Fi8 0 ni8 Vam8 50
Gi8 0 ni8 8 0 1
Rt8 ni8 0 1 noise=0

Ca1 ns1 0 1e-12
Ca2 ns2 0 1e-12
Ra1 ns1 0 0.177524466588 noise=0
Ra2 ns2 0 0.177524466588 noise=0
Ga1 ns1 0 ns2 0 -0.592192182122
Ga2 ns2 0 ns1 0 0.592192182122
Ca3 ns3 0 1e-12
Ca4 ns4 0 1e-12
Ra3 ns3 0 3.73043526058 noise=0
Ra4 ns4 0 3.73043526058 noise=0
Ga3 ns3 0 ns4 0 -1.88816876812
Ga4 ns4 0 ns3 0 1.88816876812
Ca5 ns5 0 1e-12
Ca6 ns6 0 1e-12
Ra5 ns5 0 78.3630472463 noise=0
Ra6 ns6 0 78.3630472463 noise=0
Ga5 ns5 0 ns6 0 -1.87552614083
Ga6 ns6 0 ns5 0 1.87552614083
Ca7 ns7 0 1e-12
Ca8 ns8 0 1e-12
Ra7 ns7 0 28.6294222129 noise=0
Ra8 ns8 0 28.6294222129 noise=0
Ga7 ns7 0 ns8 0 -1.8615708713
Ga8 ns8 0 ns7 0 1.8615708713
Ca9 ns9 0 1e-12
Ca10 ns10 0 1e-12
Ra9 ns9 0 934.131832031 noise=0
Ra10 ns10 0 934.131832031 noise=0
Ga9 ns9 0 ns10 0 -1.77206208419
Ga10 ns10 0 ns9 0 1.77206208419
Ca11 ns11 0 1e-12
Ca12 ns12 0 1e-12
Ra11 ns11 0 30.3138883767 noise=0
Ra12 ns12 0 30.3138883767 noise=0
Ga11 ns11 0 ns12 0 -1.74835043081
Ga12 ns12 0 ns11 0 1.74835043081
Ca13 ns13 0 1e-12
Ca14 ns14 0 1e-12
Ra13 ns13 0 29.0014618309 noise=0
Ra14 ns14 0 29.0014618309 noise=0
Ga13 ns13 0 ns14 0 -1.68453524434
Ga14 ns14 0 ns13 0 1.68453524434
Ca15 ns15 0 1e-12
Ca16 ns16 0 1e-12
Ra15 ns15 0 608.740499085 noise=0
Ra16 ns16 0 608.740499085 noise=0
Ga15 ns15 0 ns16 0 -1.60136974681
Ga16 ns16 0 ns15 0 1.60136974681
Ca17 ns17 0 1e-12
Ca18 ns18 0 1e-12
Ra17 ns17 0 28.8457454632 noise=0
Ra18 ns18 0 28.8457454632 noise=0
Ga17 ns17 0 ns18 0 -1.57343392648
Ga18 ns18 0 ns17 0 1.57343392648
Ca19 ns19 0 1e-12
Ca20 ns20 0 1e-12
Ra19 ns19 0 27.1849571621 noise=0
Ra20 ns20 0 27.1849571621 noise=0
Ga19 ns19 0 ns20 0 -1.49976985502
Ga20 ns20 0 ns19 0 1.49976985502
Ca21 ns21 0 1e-12
Ca22 ns22 0 1e-12
Ra21 ns21 0 294.868225966 noise=0
Ra22 ns22 0 294.868225966 noise=0
Ga21 ns21 0 ns22 0 -1.43272297288
Ga22 ns22 0 ns21 0 1.43272297288
Ca23 ns23 0 1e-12
Ca24 ns24 0 1e-12
Ra23 ns23 0 24.065722504 noise=0
Ra24 ns24 0 24.065722504 noise=0
Ga23 ns23 0 ns24 0 -1.39531521009
Ga24 ns24 0 ns23 0 1.39531521009
Ca25 ns25 0 1e-12
Ca26 ns26 0 1e-12
Ra25 ns25 0 27.949811121 noise=0
Ra26 ns26 0 27.949811121 noise=0
Ga25 ns25 0 ns26 0 -1.32076031205
Ga26 ns26 0 ns25 0 1.32076031205
Ca27 ns27 0 1e-12
Ca28 ns28 0 1e-12
Ra27 ns27 0 68.9019895791 noise=0
Ra28 ns28 0 68.9019895791 noise=0
Ga27 ns27 0 ns28 0 -1.26735586041
Ga28 ns28 0 ns27 0 1.26735586041
Ca29 ns29 0 1e-12
Ca30 ns30 0 1e-12
Ra29 ns29 0 17.4920890166 noise=0
Ra30 ns30 0 17.4920890166 noise=0
Ga29 ns29 0 ns30 0 -1.21455822137
Ga30 ns30 0 ns29 0 1.21455822137
Ca31 ns31 0 1e-12
Ca32 ns32 0 1e-12
Ra31 ns31 0 23.7303485873 noise=0
Ra32 ns32 0 23.7303485873 noise=0
Ga31 ns31 0 ns32 0 -1.13110590561
Ga32 ns32 0 ns31 0 1.13110590561
Ca33 ns33 0 1e-12
Ca34 ns34 0 1e-12
Ra33 ns33 0 12.6702453574 noise=0
Ra34 ns34 0 12.6702453574 noise=0
Ga33 ns33 0 ns34 0 -1.01544529945
Ga34 ns34 0 ns33 0 1.01544529945
Ca35 ns35 0 1e-12
Ca36 ns36 0 1e-12
Ra35 ns35 0 22.4497679254 noise=0
Ra36 ns36 0 22.4497679254 noise=0
Ga35 ns35 0 ns36 0 -0.947337481808
Ga36 ns36 0 ns35 0 0.947337481808
Ca37 ns37 0 1e-12
Ca38 ns38 0 1e-12
Ra37 ns37 0 19.3969089633 noise=0
Ra38 ns38 0 19.3969089633 noise=0
Ga37 ns37 0 ns38 0 -0.828769989963
Ga38 ns38 0 ns37 0 0.828769989963
Ca39 ns39 0 1e-12
Ca40 ns40 0 1e-12
Ra39 ns39 0 28.1931334636 noise=0
Ra40 ns40 0 28.1931334636 noise=0
Ga39 ns39 0 ns40 0 -0.753040704424
Ga40 ns40 0 ns39 0 0.753040704424
Ca41 ns41 0 1e-12
Ca42 ns42 0 1e-12
Ra41 ns41 0 9.58447239365 noise=0
Ra42 ns42 0 9.58447239365 noise=0
Ga41 ns41 0 ns42 0 -0.706025240203
Ga42 ns42 0 ns41 0 0.706025240203
Ca43 ns43 0 1e-12
Ca44 ns44 0 1e-12
Ra43 ns43 0 19.2217606518 noise=0
Ra44 ns44 0 19.2217606518 noise=0
Ga43 ns43 0 ns44 0 -0.584920288579
Ga44 ns44 0 ns43 0 0.584920288579
Ca45 ns45 0 1e-12
Ca46 ns46 0 1e-12
Ra45 ns45 0 12.9186134131 noise=0
Ra46 ns46 0 12.9186134131 noise=0
Ga45 ns45 0 ns46 0 -0.451995255731
Ga46 ns46 0 ns45 0 0.451995255731
Ca47 ns47 0 1e-12
Ca48 ns48 0 1e-12
Ra47 ns47 0 14.6643586754 noise=0
Ra48 ns48 0 14.6643586754 noise=0
Ga47 ns47 0 ns48 0 -0.39239765994
Ga48 ns48 0 ns47 0 0.39239765994
Ca49 ns49 0 1e-12
Ca50 ns50 0 1e-12
Ra49 ns49 0 18.5528384969 noise=0
Ra50 ns50 0 18.5528384969 noise=0
Ga49 ns49 0 ns50 0 -0.213309922964
Ga50 ns50 0 ns49 0 0.213309922964
Ca51 ns51 0 1e-12
Ca52 ns52 0 1e-12
Ra51 ns51 0 16.425306589 noise=0
Ra52 ns52 0 16.425306589 noise=0
Ga51 ns51 0 ns52 0 -0.132506240506
Ga52 ns52 0 ns51 0 0.132506240506
Ca53 ns53 0 1e-12
Ra53 ns53 0 12.9927381247 noise=0
Ca54 ns54 0 1e-12
Ra54 ns54 0 99.3047026559 noise=0
Ca55 ns55 0 1e-12
Ca56 ns56 0 1e-12
Ra55 ns55 0 116.054358759 noise=0
Ra56 ns56 0 116.054358759 noise=0
Ga55 ns55 0 ns56 0 -0.0790828435996
Ga56 ns56 0 ns55 0 0.0790828435996
Ca57 ns57 0 1e-12
Ca58 ns58 0 1e-12
Ra57 ns57 0 0.177524466588 noise=0
Ra58 ns58 0 0.177524466588 noise=0
Ga57 ns57 0 ns58 0 -0.592192182122
Ga58 ns58 0 ns57 0 0.592192182122
Ca59 ns59 0 1e-12
Ca60 ns60 0 1e-12
Ra59 ns59 0 3.73043526058 noise=0
Ra60 ns60 0 3.73043526058 noise=0
Ga59 ns59 0 ns60 0 -1.88816876812
Ga60 ns60 0 ns59 0 1.88816876812
Ca61 ns61 0 1e-12
Ca62 ns62 0 1e-12
Ra61 ns61 0 78.3630472463 noise=0
Ra62 ns62 0 78.3630472463 noise=0
Ga61 ns61 0 ns62 0 -1.87552614083
Ga62 ns62 0 ns61 0 1.87552614083
Ca63 ns63 0 1e-12
Ca64 ns64 0 1e-12
Ra63 ns63 0 28.6294222129 noise=0
Ra64 ns64 0 28.6294222129 noise=0
Ga63 ns63 0 ns64 0 -1.8615708713
Ga64 ns64 0 ns63 0 1.8615708713
Ca65 ns65 0 1e-12
Ca66 ns66 0 1e-12
Ra65 ns65 0 934.131832031 noise=0
Ra66 ns66 0 934.131832031 noise=0
Ga65 ns65 0 ns66 0 -1.77206208419
Ga66 ns66 0 ns65 0 1.77206208419
Ca67 ns67 0 1e-12
Ca68 ns68 0 1e-12
Ra67 ns67 0 30.3138883767 noise=0
Ra68 ns68 0 30.3138883767 noise=0
Ga67 ns67 0 ns68 0 -1.74835043081
Ga68 ns68 0 ns67 0 1.74835043081
Ca69 ns69 0 1e-12
Ca70 ns70 0 1e-12
Ra69 ns69 0 29.0014618309 noise=0
Ra70 ns70 0 29.0014618309 noise=0
Ga69 ns69 0 ns70 0 -1.68453524434
Ga70 ns70 0 ns69 0 1.68453524434
Ca71 ns71 0 1e-12
Ca72 ns72 0 1e-12
Ra71 ns71 0 608.740499085 noise=0
Ra72 ns72 0 608.740499085 noise=0
Ga71 ns71 0 ns72 0 -1.60136974681
Ga72 ns72 0 ns71 0 1.60136974681
Ca73 ns73 0 1e-12
Ca74 ns74 0 1e-12
Ra73 ns73 0 28.8457454632 noise=0
Ra74 ns74 0 28.8457454632 noise=0
Ga73 ns73 0 ns74 0 -1.57343392648
Ga74 ns74 0 ns73 0 1.57343392648
Ca75 ns75 0 1e-12
Ca76 ns76 0 1e-12
Ra75 ns75 0 27.1849571621 noise=0
Ra76 ns76 0 27.1849571621 noise=0
Ga75 ns75 0 ns76 0 -1.49976985502
Ga76 ns76 0 ns75 0 1.49976985502
Ca77 ns77 0 1e-12
Ca78 ns78 0 1e-12
Ra77 ns77 0 294.868225966 noise=0
Ra78 ns78 0 294.868225966 noise=0
Ga77 ns77 0 ns78 0 -1.43272297288
Ga78 ns78 0 ns77 0 1.43272297288
Ca79 ns79 0 1e-12
Ca80 ns80 0 1e-12
Ra79 ns79 0 24.065722504 noise=0
Ra80 ns80 0 24.065722504 noise=0
Ga79 ns79 0 ns80 0 -1.39531521009
Ga80 ns80 0 ns79 0 1.39531521009
Ca81 ns81 0 1e-12
Ca82 ns82 0 1e-12
Ra81 ns81 0 27.949811121 noise=0
Ra82 ns82 0 27.949811121 noise=0
Ga81 ns81 0 ns82 0 -1.32076031205
Ga82 ns82 0 ns81 0 1.32076031205
Ca83 ns83 0 1e-12
Ca84 ns84 0 1e-12
Ra83 ns83 0 68.9019895791 noise=0
Ra84 ns84 0 68.9019895791 noise=0
Ga83 ns83 0 ns84 0 -1.26735586041
Ga84 ns84 0 ns83 0 1.26735586041
Ca85 ns85 0 1e-12
Ca86 ns86 0 1e-12
Ra85 ns85 0 17.4920890166 noise=0
Ra86 ns86 0 17.4920890166 noise=0
Ga85 ns85 0 ns86 0 -1.21455822137
Ga86 ns86 0 ns85 0 1.21455822137
Ca87 ns87 0 1e-12
Ca88 ns88 0 1e-12
Ra87 ns87 0 23.7303485873 noise=0
Ra88 ns88 0 23.7303485873 noise=0
Ga87 ns87 0 ns88 0 -1.13110590561
Ga88 ns88 0 ns87 0 1.13110590561
Ca89 ns89 0 1e-12
Ca90 ns90 0 1e-12
Ra89 ns89 0 12.6702453574 noise=0
Ra90 ns90 0 12.6702453574 noise=0
Ga89 ns89 0 ns90 0 -1.01544529945
Ga90 ns90 0 ns89 0 1.01544529945
Ca91 ns91 0 1e-12
Ca92 ns92 0 1e-12
Ra91 ns91 0 22.4497679254 noise=0
Ra92 ns92 0 22.4497679254 noise=0
Ga91 ns91 0 ns92 0 -0.947337481808
Ga92 ns92 0 ns91 0 0.947337481808
Ca93 ns93 0 1e-12
Ca94 ns94 0 1e-12
Ra93 ns93 0 19.3969089633 noise=0
Ra94 ns94 0 19.3969089633 noise=0
Ga93 ns93 0 ns94 0 -0.828769989963
Ga94 ns94 0 ns93 0 0.828769989963
Ca95 ns95 0 1e-12
Ca96 ns96 0 1e-12
Ra95 ns95 0 28.1931334636 noise=0
Ra96 ns96 0 28.1931334636 noise=0
Ga95 ns95 0 ns96 0 -0.753040704424
Ga96 ns96 0 ns95 0 0.753040704424
Ca97 ns97 0 1e-12
Ca98 ns98 0 1e-12
Ra97 ns97 0 9.58447239365 noise=0
Ra98 ns98 0 9.58447239365 noise=0
Ga97 ns97 0 ns98 0 -0.706025240203
Ga98 ns98 0 ns97 0 0.706025240203
Ca99 ns99 0 1e-12
Ca100 ns100 0 1e-12
Ra99 ns99 0 19.2217606518 noise=0
Ra100 ns100 0 19.2217606518 noise=0
Ga99 ns99 0 ns100 0 -0.584920288579
Ga100 ns100 0 ns99 0 0.584920288579
Ca101 ns101 0 1e-12
Ca102 ns102 0 1e-12
Ra101 ns101 0 12.9186134131 noise=0
Ra102 ns102 0 12.9186134131 noise=0
Ga101 ns101 0 ns102 0 -0.451995255731
Ga102 ns102 0 ns101 0 0.451995255731
Ca103 ns103 0 1e-12
Ca104 ns104 0 1e-12
Ra103 ns103 0 14.6643586754 noise=0
Ra104 ns104 0 14.6643586754 noise=0
Ga103 ns103 0 ns104 0 -0.39239765994
Ga104 ns104 0 ns103 0 0.39239765994
Ca105 ns105 0 1e-12
Ca106 ns106 0 1e-12
Ra105 ns105 0 18.5528384969 noise=0
Ra106 ns106 0 18.5528384969 noise=0
Ga105 ns105 0 ns106 0 -0.213309922964
Ga106 ns106 0 ns105 0 0.213309922964
Ca107 ns107 0 1e-12
Ca108 ns108 0 1e-12
Ra107 ns107 0 16.425306589 noise=0
Ra108 ns108 0 16.425306589 noise=0
Ga107 ns107 0 ns108 0 -0.132506240506
Ga108 ns108 0 ns107 0 0.132506240506
Ca109 ns109 0 1e-12
Ra109 ns109 0 12.9927381247 noise=0
Ca110 ns110 0 1e-12
Ra110 ns110 0 99.3047026559 noise=0
Ca111 ns111 0 1e-12
Ca112 ns112 0 1e-12
Ra111 ns111 0 116.054358759 noise=0
Ra112 ns112 0 116.054358759 noise=0
Ga111 ns111 0 ns112 0 -0.0790828435996
Ga112 ns112 0 ns111 0 0.0790828435996
Ca113 ns113 0 1e-12
Ca114 ns114 0 1e-12
Ra113 ns113 0 0.177524466588 noise=0
Ra114 ns114 0 0.177524466588 noise=0
Ga113 ns113 0 ns114 0 -0.592192182122
Ga114 ns114 0 ns113 0 0.592192182122
Ca115 ns115 0 1e-12
Ca116 ns116 0 1e-12
Ra115 ns115 0 3.73043526058 noise=0
Ra116 ns116 0 3.73043526058 noise=0
Ga115 ns115 0 ns116 0 -1.88816876812
Ga116 ns116 0 ns115 0 1.88816876812
Ca117 ns117 0 1e-12
Ca118 ns118 0 1e-12
Ra117 ns117 0 78.3630472463 noise=0
Ra118 ns118 0 78.3630472463 noise=0
Ga117 ns117 0 ns118 0 -1.87552614083
Ga118 ns118 0 ns117 0 1.87552614083
Ca119 ns119 0 1e-12
Ca120 ns120 0 1e-12
Ra119 ns119 0 28.6294222129 noise=0
Ra120 ns120 0 28.6294222129 noise=0
Ga119 ns119 0 ns120 0 -1.8615708713
Ga120 ns120 0 ns119 0 1.8615708713
Ca121 ns121 0 1e-12
Ca122 ns122 0 1e-12
Ra121 ns121 0 934.131832031 noise=0
Ra122 ns122 0 934.131832031 noise=0
Ga121 ns121 0 ns122 0 -1.77206208419
Ga122 ns122 0 ns121 0 1.77206208419
Ca123 ns123 0 1e-12
Ca124 ns124 0 1e-12
Ra123 ns123 0 30.3138883767 noise=0
Ra124 ns124 0 30.3138883767 noise=0
Ga123 ns123 0 ns124 0 -1.74835043081
Ga124 ns124 0 ns123 0 1.74835043081
Ca125 ns125 0 1e-12
Ca126 ns126 0 1e-12
Ra125 ns125 0 29.0014618309 noise=0
Ra126 ns126 0 29.0014618309 noise=0
Ga125 ns125 0 ns126 0 -1.68453524434
Ga126 ns126 0 ns125 0 1.68453524434
Ca127 ns127 0 1e-12
Ca128 ns128 0 1e-12
Ra127 ns127 0 608.740499085 noise=0
Ra128 ns128 0 608.740499085 noise=0
Ga127 ns127 0 ns128 0 -1.60136974681
Ga128 ns128 0 ns127 0 1.60136974681
Ca129 ns129 0 1e-12
Ca130 ns130 0 1e-12
Ra129 ns129 0 28.8457454632 noise=0
Ra130 ns130 0 28.8457454632 noise=0
Ga129 ns129 0 ns130 0 -1.57343392648
Ga130 ns130 0 ns129 0 1.57343392648
Ca131 ns131 0 1e-12
Ca132 ns132 0 1e-12
Ra131 ns131 0 27.1849571621 noise=0
Ra132 ns132 0 27.1849571621 noise=0
Ga131 ns131 0 ns132 0 -1.49976985502
Ga132 ns132 0 ns131 0 1.49976985502
Ca133 ns133 0 1e-12
Ca134 ns134 0 1e-12
Ra133 ns133 0 294.868225966 noise=0
Ra134 ns134 0 294.868225966 noise=0
Ga133 ns133 0 ns134 0 -1.43272297288
Ga134 ns134 0 ns133 0 1.43272297288
Ca135 ns135 0 1e-12
Ca136 ns136 0 1e-12
Ra135 ns135 0 24.065722504 noise=0
Ra136 ns136 0 24.065722504 noise=0
Ga135 ns135 0 ns136 0 -1.39531521009
Ga136 ns136 0 ns135 0 1.39531521009
Ca137 ns137 0 1e-12
Ca138 ns138 0 1e-12
Ra137 ns137 0 27.949811121 noise=0
Ra138 ns138 0 27.949811121 noise=0
Ga137 ns137 0 ns138 0 -1.32076031205
Ga138 ns138 0 ns137 0 1.32076031205
Ca139 ns139 0 1e-12
Ca140 ns140 0 1e-12
Ra139 ns139 0 68.9019895791 noise=0
Ra140 ns140 0 68.9019895791 noise=0
Ga139 ns139 0 ns140 0 -1.26735586041
Ga140 ns140 0 ns139 0 1.26735586041
Ca141 ns141 0 1e-12
Ca142 ns142 0 1e-12
Ra141 ns141 0 17.4920890166 noise=0
Ra142 ns142 0 17.4920890166 noise=0
Ga141 ns141 0 ns142 0 -1.21455822137
Ga142 ns142 0 ns141 0 1.21455822137
Ca143 ns143 0 1e-12
Ca144 ns144 0 1e-12
Ra143 ns143 0 23.7303485873 noise=0
Ra144 ns144 0 23.7303485873 noise=0
Ga143 ns143 0 ns144 0 -1.13110590561
Ga144 ns144 0 ns143 0 1.13110590561
Ca145 ns145 0 1e-12
Ca146 ns146 0 1e-12
Ra145 ns145 0 12.6702453574 noise=0
Ra146 ns146 0 12.6702453574 noise=0
Ga145 ns145 0 ns146 0 -1.01544529945
Ga146 ns146 0 ns145 0 1.01544529945
Ca147 ns147 0 1e-12
Ca148 ns148 0 1e-12
Ra147 ns147 0 22.4497679254 noise=0
Ra148 ns148 0 22.4497679254 noise=0
Ga147 ns147 0 ns148 0 -0.947337481808
Ga148 ns148 0 ns147 0 0.947337481808
Ca149 ns149 0 1e-12
Ca150 ns150 0 1e-12
Ra149 ns149 0 19.3969089633 noise=0
Ra150 ns150 0 19.3969089633 noise=0
Ga149 ns149 0 ns150 0 -0.828769989963
Ga150 ns150 0 ns149 0 0.828769989963
Ca151 ns151 0 1e-12
Ca152 ns152 0 1e-12
Ra151 ns151 0 28.1931334636 noise=0
Ra152 ns152 0 28.1931334636 noise=0
Ga151 ns151 0 ns152 0 -0.753040704424
Ga152 ns152 0 ns151 0 0.753040704424
Ca153 ns153 0 1e-12
Ca154 ns154 0 1e-12
Ra153 ns153 0 9.58447239365 noise=0
Ra154 ns154 0 9.58447239365 noise=0
Ga153 ns153 0 ns154 0 -0.706025240203
Ga154 ns154 0 ns153 0 0.706025240203
Ca155 ns155 0 1e-12
Ca156 ns156 0 1e-12
Ra155 ns155 0 19.2217606518 noise=0
Ra156 ns156 0 19.2217606518 noise=0
Ga155 ns155 0 ns156 0 -0.584920288579
Ga156 ns156 0 ns155 0 0.584920288579
Ca157 ns157 0 1e-12
Ca158 ns158 0 1e-12
Ra157 ns157 0 12.9186134131 noise=0
Ra158 ns158 0 12.9186134131 noise=0
Ga157 ns157 0 ns158 0 -0.451995255731
Ga158 ns158 0 ns157 0 0.451995255731
Ca159 ns159 0 1e-12
Ca160 ns160 0 1e-12
Ra159 ns159 0 14.6643586754 noise=0
Ra160 ns160 0 14.6643586754 noise=0
Ga159 ns159 0 ns160 0 -0.39239765994
Ga160 ns160 0 ns159 0 0.39239765994
Ca161 ns161 0 1e-12
Ca162 ns162 0 1e-12
Ra161 ns161 0 18.5528384969 noise=0
Ra162 ns162 0 18.5528384969 noise=0
Ga161 ns161 0 ns162 0 -0.213309922964
Ga162 ns162 0 ns161 0 0.213309922964
Ca163 ns163 0 1e-12
Ca164 ns164 0 1e-12
Ra163 ns163 0 16.425306589 noise=0
Ra164 ns164 0 16.425306589 noise=0
Ga163 ns163 0 ns164 0 -0.132506240506
Ga164 ns164 0 ns163 0 0.132506240506
Ca165 ns165 0 1e-12
Ra165 ns165 0 12.9927381247 noise=0
Ca166 ns166 0 1e-12
Ra166 ns166 0 99.3047026559 noise=0
Ca167 ns167 0 1e-12
Ca168 ns168 0 1e-12
Ra167 ns167 0 116.054358759 noise=0
Ra168 ns168 0 116.054358759 noise=0
Ga167 ns167 0 ns168 0 -0.0790828435996
Ga168 ns168 0 ns167 0 0.0790828435996
Ca169 ns169 0 1e-12
Ca170 ns170 0 1e-12
Ra169 ns169 0 0.177524466588 noise=0
Ra170 ns170 0 0.177524466588 noise=0
Ga169 ns169 0 ns170 0 -0.592192182122
Ga170 ns170 0 ns169 0 0.592192182122
Ca171 ns171 0 1e-12
Ca172 ns172 0 1e-12
Ra171 ns171 0 3.73043526058 noise=0
Ra172 ns172 0 3.73043526058 noise=0
Ga171 ns171 0 ns172 0 -1.88816876812
Ga172 ns172 0 ns171 0 1.88816876812
Ca173 ns173 0 1e-12
Ca174 ns174 0 1e-12
Ra173 ns173 0 78.3630472463 noise=0
Ra174 ns174 0 78.3630472463 noise=0
Ga173 ns173 0 ns174 0 -1.87552614083
Ga174 ns174 0 ns173 0 1.87552614083
Ca175 ns175 0 1e-12
Ca176 ns176 0 1e-12
Ra175 ns175 0 28.6294222129 noise=0
Ra176 ns176 0 28.6294222129 noise=0
Ga175 ns175 0 ns176 0 -1.8615708713
Ga176 ns176 0 ns175 0 1.8615708713
Ca177 ns177 0 1e-12
Ca178 ns178 0 1e-12
Ra177 ns177 0 934.131832031 noise=0
Ra178 ns178 0 934.131832031 noise=0
Ga177 ns177 0 ns178 0 -1.77206208419
Ga178 ns178 0 ns177 0 1.77206208419
Ca179 ns179 0 1e-12
Ca180 ns180 0 1e-12
Ra179 ns179 0 30.3138883767 noise=0
Ra180 ns180 0 30.3138883767 noise=0
Ga179 ns179 0 ns180 0 -1.74835043081
Ga180 ns180 0 ns179 0 1.74835043081
Ca181 ns181 0 1e-12
Ca182 ns182 0 1e-12
Ra181 ns181 0 29.0014618309 noise=0
Ra182 ns182 0 29.0014618309 noise=0
Ga181 ns181 0 ns182 0 -1.68453524434
Ga182 ns182 0 ns181 0 1.68453524434
Ca183 ns183 0 1e-12
Ca184 ns184 0 1e-12
Ra183 ns183 0 608.740499085 noise=0
Ra184 ns184 0 608.740499085 noise=0
Ga183 ns183 0 ns184 0 -1.60136974681
Ga184 ns184 0 ns183 0 1.60136974681
Ca185 ns185 0 1e-12
Ca186 ns186 0 1e-12
Ra185 ns185 0 28.8457454632 noise=0
Ra186 ns186 0 28.8457454632 noise=0
Ga185 ns185 0 ns186 0 -1.57343392648
Ga186 ns186 0 ns185 0 1.57343392648
Ca187 ns187 0 1e-12
Ca188 ns188 0 1e-12
Ra187 ns187 0 27.1849571621 noise=0
Ra188 ns188 0 27.1849571621 noise=0
Ga187 ns187 0 ns188 0 -1.49976985502
Ga188 ns188 0 ns187 0 1.49976985502
Ca189 ns189 0 1e-12
Ca190 ns190 0 1e-12
Ra189 ns189 0 294.868225966 noise=0
Ra190 ns190 0 294.868225966 noise=0
Ga189 ns189 0 ns190 0 -1.43272297288
Ga190 ns190 0 ns189 0 1.43272297288
Ca191 ns191 0 1e-12
Ca192 ns192 0 1e-12
Ra191 ns191 0 24.065722504 noise=0
Ra192 ns192 0 24.065722504 noise=0
Ga191 ns191 0 ns192 0 -1.39531521009
Ga192 ns192 0 ns191 0 1.39531521009
Ca193 ns193 0 1e-12
Ca194 ns194 0 1e-12
Ra193 ns193 0 27.949811121 noise=0
Ra194 ns194 0 27.949811121 noise=0
Ga193 ns193 0 ns194 0 -1.32076031205
Ga194 ns194 0 ns193 0 1.32076031205
Ca195 ns195 0 1e-12
Ca196 ns196 0 1e-12
Ra195 ns195 0 68.9019895791 noise=0
Ra196 ns196 0 68.9019895791 noise=0
Ga195 ns195 0 ns196 0 -1.26735586041
Ga196 ns196 0 ns195 0 1.26735586041
Ca197 ns197 0 1e-12
Ca198 ns198 0 1e-12
Ra197 ns197 0 17.4920890166 noise=0
Ra198 ns198 0 17.4920890166 noise=0
Ga197 ns197 0 ns198 0 -1.21455822137
Ga198 ns198 0 ns197 0 1.21455822137
Ca199 ns199 0 1e-12
Ca200 ns200 0 1e-12
Ra199 ns199 0 23.7303485873 noise=0
Ra200 ns200 0 23.7303485873 noise=0
Ga199 ns199 0 ns200 0 -1.13110590561
Ga200 ns200 0 ns199 0 1.13110590561
Ca201 ns201 0 1e-12
Ca202 ns202 0 1e-12
Ra201 ns201 0 12.6702453574 noise=0
Ra202 ns202 0 12.6702453574 noise=0
Ga201 ns201 0 ns202 0 -1.01544529945
Ga202 ns202 0 ns201 0 1.01544529945
Ca203 ns203 0 1e-12
Ca204 ns204 0 1e-12
Ra203 ns203 0 22.4497679254 noise=0
Ra204 ns204 0 22.4497679254 noise=0
Ga203 ns203 0 ns204 0 -0.947337481808
Ga204 ns204 0 ns203 0 0.947337481808
Ca205 ns205 0 1e-12
Ca206 ns206 0 1e-12
Ra205 ns205 0 19.3969089633 noise=0
Ra206 ns206 0 19.3969089633 noise=0
Ga205 ns205 0 ns206 0 -0.828769989963
Ga206 ns206 0 ns205 0 0.828769989963
Ca207 ns207 0 1e-12
Ca208 ns208 0 1e-12
Ra207 ns207 0 28.1931334636 noise=0
Ra208 ns208 0 28.1931334636 noise=0
Ga207 ns207 0 ns208 0 -0.753040704424
Ga208 ns208 0 ns207 0 0.753040704424
Ca209 ns209 0 1e-12
Ca210 ns210 0 1e-12
Ra209 ns209 0 9.58447239365 noise=0
Ra210 ns210 0 9.58447239365 noise=0
Ga209 ns209 0 ns210 0 -0.706025240203
Ga210 ns210 0 ns209 0 0.706025240203
Ca211 ns211 0 1e-12
Ca212 ns212 0 1e-12
Ra211 ns211 0 19.2217606518 noise=0
Ra212 ns212 0 19.2217606518 noise=0
Ga211 ns211 0 ns212 0 -0.584920288579
Ga212 ns212 0 ns211 0 0.584920288579
Ca213 ns213 0 1e-12
Ca214 ns214 0 1e-12
Ra213 ns213 0 12.9186134131 noise=0
Ra214 ns214 0 12.9186134131 noise=0
Ga213 ns213 0 ns214 0 -0.451995255731
Ga214 ns214 0 ns213 0 0.451995255731
Ca215 ns215 0 1e-12
Ca216 ns216 0 1e-12
Ra215 ns215 0 14.6643586754 noise=0
Ra216 ns216 0 14.6643586754 noise=0
Ga215 ns215 0 ns216 0 -0.39239765994
Ga216 ns216 0 ns215 0 0.39239765994
Ca217 ns217 0 1e-12
Ca218 ns218 0 1e-12
Ra217 ns217 0 18.5528384969 noise=0
Ra218 ns218 0 18.5528384969 noise=0
Ga217 ns217 0 ns218 0 -0.213309922964
Ga218 ns218 0 ns217 0 0.213309922964
Ca219 ns219 0 1e-12
Ca220 ns220 0 1e-12
Ra219 ns219 0 16.425306589 noise=0
Ra220 ns220 0 16.425306589 noise=0
Ga219 ns219 0 ns220 0 -0.132506240506
Ga220 ns220 0 ns219 0 0.132506240506
Ca221 ns221 0 1e-12
Ra221 ns221 0 12.9927381247 noise=0
Ca222 ns222 0 1e-12
Ra222 ns222 0 99.3047026559 noise=0
Ca223 ns223 0 1e-12
Ca224 ns224 0 1e-12
Ra223 ns223 0 116.054358759 noise=0
Ra224 ns224 0 116.054358759 noise=0
Ga223 ns223 0 ns224 0 -0.0790828435996
Ga224 ns224 0 ns223 0 0.0790828435996
Ca225 ns225 0 1e-12
Ca226 ns226 0 1e-12
Ra225 ns225 0 0.177524466588 noise=0
Ra226 ns226 0 0.177524466588 noise=0
Ga225 ns225 0 ns226 0 -0.592192182122
Ga226 ns226 0 ns225 0 0.592192182122
Ca227 ns227 0 1e-12
Ca228 ns228 0 1e-12
Ra227 ns227 0 3.73043526058 noise=0
Ra228 ns228 0 3.73043526058 noise=0
Ga227 ns227 0 ns228 0 -1.88816876812
Ga228 ns228 0 ns227 0 1.88816876812
Ca229 ns229 0 1e-12
Ca230 ns230 0 1e-12
Ra229 ns229 0 78.3630472463 noise=0
Ra230 ns230 0 78.3630472463 noise=0
Ga229 ns229 0 ns230 0 -1.87552614083
Ga230 ns230 0 ns229 0 1.87552614083
Ca231 ns231 0 1e-12
Ca232 ns232 0 1e-12
Ra231 ns231 0 28.6294222129 noise=0
Ra232 ns232 0 28.6294222129 noise=0
Ga231 ns231 0 ns232 0 -1.8615708713
Ga232 ns232 0 ns231 0 1.8615708713
Ca233 ns233 0 1e-12
Ca234 ns234 0 1e-12
Ra233 ns233 0 934.131832031 noise=0
Ra234 ns234 0 934.131832031 noise=0
Ga233 ns233 0 ns234 0 -1.77206208419
Ga234 ns234 0 ns233 0 1.77206208419
Ca235 ns235 0 1e-12
Ca236 ns236 0 1e-12
Ra235 ns235 0 30.3138883767 noise=0
Ra236 ns236 0 30.3138883767 noise=0
Ga235 ns235 0 ns236 0 -1.74835043081
Ga236 ns236 0 ns235 0 1.74835043081
Ca237 ns237 0 1e-12
Ca238 ns238 0 1e-12
Ra237 ns237 0 29.0014618309 noise=0
Ra238 ns238 0 29.0014618309 noise=0
Ga237 ns237 0 ns238 0 -1.68453524434
Ga238 ns238 0 ns237 0 1.68453524434
Ca239 ns239 0 1e-12
Ca240 ns240 0 1e-12
Ra239 ns239 0 608.740499085 noise=0
Ra240 ns240 0 608.740499085 noise=0
Ga239 ns239 0 ns240 0 -1.60136974681
Ga240 ns240 0 ns239 0 1.60136974681
Ca241 ns241 0 1e-12
Ca242 ns242 0 1e-12
Ra241 ns241 0 28.8457454632 noise=0
Ra242 ns242 0 28.8457454632 noise=0
Ga241 ns241 0 ns242 0 -1.57343392648
Ga242 ns242 0 ns241 0 1.57343392648
Ca243 ns243 0 1e-12
Ca244 ns244 0 1e-12
Ra243 ns243 0 27.1849571621 noise=0
Ra244 ns244 0 27.1849571621 noise=0
Ga243 ns243 0 ns244 0 -1.49976985502
Ga244 ns244 0 ns243 0 1.49976985502
Ca245 ns245 0 1e-12
Ca246 ns246 0 1e-12
Ra245 ns245 0 294.868225966 noise=0
Ra246 ns246 0 294.868225966 noise=0
Ga245 ns245 0 ns246 0 -1.43272297288
Ga246 ns246 0 ns245 0 1.43272297288
Ca247 ns247 0 1e-12
Ca248 ns248 0 1e-12
Ra247 ns247 0 24.065722504 noise=0
Ra248 ns248 0 24.065722504 noise=0
Ga247 ns247 0 ns248 0 -1.39531521009
Ga248 ns248 0 ns247 0 1.39531521009
Ca249 ns249 0 1e-12
Ca250 ns250 0 1e-12
Ra249 ns249 0 27.949811121 noise=0
Ra250 ns250 0 27.949811121 noise=0
Ga249 ns249 0 ns250 0 -1.32076031205
Ga250 ns250 0 ns249 0 1.32076031205
Ca251 ns251 0 1e-12
Ca252 ns252 0 1e-12
Ra251 ns251 0 68.9019895791 noise=0
Ra252 ns252 0 68.9019895791 noise=0
Ga251 ns251 0 ns252 0 -1.26735586041
Ga252 ns252 0 ns251 0 1.26735586041
Ca253 ns253 0 1e-12
Ca254 ns254 0 1e-12
Ra253 ns253 0 17.4920890166 noise=0
Ra254 ns254 0 17.4920890166 noise=0
Ga253 ns253 0 ns254 0 -1.21455822137
Ga254 ns254 0 ns253 0 1.21455822137
Ca255 ns255 0 1e-12
Ca256 ns256 0 1e-12
Ra255 ns255 0 23.7303485873 noise=0
Ra256 ns256 0 23.7303485873 noise=0
Ga255 ns255 0 ns256 0 -1.13110590561
Ga256 ns256 0 ns255 0 1.13110590561
Ca257 ns257 0 1e-12
Ca258 ns258 0 1e-12
Ra257 ns257 0 12.6702453574 noise=0
Ra258 ns258 0 12.6702453574 noise=0
Ga257 ns257 0 ns258 0 -1.01544529945
Ga258 ns258 0 ns257 0 1.01544529945
Ca259 ns259 0 1e-12
Ca260 ns260 0 1e-12
Ra259 ns259 0 22.4497679254 noise=0
Ra260 ns260 0 22.4497679254 noise=0
Ga259 ns259 0 ns260 0 -0.947337481808
Ga260 ns260 0 ns259 0 0.947337481808
Ca261 ns261 0 1e-12
Ca262 ns262 0 1e-12
Ra261 ns261 0 19.3969089633 noise=0
Ra262 ns262 0 19.3969089633 noise=0
Ga261 ns261 0 ns262 0 -0.828769989963
Ga262 ns262 0 ns261 0 0.828769989963
Ca263 ns263 0 1e-12
Ca264 ns264 0 1e-12
Ra263 ns263 0 28.1931334636 noise=0
Ra264 ns264 0 28.1931334636 noise=0
Ga263 ns263 0 ns264 0 -0.753040704424
Ga264 ns264 0 ns263 0 0.753040704424
Ca265 ns265 0 1e-12
Ca266 ns266 0 1e-12
Ra265 ns265 0 9.58447239365 noise=0
Ra266 ns266 0 9.58447239365 noise=0
Ga265 ns265 0 ns266 0 -0.706025240203
Ga266 ns266 0 ns265 0 0.706025240203
Ca267 ns267 0 1e-12
Ca268 ns268 0 1e-12
Ra267 ns267 0 19.2217606518 noise=0
Ra268 ns268 0 19.2217606518 noise=0
Ga267 ns267 0 ns268 0 -0.584920288579
Ga268 ns268 0 ns267 0 0.584920288579
Ca269 ns269 0 1e-12
Ca270 ns270 0 1e-12
Ra269 ns269 0 12.9186134131 noise=0
Ra270 ns270 0 12.9186134131 noise=0
Ga269 ns269 0 ns270 0 -0.451995255731
Ga270 ns270 0 ns269 0 0.451995255731
Ca271 ns271 0 1e-12
Ca272 ns272 0 1e-12
Ra271 ns271 0 14.6643586754 noise=0
Ra272 ns272 0 14.6643586754 noise=0
Ga271 ns271 0 ns272 0 -0.39239765994
Ga272 ns272 0 ns271 0 0.39239765994
Ca273 ns273 0 1e-12
Ca274 ns274 0 1e-12
Ra273 ns273 0 18.5528384969 noise=0
Ra274 ns274 0 18.5528384969 noise=0
Ga273 ns273 0 ns274 0 -0.213309922964
Ga274 ns274 0 ns273 0 0.213309922964
Ca275 ns275 0 1e-12
Ca276 ns276 0 1e-12
Ra275 ns275 0 16.425306589 noise=0
Ra276 ns276 0 16.425306589 noise=0
Ga275 ns275 0 ns276 0 -0.132506240506
Ga276 ns276 0 ns275 0 0.132506240506
Ca277 ns277 0 1e-12
Ra277 ns277 0 12.9927381247 noise=0
Ca278 ns278 0 1e-12
Ra278 ns278 0 99.3047026559 noise=0
Ca279 ns279 0 1e-12
Ca280 ns280 0 1e-12
Ra279 ns279 0 116.054358759 noise=0
Ra280 ns280 0 116.054358759 noise=0
Ga279 ns279 0 ns280 0 -0.0790828435996
Ga280 ns280 0 ns279 0 0.0790828435996
Ca281 ns281 0 1e-12
Ca282 ns282 0 1e-12
Ra281 ns281 0 0.177524466588 noise=0
Ra282 ns282 0 0.177524466588 noise=0
Ga281 ns281 0 ns282 0 -0.592192182122
Ga282 ns282 0 ns281 0 0.592192182122
Ca283 ns283 0 1e-12
Ca284 ns284 0 1e-12
Ra283 ns283 0 3.73043526058 noise=0
Ra284 ns284 0 3.73043526058 noise=0
Ga283 ns283 0 ns284 0 -1.88816876812
Ga284 ns284 0 ns283 0 1.88816876812
Ca285 ns285 0 1e-12
Ca286 ns286 0 1e-12
Ra285 ns285 0 78.3630472463 noise=0
Ra286 ns286 0 78.3630472463 noise=0
Ga285 ns285 0 ns286 0 -1.87552614083
Ga286 ns286 0 ns285 0 1.87552614083
Ca287 ns287 0 1e-12
Ca288 ns288 0 1e-12
Ra287 ns287 0 28.6294222129 noise=0
Ra288 ns288 0 28.6294222129 noise=0
Ga287 ns287 0 ns288 0 -1.8615708713
Ga288 ns288 0 ns287 0 1.8615708713
Ca289 ns289 0 1e-12
Ca290 ns290 0 1e-12
Ra289 ns289 0 934.131832031 noise=0
Ra290 ns290 0 934.131832031 noise=0
Ga289 ns289 0 ns290 0 -1.77206208419
Ga290 ns290 0 ns289 0 1.77206208419
Ca291 ns291 0 1e-12
Ca292 ns292 0 1e-12
Ra291 ns291 0 30.3138883767 noise=0
Ra292 ns292 0 30.3138883767 noise=0
Ga291 ns291 0 ns292 0 -1.74835043081
Ga292 ns292 0 ns291 0 1.74835043081
Ca293 ns293 0 1e-12
Ca294 ns294 0 1e-12
Ra293 ns293 0 29.0014618309 noise=0
Ra294 ns294 0 29.0014618309 noise=0
Ga293 ns293 0 ns294 0 -1.68453524434
Ga294 ns294 0 ns293 0 1.68453524434
Ca295 ns295 0 1e-12
Ca296 ns296 0 1e-12
Ra295 ns295 0 608.740499085 noise=0
Ra296 ns296 0 608.740499085 noise=0
Ga295 ns295 0 ns296 0 -1.60136974681
Ga296 ns296 0 ns295 0 1.60136974681
Ca297 ns297 0 1e-12
Ca298 ns298 0 1e-12
Ra297 ns297 0 28.8457454632 noise=0
Ra298 ns298 0 28.8457454632 noise=0
Ga297 ns297 0 ns298 0 -1.57343392648
Ga298 ns298 0 ns297 0 1.57343392648
Ca299 ns299 0 1e-12
Ca300 ns300 0 1e-12
Ra299 ns299 0 27.1849571621 noise=0
Ra300 ns300 0 27.1849571621 noise=0
Ga299 ns299 0 ns300 0 -1.49976985502
Ga300 ns300 0 ns299 0 1.49976985502
Ca301 ns301 0 1e-12
Ca302 ns302 0 1e-12
Ra301 ns301 0 294.868225966 noise=0
Ra302 ns302 0 294.868225966 noise=0
Ga301 ns301 0 ns302 0 -1.43272297288
Ga302 ns302 0 ns301 0 1.43272297288
Ca303 ns303 0 1e-12
Ca304 ns304 0 1e-12
Ra303 ns303 0 24.065722504 noise=0
Ra304 ns304 0 24.065722504 noise=0
Ga303 ns303 0 ns304 0 -1.39531521009
Ga304 ns304 0 ns303 0 1.39531521009
Ca305 ns305 0 1e-12
Ca306 ns306 0 1e-12
Ra305 ns305 0 27.949811121 noise=0
Ra306 ns306 0 27.949811121 noise=0
Ga305 ns305 0 ns306 0 -1.32076031205
Ga306 ns306 0 ns305 0 1.32076031205
Ca307 ns307 0 1e-12
Ca308 ns308 0 1e-12
Ra307 ns307 0 68.9019895791 noise=0
Ra308 ns308 0 68.9019895791 noise=0
Ga307 ns307 0 ns308 0 -1.26735586041
Ga308 ns308 0 ns307 0 1.26735586041
Ca309 ns309 0 1e-12
Ca310 ns310 0 1e-12
Ra309 ns309 0 17.4920890166 noise=0
Ra310 ns310 0 17.4920890166 noise=0
Ga309 ns309 0 ns310 0 -1.21455822137
Ga310 ns310 0 ns309 0 1.21455822137
Ca311 ns311 0 1e-12
Ca312 ns312 0 1e-12
Ra311 ns311 0 23.7303485873 noise=0
Ra312 ns312 0 23.7303485873 noise=0
Ga311 ns311 0 ns312 0 -1.13110590561
Ga312 ns312 0 ns311 0 1.13110590561
Ca313 ns313 0 1e-12
Ca314 ns314 0 1e-12
Ra313 ns313 0 12.6702453574 noise=0
Ra314 ns314 0 12.6702453574 noise=0
Ga313 ns313 0 ns314 0 -1.01544529945
Ga314 ns314 0 ns313 0 1.01544529945
Ca315 ns315 0 1e-12
Ca316 ns316 0 1e-12
Ra315 ns315 0 22.4497679254 noise=0
Ra316 ns316 0 22.4497679254 noise=0
Ga315 ns315 0 ns316 0 -0.947337481808
Ga316 ns316 0 ns315 0 0.947337481808
Ca317 ns317 0 1e-12
Ca318 ns318 0 1e-12
Ra317 ns317 0 19.3969089633 noise=0
Ra318 ns318 0 19.3969089633 noise=0
Ga317 ns317 0 ns318 0 -0.828769989963
Ga318 ns318 0 ns317 0 0.828769989963
Ca319 ns319 0 1e-12
Ca320 ns320 0 1e-12
Ra319 ns319 0 28.1931334636 noise=0
Ra320 ns320 0 28.1931334636 noise=0
Ga319 ns319 0 ns320 0 -0.753040704424
Ga320 ns320 0 ns319 0 0.753040704424
Ca321 ns321 0 1e-12
Ca322 ns322 0 1e-12
Ra321 ns321 0 9.58447239365 noise=0
Ra322 ns322 0 9.58447239365 noise=0
Ga321 ns321 0 ns322 0 -0.706025240203
Ga322 ns322 0 ns321 0 0.706025240203
Ca323 ns323 0 1e-12
Ca324 ns324 0 1e-12
Ra323 ns323 0 19.2217606518 noise=0
Ra324 ns324 0 19.2217606518 noise=0
Ga323 ns323 0 ns324 0 -0.584920288579
Ga324 ns324 0 ns323 0 0.584920288579
Ca325 ns325 0 1e-12
Ca326 ns326 0 1e-12
Ra325 ns325 0 12.9186134131 noise=0
Ra326 ns326 0 12.9186134131 noise=0
Ga325 ns325 0 ns326 0 -0.451995255731
Ga326 ns326 0 ns325 0 0.451995255731
Ca327 ns327 0 1e-12
Ca328 ns328 0 1e-12
Ra327 ns327 0 14.6643586754 noise=0
Ra328 ns328 0 14.6643586754 noise=0
Ga327 ns327 0 ns328 0 -0.39239765994
Ga328 ns328 0 ns327 0 0.39239765994
Ca329 ns329 0 1e-12
Ca330 ns330 0 1e-12
Ra329 ns329 0 18.5528384969 noise=0
Ra330 ns330 0 18.5528384969 noise=0
Ga329 ns329 0 ns330 0 -0.213309922964
Ga330 ns330 0 ns329 0 0.213309922964
Ca331 ns331 0 1e-12
Ca332 ns332 0 1e-12
Ra331 ns331 0 16.425306589 noise=0
Ra332 ns332 0 16.425306589 noise=0
Ga331 ns331 0 ns332 0 -0.132506240506
Ga332 ns332 0 ns331 0 0.132506240506
Ca333 ns333 0 1e-12
Ra333 ns333 0 12.9927381247 noise=0
Ca334 ns334 0 1e-12
Ra334 ns334 0 99.3047026559 noise=0
Ca335 ns335 0 1e-12
Ca336 ns336 0 1e-12
Ra335 ns335 0 116.054358759 noise=0
Ra336 ns336 0 116.054358759 noise=0
Ga335 ns335 0 ns336 0 -0.0790828435996
Ga336 ns336 0 ns335 0 0.0790828435996
Ca337 ns337 0 1e-12
Ca338 ns338 0 1e-12
Ra337 ns337 0 0.177524466588 noise=0
Ra338 ns338 0 0.177524466588 noise=0
Ga337 ns337 0 ns338 0 -0.592192182122
Ga338 ns338 0 ns337 0 0.592192182122
Ca339 ns339 0 1e-12
Ca340 ns340 0 1e-12
Ra339 ns339 0 3.73043526058 noise=0
Ra340 ns340 0 3.73043526058 noise=0
Ga339 ns339 0 ns340 0 -1.88816876812
Ga340 ns340 0 ns339 0 1.88816876812
Ca341 ns341 0 1e-12
Ca342 ns342 0 1e-12
Ra341 ns341 0 78.3630472463 noise=0
Ra342 ns342 0 78.3630472463 noise=0
Ga341 ns341 0 ns342 0 -1.87552614083
Ga342 ns342 0 ns341 0 1.87552614083
Ca343 ns343 0 1e-12
Ca344 ns344 0 1e-12
Ra343 ns343 0 28.6294222129 noise=0
Ra344 ns344 0 28.6294222129 noise=0
Ga343 ns343 0 ns344 0 -1.8615708713
Ga344 ns344 0 ns343 0 1.8615708713
Ca345 ns345 0 1e-12
Ca346 ns346 0 1e-12
Ra345 ns345 0 934.131832031 noise=0
Ra346 ns346 0 934.131832031 noise=0
Ga345 ns345 0 ns346 0 -1.77206208419
Ga346 ns346 0 ns345 0 1.77206208419
Ca347 ns347 0 1e-12
Ca348 ns348 0 1e-12
Ra347 ns347 0 30.3138883767 noise=0
Ra348 ns348 0 30.3138883767 noise=0
Ga347 ns347 0 ns348 0 -1.74835043081
Ga348 ns348 0 ns347 0 1.74835043081
Ca349 ns349 0 1e-12
Ca350 ns350 0 1e-12
Ra349 ns349 0 29.0014618309 noise=0
Ra350 ns350 0 29.0014618309 noise=0
Ga349 ns349 0 ns350 0 -1.68453524434
Ga350 ns350 0 ns349 0 1.68453524434
Ca351 ns351 0 1e-12
Ca352 ns352 0 1e-12
Ra351 ns351 0 608.740499085 noise=0
Ra352 ns352 0 608.740499085 noise=0
Ga351 ns351 0 ns352 0 -1.60136974681
Ga352 ns352 0 ns351 0 1.60136974681
Ca353 ns353 0 1e-12
Ca354 ns354 0 1e-12
Ra353 ns353 0 28.8457454632 noise=0
Ra354 ns354 0 28.8457454632 noise=0
Ga353 ns353 0 ns354 0 -1.57343392648
Ga354 ns354 0 ns353 0 1.57343392648
Ca355 ns355 0 1e-12
Ca356 ns356 0 1e-12
Ra355 ns355 0 27.1849571621 noise=0
Ra356 ns356 0 27.1849571621 noise=0
Ga355 ns355 0 ns356 0 -1.49976985502
Ga356 ns356 0 ns355 0 1.49976985502
Ca357 ns357 0 1e-12
Ca358 ns358 0 1e-12
Ra357 ns357 0 294.868225966 noise=0
Ra358 ns358 0 294.868225966 noise=0
Ga357 ns357 0 ns358 0 -1.43272297288
Ga358 ns358 0 ns357 0 1.43272297288
Ca359 ns359 0 1e-12
Ca360 ns360 0 1e-12
Ra359 ns359 0 24.065722504 noise=0
Ra360 ns360 0 24.065722504 noise=0
Ga359 ns359 0 ns360 0 -1.39531521009
Ga360 ns360 0 ns359 0 1.39531521009
Ca361 ns361 0 1e-12
Ca362 ns362 0 1e-12
Ra361 ns361 0 27.949811121 noise=0
Ra362 ns362 0 27.949811121 noise=0
Ga361 ns361 0 ns362 0 -1.32076031205
Ga362 ns362 0 ns361 0 1.32076031205
Ca363 ns363 0 1e-12
Ca364 ns364 0 1e-12
Ra363 ns363 0 68.9019895791 noise=0
Ra364 ns364 0 68.9019895791 noise=0
Ga363 ns363 0 ns364 0 -1.26735586041
Ga364 ns364 0 ns363 0 1.26735586041
Ca365 ns365 0 1e-12
Ca366 ns366 0 1e-12
Ra365 ns365 0 17.4920890166 noise=0
Ra366 ns366 0 17.4920890166 noise=0
Ga365 ns365 0 ns366 0 -1.21455822137
Ga366 ns366 0 ns365 0 1.21455822137
Ca367 ns367 0 1e-12
Ca368 ns368 0 1e-12
Ra367 ns367 0 23.7303485873 noise=0
Ra368 ns368 0 23.7303485873 noise=0
Ga367 ns367 0 ns368 0 -1.13110590561
Ga368 ns368 0 ns367 0 1.13110590561
Ca369 ns369 0 1e-12
Ca370 ns370 0 1e-12
Ra369 ns369 0 12.6702453574 noise=0
Ra370 ns370 0 12.6702453574 noise=0
Ga369 ns369 0 ns370 0 -1.01544529945
Ga370 ns370 0 ns369 0 1.01544529945
Ca371 ns371 0 1e-12
Ca372 ns372 0 1e-12
Ra371 ns371 0 22.4497679254 noise=0
Ra372 ns372 0 22.4497679254 noise=0
Ga371 ns371 0 ns372 0 -0.947337481808
Ga372 ns372 0 ns371 0 0.947337481808
Ca373 ns373 0 1e-12
Ca374 ns374 0 1e-12
Ra373 ns373 0 19.3969089633 noise=0
Ra374 ns374 0 19.3969089633 noise=0
Ga373 ns373 0 ns374 0 -0.828769989963
Ga374 ns374 0 ns373 0 0.828769989963
Ca375 ns375 0 1e-12
Ca376 ns376 0 1e-12
Ra375 ns375 0 28.1931334636 noise=0
Ra376 ns376 0 28.1931334636 noise=0
Ga375 ns375 0 ns376 0 -0.753040704424
Ga376 ns376 0 ns375 0 0.753040704424
Ca377 ns377 0 1e-12
Ca378 ns378 0 1e-12
Ra377 ns377 0 9.58447239365 noise=0
Ra378 ns378 0 9.58447239365 noise=0
Ga377 ns377 0 ns378 0 -0.706025240203
Ga378 ns378 0 ns377 0 0.706025240203
Ca379 ns379 0 1e-12
Ca380 ns380 0 1e-12
Ra379 ns379 0 19.2217606518 noise=0
Ra380 ns380 0 19.2217606518 noise=0
Ga379 ns379 0 ns380 0 -0.584920288579
Ga380 ns380 0 ns379 0 0.584920288579
Ca381 ns381 0 1e-12
Ca382 ns382 0 1e-12
Ra381 ns381 0 12.9186134131 noise=0
Ra382 ns382 0 12.9186134131 noise=0
Ga381 ns381 0 ns382 0 -0.451995255731
Ga382 ns382 0 ns381 0 0.451995255731
Ca383 ns383 0 1e-12
Ca384 ns384 0 1e-12
Ra383 ns383 0 14.6643586754 noise=0
Ra384 ns384 0 14.6643586754 noise=0
Ga383 ns383 0 ns384 0 -0.39239765994
Ga384 ns384 0 ns383 0 0.39239765994
Ca385 ns385 0 1e-12
Ca386 ns386 0 1e-12
Ra385 ns385 0 18.5528384969 noise=0
Ra386 ns386 0 18.5528384969 noise=0
Ga385 ns385 0 ns386 0 -0.213309922964
Ga386 ns386 0 ns385 0 0.213309922964
Ca387 ns387 0 1e-12
Ca388 ns388 0 1e-12
Ra387 ns387 0 16.425306589 noise=0
Ra388 ns388 0 16.425306589 noise=0
Ga387 ns387 0 ns388 0 -0.132506240506
Ga388 ns388 0 ns387 0 0.132506240506
Ca389 ns389 0 1e-12
Ra389 ns389 0 12.9927381247 noise=0
Ca390 ns390 0 1e-12
Ra390 ns390 0 99.3047026559 noise=0
Ca391 ns391 0 1e-12
Ca392 ns392 0 1e-12
Ra391 ns391 0 116.054358759 noise=0
Ra392 ns392 0 116.054358759 noise=0
Ga391 ns391 0 ns392 0 -0.0790828435996
Ga392 ns392 0 ns391 0 0.0790828435996
Ca393 ns393 0 1e-12
Ca394 ns394 0 1e-12
Ra393 ns393 0 0.177524466588 noise=0
Ra394 ns394 0 0.177524466588 noise=0
Ga393 ns393 0 ns394 0 -0.592192182122
Ga394 ns394 0 ns393 0 0.592192182122
Ca395 ns395 0 1e-12
Ca396 ns396 0 1e-12
Ra395 ns395 0 3.73043526058 noise=0
Ra396 ns396 0 3.73043526058 noise=0
Ga395 ns395 0 ns396 0 -1.88816876812
Ga396 ns396 0 ns395 0 1.88816876812
Ca397 ns397 0 1e-12
Ca398 ns398 0 1e-12
Ra397 ns397 0 78.3630472463 noise=0
Ra398 ns398 0 78.3630472463 noise=0
Ga397 ns397 0 ns398 0 -1.87552614083
Ga398 ns398 0 ns397 0 1.87552614083
Ca399 ns399 0 1e-12
Ca400 ns400 0 1e-12
Ra399 ns399 0 28.6294222129 noise=0
Ra400 ns400 0 28.6294222129 noise=0
Ga399 ns399 0 ns400 0 -1.8615708713
Ga400 ns400 0 ns399 0 1.8615708713
Ca401 ns401 0 1e-12
Ca402 ns402 0 1e-12
Ra401 ns401 0 934.131832031 noise=0
Ra402 ns402 0 934.131832031 noise=0
Ga401 ns401 0 ns402 0 -1.77206208419
Ga402 ns402 0 ns401 0 1.77206208419
Ca403 ns403 0 1e-12
Ca404 ns404 0 1e-12
Ra403 ns403 0 30.3138883767 noise=0
Ra404 ns404 0 30.3138883767 noise=0
Ga403 ns403 0 ns404 0 -1.74835043081
Ga404 ns404 0 ns403 0 1.74835043081
Ca405 ns405 0 1e-12
Ca406 ns406 0 1e-12
Ra405 ns405 0 29.0014618309 noise=0
Ra406 ns406 0 29.0014618309 noise=0
Ga405 ns405 0 ns406 0 -1.68453524434
Ga406 ns406 0 ns405 0 1.68453524434
Ca407 ns407 0 1e-12
Ca408 ns408 0 1e-12
Ra407 ns407 0 608.740499085 noise=0
Ra408 ns408 0 608.740499085 noise=0
Ga407 ns407 0 ns408 0 -1.60136974681
Ga408 ns408 0 ns407 0 1.60136974681
Ca409 ns409 0 1e-12
Ca410 ns410 0 1e-12
Ra409 ns409 0 28.8457454632 noise=0
Ra410 ns410 0 28.8457454632 noise=0
Ga409 ns409 0 ns410 0 -1.57343392648
Ga410 ns410 0 ns409 0 1.57343392648
Ca411 ns411 0 1e-12
Ca412 ns412 0 1e-12
Ra411 ns411 0 27.1849571621 noise=0
Ra412 ns412 0 27.1849571621 noise=0
Ga411 ns411 0 ns412 0 -1.49976985502
Ga412 ns412 0 ns411 0 1.49976985502
Ca413 ns413 0 1e-12
Ca414 ns414 0 1e-12
Ra413 ns413 0 294.868225966 noise=0
Ra414 ns414 0 294.868225966 noise=0
Ga413 ns413 0 ns414 0 -1.43272297288
Ga414 ns414 0 ns413 0 1.43272297288
Ca415 ns415 0 1e-12
Ca416 ns416 0 1e-12
Ra415 ns415 0 24.065722504 noise=0
Ra416 ns416 0 24.065722504 noise=0
Ga415 ns415 0 ns416 0 -1.39531521009
Ga416 ns416 0 ns415 0 1.39531521009
Ca417 ns417 0 1e-12
Ca418 ns418 0 1e-12
Ra417 ns417 0 27.949811121 noise=0
Ra418 ns418 0 27.949811121 noise=0
Ga417 ns417 0 ns418 0 -1.32076031205
Ga418 ns418 0 ns417 0 1.32076031205
Ca419 ns419 0 1e-12
Ca420 ns420 0 1e-12
Ra419 ns419 0 68.9019895791 noise=0
Ra420 ns420 0 68.9019895791 noise=0
Ga419 ns419 0 ns420 0 -1.26735586041
Ga420 ns420 0 ns419 0 1.26735586041
Ca421 ns421 0 1e-12
Ca422 ns422 0 1e-12
Ra421 ns421 0 17.4920890166 noise=0
Ra422 ns422 0 17.4920890166 noise=0
Ga421 ns421 0 ns422 0 -1.21455822137
Ga422 ns422 0 ns421 0 1.21455822137
Ca423 ns423 0 1e-12
Ca424 ns424 0 1e-12
Ra423 ns423 0 23.7303485873 noise=0
Ra424 ns424 0 23.7303485873 noise=0
Ga423 ns423 0 ns424 0 -1.13110590561
Ga424 ns424 0 ns423 0 1.13110590561
Ca425 ns425 0 1e-12
Ca426 ns426 0 1e-12
Ra425 ns425 0 12.6702453574 noise=0
Ra426 ns426 0 12.6702453574 noise=0
Ga425 ns425 0 ns426 0 -1.01544529945
Ga426 ns426 0 ns425 0 1.01544529945
Ca427 ns427 0 1e-12
Ca428 ns428 0 1e-12
Ra427 ns427 0 22.4497679254 noise=0
Ra428 ns428 0 22.4497679254 noise=0
Ga427 ns427 0 ns428 0 -0.947337481808
Ga428 ns428 0 ns427 0 0.947337481808
Ca429 ns429 0 1e-12
Ca430 ns430 0 1e-12
Ra429 ns429 0 19.3969089633 noise=0
Ra430 ns430 0 19.3969089633 noise=0
Ga429 ns429 0 ns430 0 -0.828769989963
Ga430 ns430 0 ns429 0 0.828769989963
Ca431 ns431 0 1e-12
Ca432 ns432 0 1e-12
Ra431 ns431 0 28.1931334636 noise=0
Ra432 ns432 0 28.1931334636 noise=0
Ga431 ns431 0 ns432 0 -0.753040704424
Ga432 ns432 0 ns431 0 0.753040704424
Ca433 ns433 0 1e-12
Ca434 ns434 0 1e-12
Ra433 ns433 0 9.58447239365 noise=0
Ra434 ns434 0 9.58447239365 noise=0
Ga433 ns433 0 ns434 0 -0.706025240203
Ga434 ns434 0 ns433 0 0.706025240203
Ca435 ns435 0 1e-12
Ca436 ns436 0 1e-12
Ra435 ns435 0 19.2217606518 noise=0
Ra436 ns436 0 19.2217606518 noise=0
Ga435 ns435 0 ns436 0 -0.584920288579
Ga436 ns436 0 ns435 0 0.584920288579
Ca437 ns437 0 1e-12
Ca438 ns438 0 1e-12
Ra437 ns437 0 12.9186134131 noise=0
Ra438 ns438 0 12.9186134131 noise=0
Ga437 ns437 0 ns438 0 -0.451995255731
Ga438 ns438 0 ns437 0 0.451995255731
Ca439 ns439 0 1e-12
Ca440 ns440 0 1e-12
Ra439 ns439 0 14.6643586754 noise=0
Ra440 ns440 0 14.6643586754 noise=0
Ga439 ns439 0 ns440 0 -0.39239765994
Ga440 ns440 0 ns439 0 0.39239765994
Ca441 ns441 0 1e-12
Ca442 ns442 0 1e-12
Ra441 ns441 0 18.5528384969 noise=0
Ra442 ns442 0 18.5528384969 noise=0
Ga441 ns441 0 ns442 0 -0.213309922964
Ga442 ns442 0 ns441 0 0.213309922964
Ca443 ns443 0 1e-12
Ca444 ns444 0 1e-12
Ra443 ns443 0 16.425306589 noise=0
Ra444 ns444 0 16.425306589 noise=0
Ga443 ns443 0 ns444 0 -0.132506240506
Ga444 ns444 0 ns443 0 0.132506240506
Ca445 ns445 0 1e-12
Ra445 ns445 0 12.9927381247 noise=0
Ca446 ns446 0 1e-12
Ra446 ns446 0 99.3047026559 noise=0
Ca447 ns447 0 1e-12
Ca448 ns448 0 1e-12
Ra447 ns447 0 116.054358759 noise=0
Ra448 ns448 0 116.054358759 noise=0
Ga447 ns447 0 ns448 0 -0.0790828435996
Ga448 ns448 0 ns447 0 0.0790828435996

Gb1_1 ns1 0 ni1 0 -0.242230162508
Gb2_1 ns2 0 ni1 0 -5.66981737855
Gb3_1 ns3 0 ni1 0 1.70052379695
Gb4_1 ns4 0 ni1 0 1.58977849418
Gb5_1 ns5 0 ni1 0 1.86936465941
Gb6_1 ns6 0 ni1 0 0.918326016818
Gb7_1 ns7 0 ni1 0 1.86091951073
Gb8_1 ns8 0 ni1 0 -0.0696438180465
Gb9_1 ns9 0 ni1 0 1.7715070455
Gb10_1 ns10 0 ni1 0 0.919848034492
Gb11_1 ns11 0 ni1 0 -0.760413119527
Gb12_1 ns12 0 ni1 0 -1.73462525062
Gb13_1 ns13 0 ni1 0 1.66554798658
Gb14_1 ns14 0 ni1 0 -0.962084218547
Gb15_1 ns15 0 ni1 0 0.881978685923
Gb16_1 ns16 0 ni1 0 1.60046667014
Gb17_1 ns17 0 ni1 0 -1.55772849734
Gb18_1 ns18 0 ni1 0 0.747487499417
Gb19_1 ns19 0 ni1 0 -1.15723265214
Gb20_1 ns20 0 ni1 0 -1.4722884914
Gb21_1 ns21 0 ni1 0 -1.43065334637
Gb22_1 ns22 0 ni1 0 0.877735034392
Gb23_1 ns23 0 ni1 0 -0.0366302966022
Gb24_1 ns24 0 ni1 0 -1.3954618059
Gb25_1 ns25 0 ni1 0 1.30856229812
Gb26_1 ns26 0 ni1 0 0.486068116494
Gb27_1 ns27 0 ni1 0 -1.08772879245
Gb28_1 ns28 0 ni1 0 1.2550657279
Gb29_1 ns29 0 ni1 0 0.406136520382
Gb30_1 ns30 0 ni1 0 1.19813246552
Gb31_1 ns31 0 ni1 0 1.09813888731
Gb32_1 ns32 0 ni1 0 -0.927025586813
Gb33_1 ns33 0 ni1 0 -0.772633145912
Gb34_1 ns34 0 ni1 0 0.961527123453
Gb35_1 ns35 0 ni1 0 -0.623541296567
Gb36_1 ns36 0 ni1 0 0.920112973699
Gb37_1 ns37 0 ni1 0 -0.197470289704
Gb38_1 ns38 0 ni1 0 0.819693134289
Gb39_1 ns39 0 ni1 0 -0.752268145323
Gb40_1 ns40 0 ni1 0 -0.0518715051145
Gb41_1 ns41 0 ni1 0 -0.181587927011
Gb42_1 ns42 0 ni1 0 0.694608973231
Gb43_1 ns43 0 ni1 0 0.169134997258
Gb44_1 ns44 0 ni1 0 -0.574504157078
Gb45_1 ns45 0 ni1 0 -0.423994579197
Gb46_1 ns46 0 ni1 0 -0.24090789391
Gb47_1 ns47 0 ni1 0 0.374937946713
Gb48_1 ns48 0 ni1 0 -0.168660279104
Gb49_1 ns49 0 ni1 0 -0.0301538467221
Gb50_1 ns50 0 ni1 0 0.219310234788
Gb51_1 ns51 0 ni1 0 -0.12047842402
Gb52_1 ns52 0 ni1 0 0.0870596730425
Gb53_1 ns53 0 ni1 0 -0.076966070616
Gb54_1 ns54 0 ni1 0 -0.0100700165577
Gb55_1 ns55 0 ni1 0 0.0781839687698
Gb56_1 ns56 0 ni1 0 -0.016866442929
Gb57_2 ns57 0 ni2 0 -0.242230162508
Gb58_2 ns58 0 ni2 0 -5.66981737855
Gb59_2 ns59 0 ni2 0 1.70052379695
Gb60_2 ns60 0 ni2 0 1.58977849418
Gb61_2 ns61 0 ni2 0 1.86936465941
Gb62_2 ns62 0 ni2 0 0.918326016818
Gb63_2 ns63 0 ni2 0 1.86091951073
Gb64_2 ns64 0 ni2 0 -0.0696438180465
Gb65_2 ns65 0 ni2 0 1.7715070455
Gb66_2 ns66 0 ni2 0 0.919848034492
Gb67_2 ns67 0 ni2 0 -0.760413119527
Gb68_2 ns68 0 ni2 0 -1.73462525062
Gb69_2 ns69 0 ni2 0 1.66554798658
Gb70_2 ns70 0 ni2 0 -0.962084218547
Gb71_2 ns71 0 ni2 0 0.881978685923
Gb72_2 ns72 0 ni2 0 1.60046667014
Gb73_2 ns73 0 ni2 0 -1.55772849734
Gb74_2 ns74 0 ni2 0 0.747487499417
Gb75_2 ns75 0 ni2 0 -1.15723265214
Gb76_2 ns76 0 ni2 0 -1.4722884914
Gb77_2 ns77 0 ni2 0 -1.43065334637
Gb78_2 ns78 0 ni2 0 0.877735034392
Gb79_2 ns79 0 ni2 0 -0.0366302966022
Gb80_2 ns80 0 ni2 0 -1.3954618059
Gb81_2 ns81 0 ni2 0 1.30856229812
Gb82_2 ns82 0 ni2 0 0.486068116494
Gb83_2 ns83 0 ni2 0 -1.08772879245
Gb84_2 ns84 0 ni2 0 1.2550657279
Gb85_2 ns85 0 ni2 0 0.406136520382
Gb86_2 ns86 0 ni2 0 1.19813246552
Gb87_2 ns87 0 ni2 0 1.09813888731
Gb88_2 ns88 0 ni2 0 -0.927025586813
Gb89_2 ns89 0 ni2 0 -0.772633145912
Gb90_2 ns90 0 ni2 0 0.961527123453
Gb91_2 ns91 0 ni2 0 -0.623541296567
Gb92_2 ns92 0 ni2 0 0.920112973699
Gb93_2 ns93 0 ni2 0 -0.197470289704
Gb94_2 ns94 0 ni2 0 0.819693134289
Gb95_2 ns95 0 ni2 0 -0.752268145323
Gb96_2 ns96 0 ni2 0 -0.0518715051145
Gb97_2 ns97 0 ni2 0 -0.181587927011
Gb98_2 ns98 0 ni2 0 0.694608973231
Gb99_2 ns99 0 ni2 0 0.169134997258
Gb100_2 ns100 0 ni2 0 -0.574504157078
Gb101_2 ns101 0 ni2 0 -0.423994579197
Gb102_2 ns102 0 ni2 0 -0.24090789391
Gb103_2 ns103 0 ni2 0 0.374937946713
Gb104_2 ns104 0 ni2 0 -0.168660279104
Gb105_2 ns105 0 ni2 0 -0.0301538467221
Gb106_2 ns106 0 ni2 0 0.219310234788
Gb107_2 ns107 0 ni2 0 -0.12047842402
Gb108_2 ns108 0 ni2 0 0.0870596730425
Gb109_2 ns109 0 ni2 0 -0.076966070616
Gb110_2 ns110 0 ni2 0 -0.0100700165577
Gb111_2 ns111 0 ni2 0 0.0781839687698
Gb112_2 ns112 0 ni2 0 -0.016866442929
Gb113_3 ns113 0 ni3 0 -0.242230162508
Gb114_3 ns114 0 ni3 0 -5.66981737855
Gb115_3 ns115 0 ni3 0 1.70052379695
Gb116_3 ns116 0 ni3 0 1.58977849418
Gb117_3 ns117 0 ni3 0 1.86936465941
Gb118_3 ns118 0 ni3 0 0.918326016818
Gb119_3 ns119 0 ni3 0 1.86091951073
Gb120_3 ns120 0 ni3 0 -0.0696438180465
Gb121_3 ns121 0 ni3 0 1.7715070455
Gb122_3 ns122 0 ni3 0 0.919848034492
Gb123_3 ns123 0 ni3 0 -0.760413119527
Gb124_3 ns124 0 ni3 0 -1.73462525062
Gb125_3 ns125 0 ni3 0 1.66554798658
Gb126_3 ns126 0 ni3 0 -0.962084218547
Gb127_3 ns127 0 ni3 0 0.881978685923
Gb128_3 ns128 0 ni3 0 1.60046667014
Gb129_3 ns129 0 ni3 0 -1.55772849734
Gb130_3 ns130 0 ni3 0 0.747487499417
Gb131_3 ns131 0 ni3 0 -1.15723265214
Gb132_3 ns132 0 ni3 0 -1.4722884914
Gb133_3 ns133 0 ni3 0 -1.43065334637
Gb134_3 ns134 0 ni3 0 0.877735034392
Gb135_3 ns135 0 ni3 0 -0.0366302966022
Gb136_3 ns136 0 ni3 0 -1.3954618059
Gb137_3 ns137 0 ni3 0 1.30856229812
Gb138_3 ns138 0 ni3 0 0.486068116494
Gb139_3 ns139 0 ni3 0 -1.08772879245
Gb140_3 ns140 0 ni3 0 1.2550657279
Gb141_3 ns141 0 ni3 0 0.406136520382
Gb142_3 ns142 0 ni3 0 1.19813246552
Gb143_3 ns143 0 ni3 0 1.09813888731
Gb144_3 ns144 0 ni3 0 -0.927025586813
Gb145_3 ns145 0 ni3 0 -0.772633145912
Gb146_3 ns146 0 ni3 0 0.961527123453
Gb147_3 ns147 0 ni3 0 -0.623541296567
Gb148_3 ns148 0 ni3 0 0.920112973699
Gb149_3 ns149 0 ni3 0 -0.197470289704
Gb150_3 ns150 0 ni3 0 0.819693134289
Gb151_3 ns151 0 ni3 0 -0.752268145323
Gb152_3 ns152 0 ni3 0 -0.0518715051145
Gb153_3 ns153 0 ni3 0 -0.181587927011
Gb154_3 ns154 0 ni3 0 0.694608973231
Gb155_3 ns155 0 ni3 0 0.169134997258
Gb156_3 ns156 0 ni3 0 -0.574504157078
Gb157_3 ns157 0 ni3 0 -0.423994579197
Gb158_3 ns158 0 ni3 0 -0.24090789391
Gb159_3 ns159 0 ni3 0 0.374937946713
Gb160_3 ns160 0 ni3 0 -0.168660279104
Gb161_3 ns161 0 ni3 0 -0.0301538467221
Gb162_3 ns162 0 ni3 0 0.219310234788
Gb163_3 ns163 0 ni3 0 -0.12047842402
Gb164_3 ns164 0 ni3 0 0.0870596730425
Gb165_3 ns165 0 ni3 0 -0.076966070616
Gb166_3 ns166 0 ni3 0 -0.0100700165577
Gb167_3 ns167 0 ni3 0 0.0781839687698
Gb168_3 ns168 0 ni3 0 -0.016866442929
Gb169_4 ns169 0 ni4 0 -0.242230162508
Gb170_4 ns170 0 ni4 0 -5.66981737855
Gb171_4 ns171 0 ni4 0 1.70052379695
Gb172_4 ns172 0 ni4 0 1.58977849418
Gb173_4 ns173 0 ni4 0 1.86936465941
Gb174_4 ns174 0 ni4 0 0.918326016818
Gb175_4 ns175 0 ni4 0 1.86091951073
Gb176_4 ns176 0 ni4 0 -0.0696438180465
Gb177_4 ns177 0 ni4 0 1.7715070455
Gb178_4 ns178 0 ni4 0 0.919848034492
Gb179_4 ns179 0 ni4 0 -0.760413119527
Gb180_4 ns180 0 ni4 0 -1.73462525062
Gb181_4 ns181 0 ni4 0 1.66554798658
Gb182_4 ns182 0 ni4 0 -0.962084218547
Gb183_4 ns183 0 ni4 0 0.881978685923
Gb184_4 ns184 0 ni4 0 1.60046667014
Gb185_4 ns185 0 ni4 0 -1.55772849734
Gb186_4 ns186 0 ni4 0 0.747487499417
Gb187_4 ns187 0 ni4 0 -1.15723265214
Gb188_4 ns188 0 ni4 0 -1.4722884914
Gb189_4 ns189 0 ni4 0 -1.43065334637
Gb190_4 ns190 0 ni4 0 0.877735034392
Gb191_4 ns191 0 ni4 0 -0.0366302966022
Gb192_4 ns192 0 ni4 0 -1.3954618059
Gb193_4 ns193 0 ni4 0 1.30856229812
Gb194_4 ns194 0 ni4 0 0.486068116494
Gb195_4 ns195 0 ni4 0 -1.08772879245
Gb196_4 ns196 0 ni4 0 1.2550657279
Gb197_4 ns197 0 ni4 0 0.406136520382
Gb198_4 ns198 0 ni4 0 1.19813246552
Gb199_4 ns199 0 ni4 0 1.09813888731
Gb200_4 ns200 0 ni4 0 -0.927025586813
Gb201_4 ns201 0 ni4 0 -0.772633145912
Gb202_4 ns202 0 ni4 0 0.961527123453
Gb203_4 ns203 0 ni4 0 -0.623541296567
Gb204_4 ns204 0 ni4 0 0.920112973699
Gb205_4 ns205 0 ni4 0 -0.197470289704
Gb206_4 ns206 0 ni4 0 0.819693134289
Gb207_4 ns207 0 ni4 0 -0.752268145323
Gb208_4 ns208 0 ni4 0 -0.0518715051145
Gb209_4 ns209 0 ni4 0 -0.181587927011
Gb210_4 ns210 0 ni4 0 0.694608973231
Gb211_4 ns211 0 ni4 0 0.169134997258
Gb212_4 ns212 0 ni4 0 -0.574504157078
Gb213_4 ns213 0 ni4 0 -0.423994579197
Gb214_4 ns214 0 ni4 0 -0.24090789391
Gb215_4 ns215 0 ni4 0 0.374937946713
Gb216_4 ns216 0 ni4 0 -0.168660279104
Gb217_4 ns217 0 ni4 0 -0.0301538467221
Gb218_4 ns218 0 ni4 0 0.219310234788
Gb219_4 ns219 0 ni4 0 -0.12047842402
Gb220_4 ns220 0 ni4 0 0.0870596730425
Gb221_4 ns221 0 ni4 0 -0.076966070616
Gb222_4 ns222 0 ni4 0 -0.0100700165577
Gb223_4 ns223 0 ni4 0 0.0781839687698
Gb224_4 ns224 0 ni4 0 -0.016866442929
Gb225_5 ns225 0 ni5 0 -0.242230162508
Gb226_5 ns226 0 ni5 0 -5.66981737855
Gb227_5 ns227 0 ni5 0 1.70052379695
Gb228_5 ns228 0 ni5 0 1.58977849418
Gb229_5 ns229 0 ni5 0 1.86936465941
Gb230_5 ns230 0 ni5 0 0.918326016818
Gb231_5 ns231 0 ni5 0 1.86091951073
Gb232_5 ns232 0 ni5 0 -0.0696438180465
Gb233_5 ns233 0 ni5 0 1.7715070455
Gb234_5 ns234 0 ni5 0 0.919848034492
Gb235_5 ns235 0 ni5 0 -0.760413119527
Gb236_5 ns236 0 ni5 0 -1.73462525062
Gb237_5 ns237 0 ni5 0 1.66554798658
Gb238_5 ns238 0 ni5 0 -0.962084218547
Gb239_5 ns239 0 ni5 0 0.881978685923
Gb240_5 ns240 0 ni5 0 1.60046667014
Gb241_5 ns241 0 ni5 0 -1.55772849734
Gb242_5 ns242 0 ni5 0 0.747487499417
Gb243_5 ns243 0 ni5 0 -1.15723265214
Gb244_5 ns244 0 ni5 0 -1.4722884914
Gb245_5 ns245 0 ni5 0 -1.43065334637
Gb246_5 ns246 0 ni5 0 0.877735034392
Gb247_5 ns247 0 ni5 0 -0.0366302966022
Gb248_5 ns248 0 ni5 0 -1.3954618059
Gb249_5 ns249 0 ni5 0 1.30856229812
Gb250_5 ns250 0 ni5 0 0.486068116494
Gb251_5 ns251 0 ni5 0 -1.08772879245
Gb252_5 ns252 0 ni5 0 1.2550657279
Gb253_5 ns253 0 ni5 0 0.406136520382
Gb254_5 ns254 0 ni5 0 1.19813246552
Gb255_5 ns255 0 ni5 0 1.09813888731
Gb256_5 ns256 0 ni5 0 -0.927025586813
Gb257_5 ns257 0 ni5 0 -0.772633145912
Gb258_5 ns258 0 ni5 0 0.961527123453
Gb259_5 ns259 0 ni5 0 -0.623541296567
Gb260_5 ns260 0 ni5 0 0.920112973699
Gb261_5 ns261 0 ni5 0 -0.197470289704
Gb262_5 ns262 0 ni5 0 0.819693134289
Gb263_5 ns263 0 ni5 0 -0.752268145323
Gb264_5 ns264 0 ni5 0 -0.0518715051145
Gb265_5 ns265 0 ni5 0 -0.181587927011
Gb266_5 ns266 0 ni5 0 0.694608973231
Gb267_5 ns267 0 ni5 0 0.169134997258
Gb268_5 ns268 0 ni5 0 -0.574504157078
Gb269_5 ns269 0 ni5 0 -0.423994579197
Gb270_5 ns270 0 ni5 0 -0.24090789391
Gb271_5 ns271 0 ni5 0 0.374937946713
Gb272_5 ns272 0 ni5 0 -0.168660279104
Gb273_5 ns273 0 ni5 0 -0.0301538467221
Gb274_5 ns274 0 ni5 0 0.219310234788
Gb275_5 ns275 0 ni5 0 -0.12047842402
Gb276_5 ns276 0 ni5 0 0.0870596730425
Gb277_5 ns277 0 ni5 0 -0.076966070616
Gb278_5 ns278 0 ni5 0 -0.0100700165577
Gb279_5 ns279 0 ni5 0 0.0781839687698
Gb280_5 ns280 0 ni5 0 -0.016866442929
Gb281_6 ns281 0 ni6 0 -0.242230162508
Gb282_6 ns282 0 ni6 0 -5.66981737855
Gb283_6 ns283 0 ni6 0 1.70052379695
Gb284_6 ns284 0 ni6 0 1.58977849418
Gb285_6 ns285 0 ni6 0 1.86936465941
Gb286_6 ns286 0 ni6 0 0.918326016818
Gb287_6 ns287 0 ni6 0 1.86091951073
Gb288_6 ns288 0 ni6 0 -0.0696438180465
Gb289_6 ns289 0 ni6 0 1.7715070455
Gb290_6 ns290 0 ni6 0 0.919848034492
Gb291_6 ns291 0 ni6 0 -0.760413119527
Gb292_6 ns292 0 ni6 0 -1.73462525062
Gb293_6 ns293 0 ni6 0 1.66554798658
Gb294_6 ns294 0 ni6 0 -0.962084218547
Gb295_6 ns295 0 ni6 0 0.881978685923
Gb296_6 ns296 0 ni6 0 1.60046667014
Gb297_6 ns297 0 ni6 0 -1.55772849734
Gb298_6 ns298 0 ni6 0 0.747487499417
Gb299_6 ns299 0 ni6 0 -1.15723265214
Gb300_6 ns300 0 ni6 0 -1.4722884914
Gb301_6 ns301 0 ni6 0 -1.43065334637
Gb302_6 ns302 0 ni6 0 0.877735034392
Gb303_6 ns303 0 ni6 0 -0.0366302966022
Gb304_6 ns304 0 ni6 0 -1.3954618059
Gb305_6 ns305 0 ni6 0 1.30856229812
Gb306_6 ns306 0 ni6 0 0.486068116494
Gb307_6 ns307 0 ni6 0 -1.08772879245
Gb308_6 ns308 0 ni6 0 1.2550657279
Gb309_6 ns309 0 ni6 0 0.406136520382
Gb310_6 ns310 0 ni6 0 1.19813246552
Gb311_6 ns311 0 ni6 0 1.09813888731
Gb312_6 ns312 0 ni6 0 -0.927025586813
Gb313_6 ns313 0 ni6 0 -0.772633145912
Gb314_6 ns314 0 ni6 0 0.961527123453
Gb315_6 ns315 0 ni6 0 -0.623541296567
Gb316_6 ns316 0 ni6 0 0.920112973699
Gb317_6 ns317 0 ni6 0 -0.197470289704
Gb318_6 ns318 0 ni6 0 0.819693134289
Gb319_6 ns319 0 ni6 0 -0.752268145323
Gb320_6 ns320 0 ni6 0 -0.0518715051145
Gb321_6 ns321 0 ni6 0 -0.181587927011
Gb322_6 ns322 0 ni6 0 0.694608973231
Gb323_6 ns323 0 ni6 0 0.169134997258
Gb324_6 ns324 0 ni6 0 -0.574504157078
Gb325_6 ns325 0 ni6 0 -0.423994579197
Gb326_6 ns326 0 ni6 0 -0.24090789391
Gb327_6 ns327 0 ni6 0 0.374937946713
Gb328_6 ns328 0 ni6 0 -0.168660279104
Gb329_6 ns329 0 ni6 0 -0.0301538467221
Gb330_6 ns330 0 ni6 0 0.219310234788
Gb331_6 ns331 0 ni6 0 -0.12047842402
Gb332_6 ns332 0 ni6 0 0.0870596730425
Gb333_6 ns333 0 ni6 0 -0.076966070616
Gb334_6 ns334 0 ni6 0 -0.0100700165577
Gb335_6 ns335 0 ni6 0 0.0781839687698
Gb336_6 ns336 0 ni6 0 -0.016866442929
Gb337_7 ns337 0 ni7 0 -0.242230162508
Gb338_7 ns338 0 ni7 0 -5.66981737855
Gb339_7 ns339 0 ni7 0 1.70052379695
Gb340_7 ns340 0 ni7 0 1.58977849418
Gb341_7 ns341 0 ni7 0 1.86936465941
Gb342_7 ns342 0 ni7 0 0.918326016818
Gb343_7 ns343 0 ni7 0 1.86091951073
Gb344_7 ns344 0 ni7 0 -0.0696438180465
Gb345_7 ns345 0 ni7 0 1.7715070455
Gb346_7 ns346 0 ni7 0 0.919848034492
Gb347_7 ns347 0 ni7 0 -0.760413119527
Gb348_7 ns348 0 ni7 0 -1.73462525062
Gb349_7 ns349 0 ni7 0 1.66554798658
Gb350_7 ns350 0 ni7 0 -0.962084218547
Gb351_7 ns351 0 ni7 0 0.881978685923
Gb352_7 ns352 0 ni7 0 1.60046667014
Gb353_7 ns353 0 ni7 0 -1.55772849734
Gb354_7 ns354 0 ni7 0 0.747487499417
Gb355_7 ns355 0 ni7 0 -1.15723265214
Gb356_7 ns356 0 ni7 0 -1.4722884914
Gb357_7 ns357 0 ni7 0 -1.43065334637
Gb358_7 ns358 0 ni7 0 0.877735034392
Gb359_7 ns359 0 ni7 0 -0.0366302966022
Gb360_7 ns360 0 ni7 0 -1.3954618059
Gb361_7 ns361 0 ni7 0 1.30856229812
Gb362_7 ns362 0 ni7 0 0.486068116494
Gb363_7 ns363 0 ni7 0 -1.08772879245
Gb364_7 ns364 0 ni7 0 1.2550657279
Gb365_7 ns365 0 ni7 0 0.406136520382
Gb366_7 ns366 0 ni7 0 1.19813246552
Gb367_7 ns367 0 ni7 0 1.09813888731
Gb368_7 ns368 0 ni7 0 -0.927025586813
Gb369_7 ns369 0 ni7 0 -0.772633145912
Gb370_7 ns370 0 ni7 0 0.961527123453
Gb371_7 ns371 0 ni7 0 -0.623541296567
Gb372_7 ns372 0 ni7 0 0.920112973699
Gb373_7 ns373 0 ni7 0 -0.197470289704
Gb374_7 ns374 0 ni7 0 0.819693134289
Gb375_7 ns375 0 ni7 0 -0.752268145323
Gb376_7 ns376 0 ni7 0 -0.0518715051145
Gb377_7 ns377 0 ni7 0 -0.181587927011
Gb378_7 ns378 0 ni7 0 0.694608973231
Gb379_7 ns379 0 ni7 0 0.169134997258
Gb380_7 ns380 0 ni7 0 -0.574504157078
Gb381_7 ns381 0 ni7 0 -0.423994579197
Gb382_7 ns382 0 ni7 0 -0.24090789391
Gb383_7 ns383 0 ni7 0 0.374937946713
Gb384_7 ns384 0 ni7 0 -0.168660279104
Gb385_7 ns385 0 ni7 0 -0.0301538467221
Gb386_7 ns386 0 ni7 0 0.219310234788
Gb387_7 ns387 0 ni7 0 -0.12047842402
Gb388_7 ns388 0 ni7 0 0.0870596730425
Gb389_7 ns389 0 ni7 0 -0.076966070616
Gb390_7 ns390 0 ni7 0 -0.0100700165577
Gb391_7 ns391 0 ni7 0 0.0781839687698
Gb392_7 ns392 0 ni7 0 -0.016866442929
Gb393_8 ns393 0 ni8 0 -0.242230162508
Gb394_8 ns394 0 ni8 0 -5.66981737855
Gb395_8 ns395 0 ni8 0 1.70052379695
Gb396_8 ns396 0 ni8 0 1.58977849418
Gb397_8 ns397 0 ni8 0 1.86936465941
Gb398_8 ns398 0 ni8 0 0.918326016818
Gb399_8 ns399 0 ni8 0 1.86091951073
Gb400_8 ns400 0 ni8 0 -0.0696438180465
Gb401_8 ns401 0 ni8 0 1.7715070455
Gb402_8 ns402 0 ni8 0 0.919848034492
Gb403_8 ns403 0 ni8 0 -0.760413119527
Gb404_8 ns404 0 ni8 0 -1.73462525062
Gb405_8 ns405 0 ni8 0 1.66554798658
Gb406_8 ns406 0 ni8 0 -0.962084218547
Gb407_8 ns407 0 ni8 0 0.881978685923
Gb408_8 ns408 0 ni8 0 1.60046667014
Gb409_8 ns409 0 ni8 0 -1.55772849734
Gb410_8 ns410 0 ni8 0 0.747487499417
Gb411_8 ns411 0 ni8 0 -1.15723265214
Gb412_8 ns412 0 ni8 0 -1.4722884914
Gb413_8 ns413 0 ni8 0 -1.43065334637
Gb414_8 ns414 0 ni8 0 0.877735034392
Gb415_8 ns415 0 ni8 0 -0.0366302966022
Gb416_8 ns416 0 ni8 0 -1.3954618059
Gb417_8 ns417 0 ni8 0 1.30856229812
Gb418_8 ns418 0 ni8 0 0.486068116494
Gb419_8 ns419 0 ni8 0 -1.08772879245
Gb420_8 ns420 0 ni8 0 1.2550657279
Gb421_8 ns421 0 ni8 0 0.406136520382
Gb422_8 ns422 0 ni8 0 1.19813246552
Gb423_8 ns423 0 ni8 0 1.09813888731
Gb424_8 ns424 0 ni8 0 -0.927025586813
Gb425_8 ns425 0 ni8 0 -0.772633145912
Gb426_8 ns426 0 ni8 0 0.961527123453
Gb427_8 ns427 0 ni8 0 -0.623541296567
Gb428_8 ns428 0 ni8 0 0.920112973699
Gb429_8 ns429 0 ni8 0 -0.197470289704
Gb430_8 ns430 0 ni8 0 0.819693134289
Gb431_8 ns431 0 ni8 0 -0.752268145323
Gb432_8 ns432 0 ni8 0 -0.0518715051145
Gb433_8 ns433 0 ni8 0 -0.181587927011
Gb434_8 ns434 0 ni8 0 0.694608973231
Gb435_8 ns435 0 ni8 0 0.169134997258
Gb436_8 ns436 0 ni8 0 -0.574504157078
Gb437_8 ns437 0 ni8 0 -0.423994579197
Gb438_8 ns438 0 ni8 0 -0.24090789391
Gb439_8 ns439 0 ni8 0 0.374937946713
Gb440_8 ns440 0 ni8 0 -0.168660279104
Gb441_8 ns441 0 ni8 0 -0.0301538467221
Gb442_8 ns442 0 ni8 0 0.219310234788
Gb443_8 ns443 0 ni8 0 -0.12047842402
Gb444_8 ns444 0 ni8 0 0.0870596730425
Gb445_8 ns445 0 ni8 0 -0.076966070616
Gb446_8 ns446 0 ni8 0 -0.0100700165577
Gb447_8 ns447 0 ni8 0 0.0781839687698
Gb448_8 ns448 0 ni8 0 -0.016866442929

Gc1_1 0 n2 ns1 0 0.00369806103109
Gc1_2 0 n2 ns2 0 0.0104527094516
Gc1_3 0 n2 ns3 0 -0.00224636466692
Gc1_4 0 n2 ns4 0 -0.00073109990534
Gc1_5 0 n2 ns5 0 3.2555052134e-05
Gc1_6 0 n2 ns6 0 -4.21042803167e-06
Gc1_7 0 n2 ns7 0 0.000115349239321
Gc1_8 0 n2 ns8 0 4.00353470897e-05
Gc1_9 0 n2 ns9 0 5.39357528842e-07
Gc1_10 0 n2 ns10 0 -1.66528609323e-06
Gc1_11 0 n2 ns11 0 -6.66681081322e-05
Gc1_12 0 n2 ns12 0 -4.99565455639e-05
Gc1_13 0 n2 ns13 0 0.000201016483729
Gc1_14 0 n2 ns14 0 5.97964589825e-06
Gc1_15 0 n2 ns15 0 1.93916964675e-06
Gc1_16 0 n2 ns16 0 -1.82275763039e-06
Gc1_17 0 n2 ns17 0 -7.78747926129e-06
Gc1_18 0 n2 ns18 0 6.57565708722e-05
Gc1_19 0 n2 ns19 0 8.06005504227e-06
Gc1_20 0 n2 ns20 0 -0.000163723517451
Gc1_21 0 n2 ns21 0 4.43459362241e-06
Gc1_22 0 n2 ns22 0 3.75298071107e-06
Gc1_23 0 n2 ns23 0 -0.000102902705706
Gc1_24 0 n2 ns24 0 -1.43442557266e-05
Gc1_25 0 n2 ns25 0 9.97098426337e-05
Gc1_26 0 n2 ns26 0 8.17033536817e-05
Gc1_27 0 n2 ns27 0 2.44167536854e-05
Gc1_28 0 n2 ns28 0 -3.8636148896e-06
Gc1_29 0 n2 ns29 0 3.16603098128e-05
Gc1_30 0 n2 ns30 0 -0.000157490105753
Gc1_31 0 n2 ns31 0 0.000169694578529
Gc1_32 0 n2 ns32 0 1.68744093519e-05
Gc1_33 0 n2 ns33 0 0.000208437626597
Gc1_34 0 n2 ns34 0 -5.82012154143e-05
Gc1_35 0 n2 ns35 0 -0.000355941820447
Gc1_36 0 n2 ns36 0 4.51864098801e-05
Gc1_37 0 n2 ns37 0 0.000221133412274
Gc1_38 0 n2 ns38 0 3.15629145631e-05
Gc1_39 0 n2 ns39 0 -0.000104482818764
Gc1_40 0 n2 ns40 0 -0.000339092381773
Gc1_41 0 n2 ns41 0 -0.000618613746476
Gc1_42 0 n2 ns42 0 -0.000340882185462
Gc1_43 0 n2 ns43 0 0.000896137199457
Gc1_44 0 n2 ns44 0 -0.000934412959587
Gc1_45 0 n2 ns45 0 0.000400457168841
Gc1_46 0 n2 ns46 0 0.000529023457326
Gc1_47 0 n2 ns47 0 0.00316491057537
Gc1_48 0 n2 ns48 0 0.000394119210061
Gc1_49 0 n2 ns49 0 -0.00046723804503
Gc1_50 0 n2 ns50 0 0.00379838945451
Gc1_51 0 n2 ns51 0 -0.00103388252821
Gc1_52 0 n2 ns52 0 -0.00157045440381
Gc1_53 0 n2 ns53 0 -0.0108233436981
Gc1_54 0 n2 ns54 0 -0.000579659479837
Gc1_55 0 n2 ns55 0 7.60329198079e-05
Gc1_56 0 n2 ns56 0 0.000129045329924
Gc1_57 0 n2 ns57 0 -0.00150083293601
Gc1_58 0 n2 ns58 0 -0.000712029848715
Gc1_59 0 n2 ns59 0 0.000553180220668
Gc1_60 0 n2 ns60 0 0.000738508285766
Gc1_61 0 n2 ns61 0 2.35632607668e-05
Gc1_62 0 n2 ns62 0 6.87203464492e-06
Gc1_63 0 n2 ns63 0 0.00019581284379
Gc1_64 0 n2 ns64 0 3.37816861617e-05
Gc1_65 0 n2 ns65 0 -8.86295904924e-07
Gc1_66 0 n2 ns66 0 1.19188980953e-06
Gc1_67 0 n2 ns67 0 6.81293035502e-06
Gc1_68 0 n2 ns68 0 0.000152261307615
Gc1_69 0 n2 ns69 0 0.000257642898551
Gc1_70 0 n2 ns70 0 -0.000132633711811
Gc1_71 0 n2 ns71 0 -1.8802039681e-06
Gc1_72 0 n2 ns72 0 -1.45215167151e-07
Gc1_73 0 n2 ns73 0 0.000162567266235
Gc1_74 0 n2 ns74 0 -2.57926333884e-05
Gc1_75 0 n2 ns75 0 -0.000173264862543
Gc1_76 0 n2 ns76 0 -0.0002963067644
Gc1_77 0 n2 ns77 0 2.36021354259e-06
Gc1_78 0 n2 ns78 0 -6.59189384198e-06
Gc1_79 0 n2 ns79 0 -5.94273873232e-05
Gc1_80 0 n2 ns80 0 0.000192965638945
Gc1_81 0 n2 ns81 0 0.000387709353381
Gc1_82 0 n2 ns82 0 0.000206466517786
Gc1_83 0 n2 ns83 0 -1.41571240007e-05
Gc1_84 0 n2 ns84 0 -4.82287624379e-05
Gc1_85 0 n2 ns85 0 4.12078464791e-05
Gc1_86 0 n2 ns86 0 -0.0002663113761
Gc1_87 0 n2 ns87 0 0.000541635876238
Gc1_88 0 n2 ns88 0 -0.000132936869068
Gc1_89 0 n2 ns89 0 0.000736928770937
Gc1_90 0 n2 ns90 0 -5.5229880664e-05
Gc1_91 0 n2 ns91 0 -0.000608559461572
Gc1_92 0 n2 ns92 0 0.000179071000199
Gc1_93 0 n2 ns93 0 0.00059277561071
Gc1_94 0 n2 ns94 0 -0.000193668612987
Gc1_95 0 n2 ns95 0 -0.00021175019436
Gc1_96 0 n2 ns96 0 -0.000250126093253
Gc1_97 0 n2 ns97 0 -0.00114631455686
Gc1_98 0 n2 ns98 0 -0.00100554469944
Gc1_99 0 n2 ns99 0 0.000463723103531
Gc1_100 0 n2 ns100 0 -0.00112147381342
Gc1_101 0 n2 ns101 0 0.00102869127475
Gc1_102 0 n2 ns102 0 0.000652420370184
Gc1_103 0 n2 ns103 0 0.00272525155328
Gc1_104 0 n2 ns104 0 -2.99124238856e-05
Gc1_105 0 n2 ns105 0 0.000626733954415
Gc1_106 0 n2 ns106 0 0.00241184267418
Gc1_107 0 n2 ns107 0 -0.000145555388375
Gc1_108 0 n2 ns108 0 -0.00226600360126
Gc1_109 0 n2 ns109 0 -0.00679508193571
Gc1_110 0 n2 ns110 0 -0.000652169222486
Gc1_111 0 n2 ns111 0 4.34954243075e-05
Gc1_112 0 n2 ns112 0 0.000115091684013
Gc1_113 0 n2 ns113 0 0.0317479435274
Gc1_114 0 n2 ns114 0 -0.00566734254214
Gc1_115 0 n2 ns115 0 -0.000892773168243
Gc1_116 0 n2 ns116 0 0.00147228359469
Gc1_117 0 n2 ns117 0 -1.83923766583e-05
Gc1_118 0 n2 ns118 0 -3.0776397547e-05
Gc1_119 0 n2 ns119 0 -1.54176153257e-05
Gc1_120 0 n2 ns120 0 -2.64761912082e-05
Gc1_121 0 n2 ns121 0 2.43661152618e-07
Gc1_122 0 n2 ns122 0 2.18529764879e-07
Gc1_123 0 n2 ns123 0 -2.82773850367e-05
Gc1_124 0 n2 ns124 0 -0.000295720868768
Gc1_125 0 n2 ns125 0 -5.99674963906e-05
Gc1_126 0 n2 ns126 0 -0.000154048828015
Gc1_127 0 n2 ns127 0 -6.34615965248e-07
Gc1_128 0 n2 ns128 0 4.39843890546e-08
Gc1_129 0 n2 ns129 0 -0.000326051317418
Gc1_130 0 n2 ns130 0 4.2460248437e-05
Gc1_131 0 n2 ns131 0 -0.000115201033408
Gc1_132 0 n2 ns132 0 8.47285052203e-05
Gc1_133 0 n2 ns133 0 2.65225178495e-06
Gc1_134 0 n2 ns134 0 -2.39527547254e-06
Gc1_135 0 n2 ns135 0 0.000152180673408
Gc1_136 0 n2 ns136 0 -0.000387525668865
Gc1_137 0 n2 ns137 0 -4.07175490611e-05
Gc1_138 0 n2 ns138 0 -0.000212386475723
Gc1_139 0 n2 ns139 0 1.47516945652e-05
Gc1_140 0 n2 ns140 0 -4.45407115372e-05
Gc1_141 0 n2 ns141 0 -0.000314348399694
Gc1_142 0 n2 ns142 0 0.000686418383928
Gc1_143 0 n2 ns143 0 -0.000142379408116
Gc1_144 0 n2 ns144 0 -0.000164643022678
Gc1_145 0 n2 ns145 0 -0.00114106916308
Gc1_146 0 n2 ns146 0 7.48325912119e-06
Gc1_147 0 n2 ns147 0 0.000374364871754
Gc1_148 0 n2 ns148 0 0.000435372113456
Gc1_149 0 n2 ns149 0 -0.000741625635109
Gc1_150 0 n2 ns150 0 -1.61975552166e-05
Gc1_151 0 n2 ns151 0 -0.000249572115371
Gc1_152 0 n2 ns152 0 5.30643776428e-05
Gc1_153 0 n2 ns153 0 -4.56604314088e-06
Gc1_154 0 n2 ns154 0 0.0026486438625
Gc1_155 0 n2 ns155 0 -0.00104078663186
Gc1_156 0 n2 ns156 0 -0.000249590357153
Gc1_157 0 n2 ns157 0 0.00016964518514
Gc1_158 0 n2 ns158 0 -0.000973675667029
Gc1_159 0 n2 ns159 0 -1.17549588131e-05
Gc1_160 0 n2 ns160 0 -0.00206171170184
Gc1_161 0 n2 ns161 0 0.00104342764699
Gc1_162 0 n2 ns162 0 0.000181607898849
Gc1_163 0 n2 ns163 0 -0.000305659495005
Gc1_164 0 n2 ns164 0 -4.87943377142e-05
Gc1_165 0 n2 ns165 0 -0.000936710201036
Gc1_166 0 n2 ns166 0 -0.00016535698565
Gc1_167 0 n2 ns167 0 5.10584037183e-05
Gc1_168 0 n2 ns168 0 2.61906779243e-05
Gc1_169 0 n2 ns169 0 0.0227101861485
Gc1_170 0 n2 ns170 0 0.000252996112811
Gc1_171 0 n2 ns171 0 0.000313553864158
Gc1_172 0 n2 ns172 0 0.000213661539433
Gc1_173 0 n2 ns173 0 -1.14417890485e-05
Gc1_174 0 n2 ns174 0 -1.45605182577e-05
Gc1_175 0 n2 ns175 0 0.000115321621895
Gc1_176 0 n2 ns176 0 -8.80107309161e-05
Gc1_177 0 n2 ns177 0 -4.30874990824e-07
Gc1_178 0 n2 ns178 0 1.16519609065e-08
Gc1_179 0 n2 ns179 0 4.19954881774e-05
Gc1_180 0 n2 ns180 0 8.18938145387e-05
Gc1_181 0 n2 ns181 0 2.2895312422e-06
Gc1_182 0 n2 ns182 0 -0.000149815986488
Gc1_183 0 n2 ns183 0 -2.64519115581e-07
Gc1_184 0 n2 ns184 0 5.06272825587e-07
Gc1_185 0 n2 ns185 0 9.71814537257e-05
Gc1_186 0 n2 ns186 0 -6.63304566258e-05
Gc1_187 0 n2 ns187 0 -0.000161370523731
Gc1_188 0 n2 ns188 0 3.56457738963e-06
Gc1_189 0 n2 ns189 0 -4.59885355616e-06
Gc1_190 0 n2 ns190 0 1.73183418398e-06
Gc1_191 0 n2 ns191 0 1.8582819906e-05
Gc1_192 0 n2 ns192 0 0.00017731539299
Gc1_193 0 n2 ns193 0 0.000122947851871
Gc1_194 0 n2 ns194 0 -0.000129442173987
Gc1_195 0 n2 ns195 0 -3.02355471798e-05
Gc1_196 0 n2 ns196 0 2.20079820178e-05
Gc1_197 0 n2 ns197 0 -0.000202226236905
Gc1_198 0 n2 ns198 0 -0.000199884995074
Gc1_199 0 n2 ns199 0 2.45909901249e-05
Gc1_200 0 n2 ns200 0 -0.000297659277266
Gc1_201 0 n2 ns201 0 -1.90554246537e-06
Gc1_202 0 n2 ns202 0 -0.000474808312243
Gc1_203 0 n2 ns203 0 -4.05709750416e-05
Gc1_204 0 n2 ns204 0 0.000425672874659
Gc1_205 0 n2 ns205 0 1.22322159137e-05
Gc1_206 0 n2 ns206 0 -0.000323476063872
Gc1_207 0 n2 ns207 0 -0.000233078367438
Gc1_208 0 n2 ns208 0 9.21151525724e-05
Gc1_209 0 n2 ns209 0 -0.000926543194293
Gc1_210 0 n2 ns210 0 0.000295381099375
Gc1_211 0 n2 ns211 0 -0.000507832454206
Gc1_212 0 n2 ns212 0 -0.000609503115568
Gc1_213 0 n2 ns213 0 0.00105144795345
Gc1_214 0 n2 ns214 0 -0.000407394487931
Gc1_215 0 n2 ns215 0 0.00108990280673
Gc1_216 0 n2 ns216 0 -0.00151594745577
Gc1_217 0 n2 ns217 0 0.0012315442259
Gc1_218 0 n2 ns218 0 0.000287143388338
Gc1_219 0 n2 ns219 0 -0.000146926211585
Gc1_220 0 n2 ns220 0 -0.000658281939951
Gc1_221 0 n2 ns221 0 -0.000754490766589
Gc1_222 0 n2 ns222 0 -0.000455181494338
Gc1_223 0 n2 ns223 0 1.89353179857e-05
Gc1_224 0 n2 ns224 0 5.15144839499e-05
Gc1_225 0 n2 ns225 0 -0.00966172151068
Gc1_226 0 n2 ns226 0 0.000617715295529
Gc1_227 0 n2 ns227 0 -0.000189719106142
Gc1_228 0 n2 ns228 0 -0.000279520994481
Gc1_229 0 n2 ns229 0 -2.28942177952e-05
Gc1_230 0 n2 ns230 0 -1.39529156186e-05
Gc1_231 0 n2 ns231 0 -0.000259321414656
Gc1_232 0 n2 ns232 0 -5.45994262233e-05
Gc1_233 0 n2 ns233 0 8.68904101655e-07
Gc1_234 0 n2 ns234 0 -5.04552926884e-07
Gc1_235 0 n2 ns235 0 -8.57746956088e-05
Gc1_236 0 n2 ns236 0 -0.000164894642949
Gc1_237 0 n2 ns237 0 0.000310311932316
Gc1_238 0 n2 ns238 0 -0.00010835421427
Gc1_239 0 n2 ns239 0 -2.02825546609e-06
Gc1_240 0 n2 ns240 0 -2.88035490802e-07
Gc1_241 0 n2 ns241 0 0.000157510864562
Gc1_242 0 n2 ns242 0 -0.000124317490443
Gc1_243 0 n2 ns243 0 0.000114590777935
Gc1_244 0 n2 ns244 0 0.000341523587852
Gc1_245 0 n2 ns245 0 -4.11029486219e-07
Gc1_246 0 n2 ns246 0 5.58709465247e-06
Gc1_247 0 n2 ns247 0 -8.59898677202e-05
Gc1_248 0 n2 ns248 0 -0.000284721300619
Gc1_249 0 n2 ns249 0 0.000325490969875
Gc1_250 0 n2 ns250 0 0.000267354688955
Gc1_251 0 n2 ns251 0 -1.59236413009e-05
Gc1_252 0 n2 ns252 0 -3.93975738668e-05
Gc1_253 0 n2 ns253 0 -0.000305126383778
Gc1_254 0 n2 ns254 0 -0.000371657087839
Gc1_255 0 n2 ns255 0 -0.000524819480409
Gc1_256 0 n2 ns256 0 1.98940482599e-05
Gc1_257 0 n2 ns257 0 -0.00077621166762
Gc1_258 0 n2 ns258 0 0.000590387776211
Gc1_259 0 n2 ns259 0 -0.000659473976885
Gc1_260 0 n2 ns260 0 0.000178371652106
Gc1_261 0 n2 ns261 0 0.000112936792538
Gc1_262 0 n2 ns262 0 -0.000386725767731
Gc1_263 0 n2 ns263 0 1.95854659968e-05
Gc1_264 0 n2 ns264 0 0.000574141097606
Gc1_265 0 n2 ns265 0 0.00335828708546
Gc1_266 0 n2 ns266 0 0.00124133495034
Gc1_267 0 n2 ns267 0 0.00138851272202
Gc1_268 0 n2 ns268 0 -0.000920572207948
Gc1_269 0 n2 ns269 0 0.00132369687584
Gc1_270 0 n2 ns270 0 0.00258130321443
Gc1_271 0 n2 ns271 0 -0.00615030033648
Gc1_272 0 n2 ns272 0 0.000910758076294
Gc1_273 0 n2 ns273 0 -0.0018580073608
Gc1_274 0 n2 ns274 0 0.00569935780143
Gc1_275 0 n2 ns275 0 -0.00438175636761
Gc1_276 0 n2 ns276 0 -0.00320746930265
Gc1_277 0 n2 ns277 0 0.0207123632397
Gc1_278 0 n2 ns278 0 -0.000329574644999
Gc1_279 0 n2 ns279 0 8.31133489701e-05
Gc1_280 0 n2 ns280 0 -3.26485408274e-05
Gc1_281 0 n2 ns281 0 -0.0126484597542
Gc1_282 0 n2 ns282 0 0.000585895236543
Gc1_283 0 n2 ns283 0 0.000327963028486
Gc1_284 0 n2 ns284 0 0.00024080086643
Gc1_285 0 n2 ns285 0 -2.12048966015e-05
Gc1_286 0 n2 ns286 0 -9.93004443589e-06
Gc1_287 0 n2 ns287 0 -0.00027357223597
Gc1_288 0 n2 ns288 0 3.13901081183e-06
Gc1_289 0 n2 ns289 0 -1.42175584013e-06
Gc1_290 0 n2 ns290 0 5.23017769363e-07
Gc1_291 0 n2 ns291 0 9.5274004951e-06
Gc1_292 0 n2 ns292 0 0.000207241298844
Gc1_293 0 n2 ns293 0 0.000237000140479
Gc1_294 0 n2 ns294 0 -9.88605076424e-05
Gc1_295 0 n2 ns295 0 3.12550833378e-06
Gc1_296 0 n2 ns296 0 1.73444028972e-06
Gc1_297 0 n2 ns297 0 -0.000192407137966
Gc1_298 0 n2 ns298 0 5.47395411463e-05
Gc1_299 0 n2 ns299 0 0.000120413678937
Gc1_300 0 n2 ns300 0 0.0002898350722
Gc1_301 0 n2 ns301 0 6.12392087772e-06
Gc1_302 0 n2 ns302 0 -5.30009815907e-06
Gc1_303 0 n2 ns303 0 -0.000171649890657
Gc1_304 0 n2 ns304 0 0.000289998646279
Gc1_305 0 n2 ns305 0 0.00032816521901
Gc1_306 0 n2 ns306 0 0.000102839135754
Gc1_307 0 n2 ns307 0 -2.09264100463e-05
Gc1_308 0 n2 ns308 0 4.4571816624e-05
Gc1_309 0 n2 ns309 0 -4.44075372091e-05
Gc1_310 0 n2 ns310 0 0.000649982552169
Gc1_311 0 n2 ns311 0 -0.000317639088581
Gc1_312 0 n2 ns312 0 0.000208207991826
Gc1_313 0 n2 ns313 0 0.00172281003269
Gc1_314 0 n2 ns314 0 0.000679346469732
Gc1_315 0 n2 ns315 0 -0.000142080687521
Gc1_316 0 n2 ns316 0 0.000364004965674
Gc1_317 0 n2 ns317 0 -0.000712564159947
Gc1_318 0 n2 ns318 0 -4.17447664382e-05
Gc1_319 0 n2 ns319 0 0.000336362298967
Gc1_320 0 n2 ns320 0 0.000236315056839
Gc1_321 0 n2 ns321 0 0.00121220443255
Gc1_322 0 n2 ns322 0 -0.00411692024667
Gc1_323 0 n2 ns323 0 -0.000132273682201
Gc1_324 0 n2 ns324 0 -0.00114382229382
Gc1_325 0 n2 ns325 0 0.000860023698305
Gc1_326 0 n2 ns326 0 -0.00245877524473
Gc1_327 0 n2 ns327 0 -5.32256664087e-05
Gc1_328 0 n2 ns328 0 0.0012648311598
Gc1_329 0 n2 ns329 0 0.0023214853408
Gc1_330 0 n2 ns330 0 0.00205859599595
Gc1_331 0 n2 ns331 0 0.00321799582808
Gc1_332 0 n2 ns332 0 0.00155576731052
Gc1_333 0 n2 ns333 0 0.00445567155029
Gc1_334 0 n2 ns334 0 0.000608808856709
Gc1_335 0 n2 ns335 0 -9.1384099696e-05
Gc1_336 0 n2 ns336 0 -0.000102851709794
Gc1_337 0 n2 ns337 0 0.00409734366931
Gc1_338 0 n2 ns338 0 7.53274624201e-05
Gc1_339 0 n2 ns339 0 -0.0001925276575
Gc1_340 0 n2 ns340 0 -0.000281888294167
Gc1_341 0 n2 ns341 0 1.15191095232e-05
Gc1_342 0 n2 ns342 0 2.80361658913e-05
Gc1_343 0 n2 ns343 0 4.65418804038e-05
Gc1_344 0 n2 ns344 0 3.30192256893e-05
Gc1_345 0 n2 ns345 0 -1.40483504293e-07
Gc1_346 0 n2 ns346 0 -2.33157347819e-07
Gc1_347 0 n2 ns347 0 8.3660109655e-06
Gc1_348 0 n2 ns348 0 -0.000267058507058
Gc1_349 0 n2 ns349 0 -9.07101515215e-05
Gc1_350 0 n2 ns350 0 -0.000114723127044
Gc1_351 0 n2 ns351 0 9.53180468036e-07
Gc1_352 0 n2 ns352 0 1.66924929894e-07
Gc1_353 0 n2 ns353 0 0.000297065079272
Gc1_354 0 n2 ns354 0 -3.37958887128e-05
Gc1_355 0 n2 ns355 0 0.000128456600626
Gc1_356 0 n2 ns356 0 -0.000124799703635
Gc1_357 0 n2 ns357 0 1.80547421221e-07
Gc1_358 0 n2 ns358 0 -3.69319149617e-06
Gc1_359 0 n2 ns359 0 0.000179774225755
Gc1_360 0 n2 ns360 0 -0.000432063701159
Gc1_361 0 n2 ns361 0 2.59763628944e-05
Gc1_362 0 n2 ns362 0 -0.000219573337906
Gc1_363 0 n2 ns363 0 -1.92926076886e-06
Gc1_364 0 n2 ns364 0 1.02210467797e-05
Gc1_365 0 n2 ns365 0 -1.04569665499e-06
Gc1_366 0 n2 ns366 0 -0.00083492949017
Gc1_367 0 n2 ns367 0 0.000157715751775
Gc1_368 0 n2 ns368 0 0.000414545927534
Gc1_369 0 n2 ns369 0 -0.00160918062618
Gc1_370 0 n2 ns370 0 -0.000276104394061
Gc1_371 0 n2 ns371 0 0.000142011580891
Gc1_372 0 n2 ns372 0 0.000546320755486
Gc1_373 0 n2 ns373 0 0.000525648113556
Gc1_374 0 n2 ns374 0 0.000188863922737
Gc1_375 0 n2 ns375 0 0.000372140555034
Gc1_376 0 n2 ns376 0 -0.000194985837207
Gc1_377 0 n2 ns377 0 -0.000740162367362
Gc1_378 0 n2 ns378 0 0.0022425316445
Gc1_379 0 n2 ns379 0 -0.000798006865506
Gc1_380 0 n2 ns380 0 -0.000246905585307
Gc1_381 0 n2 ns381 0 -0.00181660719123
Gc1_382 0 n2 ns382 0 0.00180810924652
Gc1_383 0 n2 ns383 0 -0.0012087729968
Gc1_384 0 n2 ns384 0 0.00117321064183
Gc1_385 0 n2 ns385 0 0.00145331325472
Gc1_386 0 n2 ns386 0 -0.000441792489436
Gc1_387 0 n2 ns387 0 0.00152084955402
Gc1_388 0 n2 ns388 0 -0.000928296053423
Gc1_389 0 n2 ns389 0 0.00176741033471
Gc1_390 0 n2 ns390 0 0.000105947790536
Gc1_391 0 n2 ns391 0 -4.3779143787e-05
Gc1_392 0 n2 ns392 0 2.9404718998e-05
Gc1_393 0 n2 ns393 0 -0.000712891644551
Gc1_394 0 n2 ns394 0 -0.000223360699531
Gc1_395 0 n2 ns395 0 0.000253241783296
Gc1_396 0 n2 ns396 0 0.000131396910427
Gc1_397 0 n2 ns397 0 -2.17024156986e-07
Gc1_398 0 n2 ns398 0 1.61885920977e-05
Gc1_399 0 n2 ns399 0 -3.36215959114e-05
Gc1_400 0 n2 ns400 0 7.31846856361e-05
Gc1_401 0 n2 ns401 0 5.29574467417e-08
Gc1_402 0 n2 ns402 0 1.50539720742e-07
Gc1_403 0 n2 ns403 0 6.45795686073e-05
Gc1_404 0 n2 ns404 0 0.000124457188913
Gc1_405 0 n2 ns405 0 -5.2077960216e-05
Gc1_406 0 n2 ns406 0 -9.00033810885e-05
Gc1_407 0 n2 ns407 0 1.98103925914e-08
Gc1_408 0 n2 ns408 0 -1.33386402439e-06
Gc1_409 0 n2 ns409 0 -9.1532224808e-05
Gc1_410 0 n2 ns410 0 9.72016315306e-05
Gc1_411 0 n2 ns411 0 0.000122148250941
Gc1_412 0 n2 ns412 0 -4.01991776859e-05
Gc1_413 0 n2 ns413 0 -6.61082151308e-06
Gc1_414 0 n2 ns414 0 3.30653471385e-06
Gc1_415 0 n2 ns415 0 1.33371448039e-05
Gc1_416 0 n2 ns416 0 0.00019413014861
Gc1_417 0 n2 ns417 0 9.61870045224e-05
Gc1_418 0 n2 ns418 0 -0.000208595143738
Gc1_419 0 n2 ns419 0 2.7401307316e-05
Gc1_420 0 n2 ns420 0 -3.77953777512e-05
Gc1_421 0 n2 ns421 0 0.000241617432218
Gc1_422 0 n2 ns422 0 0.000157219759174
Gc1_423 0 n2 ns423 0 2.80094502816e-05
Gc1_424 0 n2 ns424 0 0.000131200188841
Gc1_425 0 n2 ns425 0 0.000111522044076
Gc1_426 0 n2 ns426 0 -0.000695226331731
Gc1_427 0 n2 ns427 0 0.000119320283825
Gc1_428 0 n2 ns428 0 0.000189587806302
Gc1_429 0 n2 ns429 0 1.96324455686e-05
Gc1_430 0 n2 ns430 0 0.000366493539643
Gc1_431 0 n2 ns431 0 0.000188975086354
Gc1_432 0 n2 ns432 0 -0.000143575537976
Gc1_433 0 n2 ns433 0 -0.00110363520368
Gc1_434 0 n2 ns434 0 2.04437484336e-05
Gc1_435 0 n2 ns435 0 -0.00064668442435
Gc1_436 0 n2 ns436 0 -0.000330883108359
Gc1_437 0 n2 ns437 0 -0.00128365506501
Gc1_438 0 n2 ns438 0 0.000172293676888
Gc1_439 0 n2 ns439 0 -0.000536367293194
Gc1_440 0 n2 ns440 0 0.000866856088156
Gc1_441 0 n2 ns441 0 0.00142601029278
Gc1_442 0 n2 ns442 0 5.91964808875e-06
Gc1_443 0 n2 ns443 0 0.0011063320393
Gc1_444 0 n2 ns444 0 -0.00024784266722
Gc1_445 0 n2 ns445 0 0.00104576635329
Gc1_446 0 n2 ns446 0 0.00037466222517
Gc1_447 0 n2 ns447 0 -3.4030159137e-05
Gc1_448 0 n2 ns448 0 -1.74255837276e-05
Gd1_1 0 n2 ni1 0 -0.00411277433817
Gd1_2 0 n2 ni2 0 0.00504122796507
Gd1_3 0 n2 ni3 0 0.00314464607336
Gd1_4 0 n2 ni4 0 -0.000949927881092
Gd1_5 0 n2 ni5 0 -0.000469964997314
Gd1_6 0 n2 ni6 0 -0.000111447854493
Gd1_7 0 n2 ni7 0 -0.00018079886118
Gd1_8 0 n2 ni8 0 0.000202727455259
Gc2_1 0 n4 ns1 0 -0.00150083634578
Gc2_2 0 n4 ns2 0 -0.000712029687613
Gc2_3 0 n4 ns3 0 0.000553181219671
Gc2_4 0 n4 ns4 0 0.000738507811836
Gc2_5 0 n4 ns5 0 2.35632438805e-05
Gc2_6 0 n4 ns6 0 6.8720215469e-06
Gc2_7 0 n4 ns7 0 0.000195812866605
Gc2_8 0 n4 ns8 0 3.37818366334e-05
Gc2_9 0 n4 ns9 0 -8.86293633062e-07
Gc2_10 0 n4 ns10 0 1.19189605664e-06
Gc2_11 0 n4 ns11 0 6.81288021792e-06
Gc2_12 0 n4 ns12 0 0.000152261313912
Gc2_13 0 n4 ns13 0 0.000257642790124
Gc2_14 0 n4 ns14 0 -0.000132633772678
Gc2_15 0 n4 ns15 0 -1.8802072958e-06
Gc2_16 0 n4 ns16 0 -1.45221507166e-07
Gc2_17 0 n4 ns17 0 0.000162567373706
Gc2_18 0 n4 ns18 0 -2.57925740819e-05
Gc2_19 0 n4 ns19 0 -0.000173264680285
Gc2_20 0 n4 ns20 0 -0.000296306765568
Gc2_21 0 n4 ns21 0 2.3602090831e-06
Gc2_22 0 n4 ns22 0 -6.59188386061e-06
Gc2_23 0 n4 ns23 0 -5.942759225e-05
Gc2_24 0 n4 ns24 0 0.000192965871461
Gc2_25 0 n4 ns25 0 0.000387709516024
Gc2_26 0 n4 ns26 0 0.00020646650028
Gc2_27 0 n4 ns27 0 -1.41570320889e-05
Gc2_28 0 n4 ns28 0 -4.82288305765e-05
Gc2_29 0 n4 ns29 0 4.12076910095e-05
Gc2_30 0 n4 ns30 0 -0.000266311403732
Gc2_31 0 n4 ns31 0 0.000541635758719
Gc2_32 0 n4 ns32 0 -0.000132937037806
Gc2_33 0 n4 ns33 0 0.000736930143488
Gc2_34 0 n4 ns34 0 -5.52310126963e-05
Gc2_35 0 n4 ns35 0 -0.000608560433601
Gc2_36 0 n4 ns36 0 0.000179071085127
Gc2_37 0 n4 ns37 0 0.000592775850633
Gc2_38 0 n4 ns38 0 -0.000193669148582
Gc2_39 0 n4 ns39 0 -0.000211749773666
Gc2_40 0 n4 ns40 0 -0.000250126031673
Gc2_41 0 n4 ns41 0 -0.00114631790657
Gc2_42 0 n4 ns42 0 -0.00100554679589
Gc2_43 0 n4 ns43 0 0.000463724356143
Gc2_44 0 n4 ns44 0 -0.00112147614591
Gc2_45 0 n4 ns45 0 0.00102869330785
Gc2_46 0 n4 ns46 0 0.00065242001734
Gc2_47 0 n4 ns47 0 0.00272525397585
Gc2_48 0 n4 ns48 0 -2.99137776077e-05
Gc2_49 0 n4 ns49 0 0.00062673288111
Gc2_50 0 n4 ns50 0 0.00241184488656
Gc2_51 0 n4 ns51 0 -0.000145558305707
Gc2_52 0 n4 ns52 0 -0.00226600192637
Gc2_53 0 n4 ns53 0 -0.00679508499766
Gc2_54 0 n4 ns54 0 -0.000652170465316
Gc2_55 0 n4 ns55 0 4.34952899893e-05
Gc2_56 0 n4 ns56 0 0.000115091772052
Gc2_57 0 n4 ns57 0 0.0152228745686
Gc2_58 0 n4 ns58 0 0.0102379426874
Gc2_59 0 n4 ns59 0 -0.00245573485977
Gc2_60 0 n4 ns60 0 -0.000975381725303
Gc2_61 0 n4 ns61 0 2.23574114911e-05
Gc2_62 0 n4 ns62 0 -1.32731486962e-05
Gc2_63 0 n4 ns63 0 0.000179688408509
Gc2_64 0 n4 ns64 0 -9.55735165204e-06
Gc2_65 0 n4 ns65 0 3.77239204795e-06
Gc2_66 0 n4 ns66 0 1.37429729447e-06
Gc2_67 0 n4 ns67 0 -1.98621823563e-05
Gc2_68 0 n4 ns68 0 -4.97960601103e-05
Gc2_69 0 n4 ns69 0 0.000177298841876
Gc2_70 0 n4 ns70 0 -7.22002415793e-05
Gc2_71 0 n4 ns71 0 3.71857027148e-06
Gc2_72 0 n4 ns72 0 5.1036972257e-06
Gc2_73 0 n4 ns73 0 1.8978317079e-05
Gc2_74 0 n4 ns74 0 2.55522886304e-06
Gc2_75 0 n4 ns75 0 -6.82032346952e-05
Gc2_76 0 n4 ns76 0 -0.000113290134885
Gc2_77 0 n4 ns77 0 -1.29116316625e-05
Gc2_78 0 n4 ns78 0 1.0573404224e-05
Gc2_79 0 n4 ns79 0 -4.61204629269e-05
Gc2_80 0 n4 ns80 0 8.99487846215e-05
Gc2_81 0 n4 ns81 0 0.000111145833735
Gc2_82 0 n4 ns82 0 -6.23087457192e-05
Gc2_83 0 n4 ns83 0 -2.38204864401e-05
Gc2_84 0 n4 ns84 0 5.23756849373e-05
Gc2_85 0 n4 ns85 0 -0.000207753324369
Gc2_86 0 n4 ns86 0 -0.000316765615172
Gc2_87 0 n4 ns87 0 0.000100379864386
Gc2_88 0 n4 ns88 0 -0.00023206233766
Gc2_89 0 n4 ns89 0 5.69183779808e-06
Gc2_90 0 n4 ns90 0 -0.000575463759111
Gc2_91 0 n4 ns91 0 -0.000285587853092
Gc2_92 0 n4 ns92 0 0.000395601522847
Gc2_93 0 n4 ns93 0 2.0500038695e-05
Gc2_94 0 n4 ns94 0 -0.000222861126573
Gc2_95 0 n4 ns95 0 -0.000237840980644
Gc2_96 0 n4 ns96 0 -0.000203090285678
Gc2_97 0 n4 ns97 0 -0.00109165696763
Gc2_98 0 n4 ns98 0 0.000256326481441
Gc2_99 0 n4 ns99 0 0.000343286522172
Gc2_100 0 n4 ns100 0 -0.0009873858949
Gc2_101 0 n4 ns101 0 0.000842369281475
Gc2_102 0 n4 ns102 0 -1.14012938472e-05
Gc2_103 0 n4 ns103 0 0.00305298159007
Gc2_104 0 n4 ns104 0 -0.000484653588901
Gc2_105 0 n4 ns105 0 -0.000125605325026
Gc2_106 0 n4 ns106 0 0.00327022176338
Gc2_107 0 n4 ns107 0 -0.0013460689684
Gc2_108 0 n4 ns108 0 -0.00157035366545
Gc2_109 0 n4 ns109 0 -0.0100639547745
Gc2_110 0 n4 ns110 0 -0.000505576694458
Gc2_111 0 n4 ns111 0 6.28444570784e-05
Gc2_112 0 n4 ns112 0 6.68976461175e-05
Gc2_113 0 n4 ns113 0 0.0226511895128
Gc2_114 0 n4 ns114 0 0.000257076300197
Gc2_115 0 n4 ns115 0 0.00031375956115
Gc2_116 0 n4 ns116 0 0.000212387976176
Gc2_117 0 n4 ns117 0 -1.13828452161e-05
Gc2_118 0 n4 ns118 0 -1.45291708328e-05
Gc2_119 0 n4 ns119 0 0.00011528832745
Gc2_120 0 n4 ns120 0 -8.7910169235e-05
Gc2_121 0 n4 ns121 0 -4.24100366093e-07
Gc2_122 0 n4 ns122 0 2.57508089928e-08
Gc2_123 0 n4 ns123 0 4.22397829851e-05
Gc2_124 0 n4 ns124 0 8.22028649821e-05
Gc2_125 0 n4 ns125 0 2.54737830022e-06
Gc2_126 0 n4 ns126 0 -0.000149723812957
Gc2_127 0 n4 ns127 0 -2.63855328509e-07
Gc2_128 0 n4 ns128 0 5.30907931508e-07
Gc2_129 0 n4 ns129 0 9.74670925133e-05
Gc2_130 0 n4 ns130 0 -6.65740747955e-05
Gc2_131 0 n4 ns131 0 -0.000161382096396
Gc2_132 0 n4 ns132 0 3.30372977483e-06
Gc2_133 0 n4 ns133 0 -4.64523966318e-06
Gc2_134 0 n4 ns134 0 1.74800076898e-06
Gc2_135 0 n4 ns135 0 1.86769183004e-05
Gc2_136 0 n4 ns136 0 0.000177719125174
Gc2_137 0 n4 ns137 0 0.000123322552595
Gc2_138 0 n4 ns138 0 -0.000129264040101
Gc2_139 0 n4 ns139 0 -3.02655229688e-05
Gc2_140 0 n4 ns140 0 2.21821969651e-05
Gc2_141 0 n4 ns141 0 -0.000202368413196
Gc2_142 0 n4 ns142 0 -0.000200897389948
Gc2_143 0 n4 ns143 0 2.48147240686e-05
Gc2_144 0 n4 ns144 0 -0.000297788998967
Gc2_145 0 n4 ns145 0 -6.12304519604e-07
Gc2_146 0 n4 ns146 0 -0.000476087598351
Gc2_147 0 n4 ns147 0 -4.14267901017e-05
Gc2_148 0 n4 ns148 0 0.000425640911354
Gc2_149 0 n4 ns149 0 1.27394568078e-05
Gc2_150 0 n4 ns150 0 -0.000324163805592
Gc2_151 0 n4 ns151 0 -0.000232879794245
Gc2_152 0 n4 ns152 0 9.17384309721e-05
Gc2_153 0 n4 ns153 0 -0.000928693527406
Gc2_154 0 n4 ns154 0 0.000293814805434
Gc2_155 0 n4 ns155 0 -0.000506825242905
Gc2_156 0 n4 ns156 0 -0.000610192239648
Gc2_157 0 n4 ns157 0 0.00105222691792
Gc2_158 0 n4 ns158 0 -0.000406719574695
Gc2_159 0 n4 ns159 0 0.00109166610467
Gc2_160 0 n4 ns160 0 -0.0015148619021
Gc2_161 0 n4 ns161 0 0.00122937677166
Gc2_162 0 n4 ns162 0 0.000287536097154
Gc2_163 0 n4 ns163 0 -0.000149039665828
Gc2_164 0 n4 ns164 0 -0.000657366860858
Gc2_165 0 n4 ns165 0 -0.000757121036351
Gc2_166 0 n4 ns166 0 -0.000454976566239
Gc2_167 0 n4 ns167 0 1.89400563911e-05
Gc2_168 0 n4 ns168 0 5.1429927783e-05
Gc2_169 0 n4 ns169 0 0.0162265823181
Gc2_170 0 n4 ns170 0 -0.00290424643424
Gc2_171 0 n4 ns171 0 -0.000318656498967
Gc2_172 0 n4 ns172 0 0.00100347470728
Gc2_173 0 n4 ns173 0 2.91346667942e-08
Gc2_174 0 n4 ns174 0 -9.72618579984e-06
Gc2_175 0 n4 ns175 0 0.000115167260522
Gc2_176 0 n4 ns176 0 -9.78262182226e-06
Gc2_177 0 n4 ns177 0 -3.20049608245e-06
Gc2_178 0 n4 ns178 0 -2.35905308085e-06
Gc2_179 0 n4 ns179 0 -1.37137701917e-05
Gc2_180 0 n4 ns180 0 -0.000156417117927
Gc2_181 0 n4 ns181 0 8.22814075283e-05
Gc2_182 0 n4 ns182 0 -0.000161815580161
Gc2_183 0 n4 ns183 0 -2.51949112957e-06
Gc2_184 0 n4 ns184 0 -7.05993602523e-06
Gc2_185 0 n4 ns185 0 -0.000163901664466
Gc2_186 0 n4 ns186 0 1.919694761e-05
Gc2_187 0 n4 ns187 0 -0.000152775082257
Gc2_188 0 n4 ns188 0 -8.09313958229e-05
Gc2_189 0 n4 ns189 0 2.0184418756e-05
Gc2_190 0 n4 ns190 0 -9.65584278696e-06
Gc2_191 0 n4 ns191 0 8.76457344215e-05
Gc2_192 0 n4 ns192 0 -0.00019236810901
Gc2_193 0 n4 ns193 0 0.000159939824992
Gc2_194 0 n4 ns194 0 -1.66144004242e-05
Gc2_195 0 n4 ns195 0 4.3053223985e-05
Gc2_196 0 n4 ns196 0 -0.000102198170849
Gc2_197 0 n4 ns197 0 -0.000148628124684
Gc2_198 0 n4 ns198 0 0.000448250796228
Gc2_199 0 n4 ns199 0 0.000158098066742
Gc2_200 0 n4 ns200 0 -9.86568912802e-05
Gc2_201 0 n4 ns201 0 -0.000318073602041
Gc2_202 0 n4 ns202 0 0.000123268445041
Gc2_203 0 n4 ns203 0 -1.38524481664e-05
Gc2_204 0 n4 ns204 0 0.000313168543153
Gc2_205 0 n4 ns205 0 -6.37500985904e-05
Gc2_206 0 n4 ns206 0 -9.04978328799e-05
Gc2_207 0 n4 ns207 0 -0.000303355110595
Gc2_208 0 n4 ns208 0 -3.02031837208e-05
Gc2_209 0 n4 ns209 0 -0.000486259384807
Gc2_210 0 n4 ns210 0 0.000714371485811
Gc2_211 0 n4 ns211 0 -0.00043999261856
Gc2_212 0 n4 ns212 0 -0.000774921954807
Gc2_213 0 n4 ns213 0 0.000871592222131
Gc2_214 0 n4 ns214 0 -6.54507813513e-05
Gc2_215 0 n4 ns215 0 0.00150257473437
Gc2_216 0 n4 ns216 0 -0.00125654999482
Gc2_217 0 n4 ns217 0 0.00114353643125
Gc2_218 0 n4 ns218 0 0.00115298566484
Gc2_219 0 n4 ns219 0 -0.000214340277461
Gc2_220 0 n4 ns220 0 -0.00129388909763
Gc2_221 0 n4 ns221 0 -0.00352640070447
Gc2_222 0 n4 ns222 0 -0.000541183640441
Gc2_223 0 n4 ns223 0 4.33962937286e-05
Gc2_224 0 n4 ns224 0 7.30324693031e-05
Gc2_225 0 n4 ns225 0 -0.0126554205655
Gc2_226 0 n4 ns226 0 0.000588768052282
Gc2_227 0 n4 ns227 0 0.000327639723403
Gc2_228 0 n4 ns228 0 0.000240251125313
Gc2_229 0 n4 ns229 0 -2.11995694965e-05
Gc2_230 0 n4 ns230 0 -9.91490569251e-06
Gc2_231 0 n4 ns231 0 -0.000273638518861
Gc2_232 0 n4 ns232 0 2.9943678674e-06
Gc2_233 0 n4 ns233 0 -1.42597687832e-06
Gc2_234 0 n4 ns234 0 5.23320896656e-07
Gc2_235 0 n4 ns235 0 9.53029257685e-06
Gc2_236 0 n4 ns236 0 0.000207127822904
Gc2_237 0 n4 ns237 0 0.000237167848661
Gc2_238 0 n4 ns238 0 -9.88891036308e-05
Gc2_239 0 n4 ns239 0 3.12988331198e-06
Gc2_240 0 n4 ns240 0 1.73141820751e-06
Gc2_241 0 n4 ns241 0 -0.000192347724289
Gc2_242 0 n4 ns242 0 5.47382792491e-05
Gc2_243 0 n4 ns243 0 0.00012029289273
Gc2_244 0 n4 ns244 0 0.000290061063976
Gc2_245 0 n4 ns245 0 6.10825970771e-06
Gc2_246 0 n4 ns246 0 -5.30596222768e-06
Gc2_247 0 n4 ns247 0 -0.000171597747416
Gc2_248 0 n4 ns248 0 0.000289904230848
Gc2_249 0 n4 ns249 0 0.000328307629333
Gc2_250 0 n4 ns250 0 0.000102998441453
Gc2_251 0 n4 ns251 0 -2.08724904254e-05
Gc2_252 0 n4 ns252 0 4.45140807171e-05
Gc2_253 0 n4 ns253 0 -4.39907947317e-05
Gc2_254 0 n4 ns254 0 0.000649895657319
Gc2_255 0 n4 ns255 0 -0.000317779438102
Gc2_256 0 n4 ns256 0 0.000208029226967
Gc2_257 0 n4 ns257 0 0.00172349067931
Gc2_258 0 n4 ns258 0 0.000679334502299
Gc2_259 0 n4 ns259 0 -0.000142167447057
Gc2_260 0 n4 ns260 0 0.000363804655354
Gc2_261 0 n4 ns261 0 -0.000712277610681
Gc2_262 0 n4 ns262 0 -4.14707718258e-05
Gc2_263 0 n4 ns263 0 0.00033621347674
Gc2_264 0 n4 ns264 0 0.000236772661527
Gc2_265 0 n4 ns265 0 0.0012125835237
Gc2_266 0 n4 ns266 0 -0.00411906755247
Gc2_267 0 n4 ns267 0 -0.000132190869348
Gc2_268 0 n4 ns268 0 -0.00114373003795
Gc2_269 0 n4 ns269 0 0.000860686840001
Gc2_270 0 n4 ns270 0 -0.00245795106842
Gc2_271 0 n4 ns271 0 -5.326101649e-05
Gc2_272 0 n4 ns272 0 0.00126581764366
Gc2_273 0 n4 ns273 0 0.00232157258297
Gc2_274 0 n4 ns274 0 0.00205769741145
Gc2_275 0 n4 ns275 0 0.00321778026822
Gc2_276 0 n4 ns276 0 0.00155491908494
Gc2_277 0 n4 ns277 0 0.00445670443093
Gc2_278 0 n4 ns278 0 0.000608525177862
Gc2_279 0 n4 ns279 0 -9.1395666099e-05
Gc2_280 0 n4 ns280 0 -0.00010272195399
Gc2_281 0 n4 ns281 0 -0.00729026421527
Gc2_282 0 n4 ns282 0 -0.000258425324532
Gc2_283 0 n4 ns283 0 -0.000180797194688
Gc2_284 0 n4 ns284 0 -0.000113501968685
Gc2_285 0 n4 ns285 0 -1.74097609599e-05
Gc2_286 0 n4 ns286 0 -3.32163548727e-06
Gc2_287 0 n4 ns287 0 -0.000275694758993
Gc2_288 0 n4 ns288 0 -1.10137275123e-05
Gc2_289 0 n4 ns289 0 4.71336999647e-06
Gc2_290 0 n4 ns290 0 3.51765760354e-06
Gc2_291 0 n4 ns291 0 -2.53760375826e-05
Gc2_292 0 n4 ns292 0 -0.000137896245024
Gc2_293 0 n4 ns293 0 0.000270808123075
Gc2_294 0 n4 ns294 0 -0.00018468253216
Gc2_295 0 n4 ns295 0 -4.61977463294e-06
Gc2_296 0 n4 ns296 0 -1.12265516685e-05
Gc2_297 0 n4 ns297 0 0.00014982024781
Gc2_298 0 n4 ns298 0 -4.94715315477e-05
Gc2_299 0 n4 ns299 0 0.000211015439689
Gc2_300 0 n4 ns300 0 0.000289872121437
Gc2_301 0 n4 ns301 0 -2.73481805763e-05
Gc2_302 0 n4 ns302 0 1.53901462156e-05
Gc2_303 0 n4 ns303 0 -4.31805075642e-06
Gc2_304 0 n4 ns304 0 -0.000231976267844
Gc2_305 0 n4 ns305 0 0.000403837512631
Gc2_306 0 n4 ns306 0 0.000104618644261
Gc2_307 0 n4 ns307 0 5.25061131862e-05
Gc2_308 0 n4 ns308 0 -0.000121125800891
Gc2_309 0 n4 ns309 0 -5.35640081024e-05
Gc2_310 0 n4 ns310 0 -0.00045025015966
Gc2_311 0 n4 ns311 0 -0.00050207073712
Gc2_312 0 n4 ns312 0 8.26430658264e-05
Gc2_313 0 n4 ns313 0 -0.00138709120553
Gc2_314 0 n4 ns314 0 -0.00043626809257
Gc2_315 0 n4 ns315 0 -0.000657882363948
Gc2_316 0 n4 ns316 0 0.000373090479051
Gc2_317 0 n4 ns317 0 0.000340042132891
Gc2_318 0 n4 ns318 0 -2.57289841911e-05
Gc2_319 0 n4 ns319 0 0.000195902211657
Gc2_320 0 n4 ns320 0 0.0003249386078
Gc2_321 0 n4 ns321 0 0.0022818967757
Gc2_322 0 n4 ns322 0 0.00341304829494
Gc2_323 0 n4 ns323 0 0.000637614461182
Gc2_324 0 n4 ns324 0 -0.000932062329737
Gc2_325 0 n4 ns325 0 -1.75250677345e-05
Gc2_326 0 n4 ns326 0 0.00474196042268
Gc2_327 0 n4 ns327 0 -0.00693096430312
Gc2_328 0 n4 ns328 0 0.0019585980884
Gc2_329 0 n4 ns329 0 -0.00179584722234
Gc2_330 0 n4 ns330 0 0.00441459175241
Gc2_331 0 n4 ns331 0 -0.0051271866824
Gc2_332 0 n4 ns332 0 -0.00466612352263
Gc2_333 0 n4 ns333 0 0.0197683260162
Gc2_334 0 n4 ns334 0 -0.000394760283214
Gc2_335 0 n4 ns335 0 9.46163595335e-05
Gc2_336 0 n4 ns336 0 7.09160241694e-05
Gc2_337 0 n4 ns337 0 -0.000733989784565
Gc2_338 0 n4 ns338 0 -0.000221638263253
Gc2_339 0 n4 ns339 0 0.000253494793638
Gc2_340 0 n4 ns340 0 0.000131180778036
Gc2_341 0 n4 ns341 0 -2.20810513126e-07
Gc2_342 0 n4 ns342 0 1.61374342596e-05
Gc2_343 0 n4 ns343 0 -3.38400967191e-05
Gc2_344 0 n4 ns344 0 7.30227327851e-05
Gc2_345 0 n4 ns345 0 5.17453604586e-08
Gc2_346 0 n4 ns346 0 1.5725020808e-07
Gc2_347 0 n4 ns347 0 6.46504156831e-05
Gc2_348 0 n4 ns348 0 0.000124841133167
Gc2_349 0 n4 ns349 0 -5.17911419128e-05
Gc2_350 0 n4 ns350 0 -8.98810829068e-05
Gc2_351 0 n4 ns351 0 2.52198682593e-08
Gc2_352 0 n4 ns352 0 -1.33789563188e-06
Gc2_353 0 n4 ns353 0 -9.18622697583e-05
Gc2_354 0 n4 ns354 0 9.73568241626e-05
Gc2_355 0 n4 ns355 0 0.000122058547061
Gc2_356 0 n4 ns356 0 -3.97701849494e-05
Gc2_357 0 n4 ns357 0 -6.60400032602e-06
Gc2_358 0 n4 ns358 0 3.30414590975e-06
Gc2_359 0 n4 ns359 0 1.31289713151e-05
Gc2_360 0 n4 ns360 0 0.000194725151055
Gc2_361 0 n4 ns361 0 9.64034745865e-05
Gc2_362 0 n4 ns362 0 -0.000208345081493
Gc2_363 0 n4 ns363 0 2.73715105519e-05
Gc2_364 0 n4 ns364 0 -3.7729310028e-05
Gc2_365 0 n4 ns365 0 0.000241751944307
Gc2_366 0 n4 ns366 0 0.000157883810114
Gc2_367 0 n4 ns367 0 2.75567200961e-05
Gc2_368 0 n4 ns368 0 0.000130809894876
Gc2_369 0 n4 ns369 0 0.000114246166565
Gc2_370 0 n4 ns370 0 -0.000695420138377
Gc2_371 0 n4 ns371 0 0.00011901556436
Gc2_372 0 n4 ns372 0 0.000188874202395
Gc2_373 0 n4 ns373 0 1.90602597818e-05
Gc2_374 0 n4 ns374 0 0.000366364572317
Gc2_375 0 n4 ns375 0 0.000188703557749
Gc2_376 0 n4 ns376 0 -0.000143158646992
Gc2_377 0 n4 ns377 0 -0.00110329535532
Gc2_378 0 n4 ns378 0 1.65990624676e-05
Gc2_379 0 n4 ns379 0 -0.000646293001097
Gc2_380 0 n4 ns380 0 -0.000330619078001
Gc2_381 0 n4 ns381 0 -0.00128197768652
Gc2_382 0 n4 ns382 0 0.000170980663147
Gc2_383 0 n4 ns383 0 -0.000536350814461
Gc2_384 0 n4 ns384 0 0.000867322627112
Gc2_385 0 n4 ns385 0 0.00142266069139
Gc2_386 0 n4 ns386 0 4.43055725029e-06
Gc2_387 0 n4 ns387 0 0.00110385144611
Gc2_388 0 n4 ns388 0 -0.000245422824099
Gc2_389 0 n4 ns389 0 0.0010463496488
Gc2_390 0 n4 ns390 0 0.000374512103743
Gc2_391 0 n4 ns391 0 -3.41196668338e-05
Gc2_392 0 n4 ns392 0 -1.76165151439e-05
Gc2_393 0 n4 ns393 0 -0.00295378151157
Gc2_394 0 n4 ns394 0 0.000693701850963
Gc2_395 0 n4 ns395 0 -7.51054372629e-05
Gc2_396 0 n4 ns396 0 -0.000151998779279
Gc2_397 0 n4 ns397 0 -2.52960211893e-06
Gc2_398 0 n4 ns398 0 1.66989831648e-05
Gc2_399 0 n4 ns399 0 -0.000108906178228
Gc2_400 0 n4 ns400 0 3.40412708238e-05
Gc2_401 0 n4 ns401 0 -4.40632726761e-06
Gc2_402 0 n4 ns402 0 -4.11234678439e-06
Gc2_403 0 n4 ns403 0 2.00290931522e-06
Gc2_404 0 n4 ns404 0 -0.000182877566118
Gc2_405 0 n4 ns405 0 6.05376365416e-05
Gc2_406 0 n4 ns406 0 -0.000175912992237
Gc2_407 0 n4 ns407 0 4.34129687021e-06
Gc2_408 0 n4 ns408 0 1.08969947471e-05
Gc2_409 0 n4 ns409 0 0.000197481036365
Gc2_410 0 n4 ns410 0 -2.37865664095e-05
Gc2_411 0 n4 ns411 0 0.000192540820439
Gc2_412 0 n4 ns412 0 4.62276510281e-05
Gc2_413 0 n4 ns413 0 2.56829275836e-05
Gc2_414 0 n4 ns414 0 -1.39805354911e-05
Gc2_415 0 n4 ns415 0 8.30783661322e-05
Gc2_416 0 n4 ns416 0 -0.000305735376805
Gc2_417 0 n4 ns417 0 0.000218304986974
Gc2_418 0 n4 ns418 0 -0.00011148521247
Gc2_419 0 n4 ns419 0 -6.73764736944e-05
Gc2_420 0 n4 ns420 0 9.28990642603e-05
Gc2_421 0 n4 ns421 0 -0.000148415456944
Gc2_422 0 n4 ns422 0 -0.000412879474742
Gc2_423 0 n4 ns423 0 -2.44103079358e-05
Gc2_424 0 n4 ns424 0 0.000591866237994
Gc2_425 0 n4 ns425 0 -0.000450193257323
Gc2_426 0 n4 ns426 0 0.000604159508221
Gc2_427 0 n4 ns427 0 5.4562996005e-05
Gc2_428 0 n4 ns428 0 0.000795721117988
Gc2_429 0 n4 ns429 0 -4.94621470705e-05
Gc2_430 0 n4 ns430 0 4.71602626525e-05
Gc2_431 0 n4 ns431 0 0.00052735616285
Gc2_432 0 n4 ns432 0 -1.86246027367e-05
Gc2_433 0 n4 ns433 0 0.000719757198574
Gc2_434 0 n4 ns434 0 -0.000662006781434
Gc2_435 0 n4 ns435 0 -0.000710401382465
Gc2_436 0 n4 ns436 0 -0.000958716474241
Gc2_437 0 n4 ns437 0 -0.000589183765635
Gc2_438 0 n4 ns438 0 7.36992926372e-05
Gc2_439 0 n4 ns439 0 -0.000972452605325
Gc2_440 0 n4 ns440 0 0.00185748839124
Gc2_441 0 n4 ns441 0 0.00222410920186
Gc2_442 0 n4 ns442 0 0.000745956931016
Gc2_443 0 n4 ns443 0 0.00243420576994
Gc2_444 0 n4 ns444 0 5.46264004929e-05
Gc2_445 0 n4 ns445 0 0.00325226916723
Gc2_446 0 n4 ns446 0 0.000424212885871
Gc2_447 0 n4 ns447 0 -6.74321287756e-05
Gc2_448 0 n4 ns448 0 -2.66538111887e-05
Gd2_1 0 n4 ni1 0 0.00504122901047
Gd2_2 0 n4 ni2 0 -0.00579869172364
Gd2_3 0 n4 ni3 0 -0.00094960588339
Gd2_4 0 n4 ni4 0 0.00386358684348
Gd2_5 0 n4 ni5 0 -0.00011454735358
Gd2_6 0 n4 ni6 0 9.70893608501e-05
Gd2_7 0 n4 ni7 0 0.000200901114833
Gd2_8 0 n4 ni8 0 -0.000463495795991
Gc3_1 0 n6 ns1 0 0.0317479028697
Gc3_2 0 n6 ns2 0 -0.00566734190449
Gc3_3 0 n6 ns3 0 -0.000892772038531
Gc3_4 0 n6 ns4 0 0.00147228396924
Gc3_5 0 n6 ns5 0 -1.83923556145e-05
Gc3_6 0 n6 ns6 0 -3.0776451742e-05
Gc3_7 0 n6 ns7 0 -1.54179701041e-05
Gc3_8 0 n6 ns8 0 -2.64760823991e-05
Gc3_9 0 n6 ns9 0 2.43660798753e-07
Gc3_10 0 n6 ns10 0 2.18523857002e-07
Gc3_11 0 n6 ns11 0 -2.82772418145e-05
Gc3_12 0 n6 ns12 0 -0.000295720780004
Gc3_13 0 n6 ns13 0 -5.99674136074e-05
Gc3_14 0 n6 ns14 0 -0.000154048790259
Gc3_15 0 n6 ns15 0 -6.3462220745e-07
Gc3_16 0 n6 ns16 0 4.399243303e-08
Gc3_17 0 n6 ns17 0 -0.000326050945388
Gc3_18 0 n6 ns18 0 4.24605321567e-05
Gc3_19 0 n6 ns19 0 -0.000115200462827
Gc3_20 0 n6 ns20 0 8.47284381619e-05
Gc3_21 0 n6 ns21 0 2.652247751e-06
Gc3_22 0 n6 ns22 0 -2.39526879218e-06
Gc3_23 0 n6 ns23 0 0.000152180890715
Gc3_24 0 n6 ns24 0 -0.000387525498946
Gc3_25 0 n6 ns25 0 -4.07169103394e-05
Gc3_26 0 n6 ns26 0 -0.000212386259958
Gc3_27 0 n6 ns27 0 1.47517802874e-05
Gc3_28 0 n6 ns28 0 -4.45406843674e-05
Gc3_29 0 n6 ns29 0 -0.000314348238851
Gc3_30 0 n6 ns30 0 0.000686418103192
Gc3_31 0 n6 ns31 0 -0.000142379572055
Gc3_32 0 n6 ns32 0 -0.00016464304769
Gc3_33 0 n6 ns33 0 -0.00114106941741
Gc3_34 0 n6 ns34 0 7.48050643104e-06
Gc3_35 0 n6 ns35 0 0.000374363373931
Gc3_36 0 n6 ns36 0 0.000435375527264
Gc3_37 0 n6 ns37 0 -0.000741624447798
Gc3_38 0 n6 ns38 0 -1.6197792118e-05
Gc3_39 0 n6 ns39 0 -0.000249571326038
Gc3_40 0 n6 ns40 0 5.306410456e-05
Gc3_41 0 n6 ns41 0 -4.56677175149e-06
Gc3_42 0 n6 ns42 0 0.00264864650003
Gc3_43 0 n6 ns43 0 -0.00104079027009
Gc3_44 0 n6 ns44 0 -0.000249595157743
Gc3_45 0 n6 ns45 0 0.000169647856846
Gc3_46 0 n6 ns46 0 -0.000973664297
Gc3_47 0 n6 ns47 0 -1.17562562524e-05
Gc3_48 0 n6 ns48 0 -0.0020617039407
Gc3_49 0 n6 ns49 0 0.00104342761057
Gc3_50 0 n6 ns50 0 0.000181602407486
Gc3_51 0 n6 ns51 0 -0.00030566651504
Gc3_52 0 n6 ns52 0 -4.88012985773e-05
Gc3_53 0 n6 ns53 0 -0.000936713905129
Gc3_54 0 n6 ns54 0 -0.000165358155141
Gc3_55 0 n6 ns55 0 5.10585057075e-05
Gc3_56 0 n6 ns56 0 2.61912715295e-05
Gc3_57 0 n6 ns57 0 0.0226511000296
Gc3_58 0 n6 ns58 0 0.000257086904167
Gc3_59 0 n6 ns59 0 0.000313762208304
Gc3_60 0 n6 ns60 0 0.000212388476909
Gc3_61 0 n6 ns61 0 -1.13829077095e-05
Gc3_62 0 n6 ns62 0 -1.45292488164e-05
Gc3_63 0 n6 ns63 0 0.00011528843495
Gc3_64 0 n6 ns64 0 -8.79100076168e-05
Gc3_65 0 n6 ns65 0 -4.24090841631e-07
Gc3_66 0 n6 ns66 0 2.57571471813e-08
Gc3_67 0 n6 ns67 0 4.22394338045e-05
Gc3_68 0 n6 ns68 0 8.22030053124e-05
Gc3_69 0 n6 ns69 0 2.54686817037e-06
Gc3_70 0 n6 ns70 0 -0.000149724009724
Gc3_71 0 n6 ns71 0 -2.63862853588e-07
Gc3_72 0 n6 ns72 0 5.30879300257e-07
Gc3_73 0 n6 ns73 0 9.74670775006e-05
Gc3_74 0 n6 ns74 0 -6.65740701292e-05
Gc3_75 0 n6 ns75 0 -0.000161382347163
Gc3_76 0 n6 ns76 0 3.30399389121e-06
Gc3_77 0 n6 ns77 0 -4.64524242857e-06
Gc3_78 0 n6 ns78 0 1.74803628571e-06
Gc3_79 0 n6 ns79 0 1.86756469921e-05
Gc3_80 0 n6 ns80 0 0.000177720183388
Gc3_81 0 n6 ns81 0 0.000123322240312
Gc3_82 0 n6 ns82 0 -0.000129264425465
Gc3_83 0 n6 ns83 0 -3.02654075559e-05
Gc3_84 0 n6 ns84 0 2.21818659988e-05
Gc3_85 0 n6 ns85 0 -0.00020236895796
Gc3_86 0 n6 ns86 0 -0.00020089761583
Gc3_87 0 n6 ns87 0 2.48146361602e-05
Gc3_88 0 n6 ns88 0 -0.000297789096923
Gc3_89 0 n6 ns89 0 -6.06896035166e-07
Gc3_90 0 n6 ns90 0 -0.000476088692434
Gc3_91 0 n6 ns91 0 -4.14305239523e-05
Gc3_92 0 n6 ns92 0 0.000425639479038
Gc3_93 0 n6 ns93 0 1.27391410344e-05
Gc3_94 0 n6 ns94 0 -0.000324163236598
Gc3_95 0 n6 ns95 0 -0.000232881006592
Gc3_96 0 n6 ns96 0 9.17388339143e-05
Gc3_97 0 n6 ns97 0 -0.000928693493238
Gc3_98 0 n6 ns98 0 0.000293801154066
Gc3_99 0 n6 ns99 0 -0.000506815492062
Gc3_100 0 n6 ns100 0 -0.000610196731288
Gc3_101 0 n6 ns101 0 0.00105222718805
Gc3_102 0 n6 ns102 0 -0.000406724293967
Gc3_103 0 n6 ns103 0 0.00109166927642
Gc3_104 0 n6 ns104 0 -0.00151486373028
Gc3_105 0 n6 ns105 0 0.00122937078509
Gc3_106 0 n6 ns106 0 0.000287540507467
Gc3_107 0 n6 ns107 0 -0.000149053123068
Gc3_108 0 n6 ns108 0 -0.000657361944569
Gc3_109 0 n6 ns109 0 -0.000757133279405
Gc3_110 0 n6 ns110 0 -0.000454975098948
Gc3_111 0 n6 ns111 0 1.89400867473e-05
Gc3_112 0 n6 ns112 0 5.14290696961e-05
Gc3_113 0 n6 ns113 0 0.00373692429718
Gc3_114 0 n6 ns114 0 0.0104309678185
Gc3_115 0 n6 ns115 0 -0.00224997764108
Gc3_116 0 n6 ns116 0 -0.000725209441721
Gc3_117 0 n6 ns117 0 3.25280833094e-05
Gc3_118 0 n6 ns118 0 -4.27077748287e-06
Gc3_119 0 n6 ns119 0 0.00011495989905
Gc3_120 0 n6 ns120 0 4.05223000798e-05
Gc3_121 0 n6 ns121 0 5.47786109482e-07
Gc3_122 0 n6 ns122 0 -1.66722808931e-06
Gc3_123 0 n6 ns123 0 -6.70658171643e-05
Gc3_124 0 n6 ns124 0 -5.11542699068e-05
Gc3_125 0 n6 ns125 0 0.000201018232398
Gc3_126 0 n6 ns126 0 6.02700161672e-06
Gc3_127 0 n6 ns127 0 1.94547064219e-06
Gc3_128 0 n6 ns128 0 -1.8113440083e-06
Gc3_129 0 n6 ns129 0 -9.13136501336e-06
Gc3_130 0 n6 ns130 0 6.64976986729e-05
Gc3_131 0 n6 ns131 0 8.40732650539e-06
Gc3_132 0 n6 ns132 0 -0.000163465634067
Gc3_133 0 n6 ns133 0 4.42166631063e-06
Gc3_134 0 n6 ns134 0 3.76468360733e-06
Gc3_135 0 n6 ns135 0 -0.000102686468644
Gc3_136 0 n6 ns136 0 -1.65089988443e-05
Gc3_137 0 n6 ns137 0 9.907865917e-05
Gc3_138 0 n6 ns138 0 8.14202926101e-05
Gc3_139 0 n6 ns139 0 2.45097074449e-05
Gc3_140 0 n6 ns140 0 -3.81918954311e-06
Gc3_141 0 n6 ns141 0 3.16589684421e-05
Gc3_142 0 n6 ns142 0 -0.000154884541009
Gc3_143 0 n6 ns143 0 0.000168715592472
Gc3_144 0 n6 ns144 0 1.74351679377e-05
Gc3_145 0 n6 ns145 0 0.000203569784359
Gc3_146 0 n6 ns146 0 -5.68636278758e-05
Gc3_147 0 n6 ns147 0 -0.000354550736732
Gc3_148 0 n6 ns148 0 4.54067790335e-05
Gc3_149 0 n6 ns149 0 0.000218504410913
Gc3_150 0 n6 ns150 0 3.34743756058e-05
Gc3_151 0 n6 ns151 0 -0.000103736810434
Gc3_152 0 n6 ns152 0 -0.00033964050449
Gc3_153 0 n6 ns153 0 -0.000613866114946
Gc3_154 0 n6 ns154 0 -0.000330223507865
Gc3_155 0 n6 ns155 0 0.000894717373124
Gc3_156 0 n6 ns156 0 -0.000932479991433
Gc3_157 0 n6 ns157 0 0.000395292471778
Gc3_158 0 n6 ns158 0 0.000530845618145
Gc3_159 0 n6 ns159 0 0.00316039425092
Gc3_160 0 n6 ns160 0 0.000396786906155
Gc3_161 0 n6 ns161 0 -0.000469581579885
Gc3_162 0 n6 ns162 0 0.00379848357872
Gc3_163 0 n6 ns163 0 -0.00103677579744
Gc3_164 0 n6 ns164 0 -0.00156956111746
Gc3_165 0 n6 ns165 0 -0.0108286067483
Gc3_166 0 n6 ns166 0 -0.000579136972561
Gc3_167 0 n6 ns167 0 7.61037112245e-05
Gc3_168 0 n6 ns168 0 0.000129226954642
Gc3_169 0 n6 ns169 0 -0.00151417079328
Gc3_170 0 n6 ns170 0 -0.000697962221192
Gc3_171 0 n6 ns171 0 0.000556258472572
Gc3_172 0 n6 ns172 0 0.000735343334177
Gc3_173 0 n6 ns173 0 2.36105943475e-05
Gc3_174 0 n6 ns174 0 6.94392589934e-06
Gc3_175 0 n6 ns175 0 0.0001960705637
Gc3_176 0 n6 ns176 0 3.38734217303e-05
Gc3_177 0 n6 ns177 0 -8.99333170921e-07
Gc3_178 0 n6 ns178 0 1.17406784428e-06
Gc3_179 0 n6 ns179 0 6.86930281848e-06
Gc3_180 0 n6 ns180 0 0.000153113407445
Gc3_181 0 n6 ns181 0 0.000257900109149
Gc3_182 0 n6 ns182 0 -0.000132372024258
Gc3_183 0 n6 ns183 0 -1.88042514405e-06
Gc3_184 0 n6 ns184 0 -1.73776366917e-07
Gc3_185 0 n6 ns185 0 0.000163428431781
Gc3_186 0 n6 ns186 0 -2.59504983526e-05
Gc3_187 0 n6 ns187 0 -0.000173244064621
Gc3_188 0 n6 ns188 0 -0.000296671436484
Gc3_189 0 n6 ns189 0 2.41256714023e-06
Gc3_190 0 n6 ns190 0 -6.60852639822e-06
Gc3_191 0 n6 ns191 0 -5.99156205102e-05
Gc3_192 0 n6 ns192 0 0.000194045744801
Gc3_193 0 n6 ns193 0 0.000387891117562
Gc3_194 0 n6 ns194 0 0.000206981594434
Gc3_195 0 n6 ns195 0 -1.41440665311e-05
Gc3_196 0 n6 ns196 0 -4.83691482031e-05
Gc3_197 0 n6 ns197 0 4.20656760748e-05
Gc3_198 0 n6 ns198 0 -0.000267824882673
Gc3_199 0 n6 ns199 0 0.000542467282265
Gc3_200 0 n6 ns200 0 -0.000132294695172
Gc3_201 0 n6 ns201 0 0.000739504480832
Gc3_202 0 n6 ns202 0 -5.39134352701e-05
Gc3_203 0 n6 ns203 0 -0.000609253806495
Gc3_204 0 n6 ns204 0 0.000177873004846
Gc3_205 0 n6 ns205 0 0.00059429977289
Gc3_206 0 n6 ns206 0 -0.000193756589342
Gc3_207 0 n6 ns207 0 -0.000211802976589
Gc3_208 0 n6 ns208 0 -0.000250031926452
Gc3_209 0 n6 ns209 0 -0.00114700237612
Gc3_210 0 n6 ns210 0 -0.00101128818163
Gc3_211 0 n6 ns211 0 0.00046517534942
Gc3_212 0 n6 ns212 0 -0.00112171168389
Gc3_213 0 n6 ns213 0 0.00103002716728
Gc3_214 0 n6 ns214 0 0.000651035177163
Gc3_215 0 n6 ns215 0 0.00272654189809
Gc3_216 0 n6 ns216 0 -3.06080290101e-05
Gc3_217 0 n6 ns217 0 0.000626997896911
Gc3_218 0 n6 ns218 0 0.00241232161918
Gc3_219 0 n6 ns219 0 -0.000142921554989
Gc3_220 0 n6 ns220 0 -0.00226438738646
Gc3_221 0 n6 ns221 0 -0.00679025774075
Gc3_222 0 n6 ns222 0 -0.0006523431283
Gc3_223 0 n6 ns223 0 4.3452301513e-05
Gc3_224 0 n6 ns224 0 0.000114964428917
Gc3_225 0 n6 ns225 0 0.00410510135887
Gc3_226 0 n6 ns226 0 7.3969538696e-05
Gc3_227 0 n6 ns227 0 -0.00019290859757
Gc3_228 0 n6 ns228 0 -0.000281569058017
Gc3_229 0 n6 ns229 0 1.15492434246e-05
Gc3_230 0 n6 ns230 0 2.80588641744e-05
Gc3_231 0 n6 ns231 0 4.6595664315e-05
Gc3_232 0 n6 ns232 0 3.30220489974e-05
Gc3_233 0 n6 ns233 0 -1.3975964515e-07
Gc3_234 0 n6 ns234 0 -2.3262570258e-07
Gc3_235 0 n6 ns235 0 8.17838412287e-06
Gc3_236 0 n6 ns236 0 -0.000267802019846
Gc3_237 0 n6 ns237 0 -9.08757557896e-05
Gc3_238 0 n6 ns238 0 -0.000114995905624
Gc3_239 0 n6 ns239 0 9.5356114839e-07
Gc3_240 0 n6 ns240 0 1.65870318137e-07
Gc3_241 0 n6 ns241 0 0.000297755114514
Gc3_242 0 n6 ns242 0 -3.40126065225e-05
Gc3_243 0 n6 ns243 0 0.000128552465434
Gc3_244 0 n6 ns244 0 -0.000124974548348
Gc3_245 0 n6 ns245 0 1.84337627927e-07
Gc3_246 0 n6 ns246 0 -3.70047216758e-06
Gc3_247 0 n6 ns247 0 0.000179930060709
Gc3_248 0 n6 ns248 0 -0.000433279568062
Gc3_249 0 n6 ns249 0 2.60079022374e-05
Gc3_250 0 n6 ns250 0 -0.000219770581139
Gc3_251 0 n6 ns251 0 -1.92004208708e-06
Gc3_252 0 n6 ns252 0 1.02552947113e-05
Gc3_253 0 n6 ns253 0 -1.09656867224e-06
Gc3_254 0 n6 ns254 0 -0.000836228769261
Gc3_255 0 n6 ns255 0 0.000157977811689
Gc3_256 0 n6 ns256 0 0.000415009388453
Gc3_257 0 n6 ns257 0 -0.00161092369213
Gc3_258 0 n6 ns258 0 -0.000276259389037
Gc3_259 0 n6 ns259 0 0.000142057201303
Gc3_260 0 n6 ns260 0 0.000547163940317
Gc3_261 0 n6 ns261 0 0.000525890716072
Gc3_262 0 n6 ns262 0 0.000189087903116
Gc3_263 0 n6 ns263 0 0.00037248349481
Gc3_264 0 n6 ns264 0 -0.00019529708323
Gc3_265 0 n6 ns265 0 -0.000740118891355
Gc3_266 0 n6 ns266 0 0.00224474161192
Gc3_267 0 n6 ns267 0 -0.0007983471612
Gc3_268 0 n6 ns268 0 -0.000247464251814
Gc3_269 0 n6 ns269 0 -0.00181778507417
Gc3_270 0 n6 ns270 0 0.00180957900411
Gc3_271 0 n6 ns271 0 -0.00120937830192
Gc3_272 0 n6 ns272 0 0.00117387848649
Gc3_273 0 n6 ns273 0 0.00145363986381
Gc3_274 0 n6 ns274 0 -0.0004416158869
Gc3_275 0 n6 ns275 0 0.0015204812495
Gc3_276 0 n6 ns276 0 -0.000929480864747
Gc3_277 0 n6 ns277 0 0.00176545951587
Gc3_278 0 n6 ns278 0 0.000106015269171
Gc3_279 0 n6 ns279 0 -4.38083463129e-05
Gc3_280 0 n6 ns280 0 2.94829197676e-05
Gc3_281 0 n6 ns281 0 -0.000744609710124
Gc3_282 0 n6 ns282 0 -0.000221942877758
Gc3_283 0 n6 ns283 0 0.000254143727077
Gc3_284 0 n6 ns284 0 0.000131767220451
Gc3_285 0 n6 ns285 0 -2.34133356283e-07
Gc3_286 0 n6 ns286 0 1.61555249505e-05
Gc3_287 0 n6 ns287 0 -3.38837347592e-05
Gc3_288 0 n6 ns288 0 7.3173069037e-05
Gc3_289 0 n6 ns289 0 6.05665433097e-08
Gc3_290 0 n6 ns290 0 1.64268013503e-07
Gc3_291 0 n6 ns291 0 6.48773851753e-05
Gc3_292 0 n6 ns292 0 0.000125412987009
Gc3_293 0 n6 ns293 0 -5.18517650484e-05
Gc3_294 0 n6 ns294 0 -8.99372189604e-05
Gc3_295 0 n6 ns295 0 2.09684289225e-08
Gc3_296 0 n6 ns296 0 -1.35468678061e-06
Gc3_297 0 n6 ns297 0 -9.23891994221e-05
Gc3_298 0 n6 ns298 0 9.76948590841e-05
Gc3_299 0 n6 ns299 0 0.000122173222444
Gc3_300 0 n6 ns300 0 -3.97925229361e-05
Gc3_301 0 n6 ns301 0 -6.65168337042e-06
Gc3_302 0 n6 ns302 0 3.32496086694e-06
Gc3_303 0 n6 ns303 0 1.31117103296e-05
Gc3_304 0 n6 ns304 0 0.000195720718001
Gc3_305 0 n6 ns305 0 9.64964821342e-05
Gc3_306 0 n6 ns306 0 -0.000208540854653
Gc3_307 0 n6 ns307 0 2.74966816749e-05
Gc3_308 0 n6 ns308 0 -3.79026214347e-05
Gc3_309 0 n6 ns309 0 0.000242233071514
Gc3_310 0 n6 ns310 0 0.000158984234294
Gc3_311 0 n6 ns311 0 2.71568817319e-05
Gc3_312 0 n6 ns312 0 0.000130630970069
Gc3_313 0 n6 ns313 0 0.000115271769661
Gc3_314 0 n6 ns314 0 -0.000695990683216
Gc3_315 0 n6 ns315 0 0.000118540961526
Gc3_316 0 n6 ns316 0 0.000188401469348
Gc3_317 0 n6 ns317 0 1.89381826262e-05
Gc3_318 0 n6 ns318 0 0.000366009951109
Gc3_319 0 n6 ns319 0 0.000188898903766
Gc3_320 0 n6 ns320 0 -0.000143078274145
Gc3_321 0 n6 ns321 0 -0.00110509121193
Gc3_322 0 n6 ns322 0 1.68219996356e-05
Gc3_323 0 n6 ns323 0 -0.000646017227225
Gc3_324 0 n6 ns324 0 -0.000330924917501
Gc3_325 0 n6 ns325 0 -0.00128293229304
Gc3_326 0 n6 ns326 0 0.000171007611578
Gc3_327 0 n6 ns327 0 -0.000536781175482
Gc3_328 0 n6 ns328 0 0.000867140540097
Gc3_329 0 n6 ns329 0 0.0014230201684
Gc3_330 0 n6 ns330 0 4.26201314088e-06
Gc3_331 0 n6 ns331 0 0.00110437369521
Gc3_332 0 n6 ns332 0 -0.000246138919909
Gc3_333 0 n6 ns333 0 0.00104592081712
Gc3_334 0 n6 ns334 0 0.000374585052266
Gc3_335 0 n6 ns335 0 -3.40886216981e-05
Gc3_336 0 n6 ns336 0 -1.75484541594e-05
Gc3_337 0 n6 ns337 0 -0.00964328212767
Gc3_338 0 n6 ns338 0 0.000616984077227
Gc3_339 0 n6 ns339 0 -0.000189965886386
Gc3_340 0 n6 ns340 0 -0.000279534003263
Gc3_341 0 n6 ns341 0 -2.28295057602e-05
Gc3_342 0 n6 ns342 0 -1.39628248234e-05
Gc3_343 0 n6 ns343 0 -0.00025867423096
Gc3_344 0 n6 ns344 0 -5.47103609482e-05
Gc3_345 0 n6 ns345 0 8.72757624025e-07
Gc3_346 0 n6 ns346 0 -5.0404788795e-07
Gc3_347 0 n6 ns347 0 -8.58858836365e-05
Gc3_348 0 n6 ns348 0 -0.000165106711224
Gc3_349 0 n6 ns349 0 0.000309708866005
Gc3_350 0 n6 ns350 0 -0.000107831623835
Gc3_351 0 n6 ns351 0 -2.0311366627e-06
Gc3_352 0 n6 ns352 0 -2.94443479633e-07
Gc3_353 0 n6 ns353 0 0.000157747179865
Gc3_354 0 n6 ns354 0 -0.00012446182061
Gc3_355 0 n6 ns355 0 0.000114040575641
Gc3_356 0 n6 ns356 0 0.000340895817788
Gc3_357 0 n6 ns357 0 -4.24926324953e-07
Gc3_358 0 n6 ns358 0 5.58894783552e-06
Gc3_359 0 n6 ns359 0 -8.58525019991e-05
Gc3_360 0 n6 ns360 0 -0.000285082680114
Gc3_361 0 n6 ns361 0 0.000324508674464
Gc3_362 0 n6 ns362 0 0.000267276362427
Gc3_363 0 n6 ns363 0 -1.58872569382e-05
Gc3_364 0 n6 ns364 0 -3.94181488823e-05
Gc3_365 0 n6 ns365 0 -0.00030510857131
Gc3_366 0 n6 ns366 0 -0.000372558300297
Gc3_367 0 n6 ns367 0 -0.000523914068529
Gc3_368 0 n6 ns368 0 1.91833437566e-05
Gc3_369 0 n6 ns369 0 -0.000778196499484
Gc3_370 0 n6 ns370 0 0.000589706953457
Gc3_371 0 n6 ns371 0 -0.000658673185971
Gc3_372 0 n6 ns372 0 0.000177080979484
Gc3_373 0 n6 ns373 0 0.000114066008977
Gc3_374 0 n6 ns374 0 -0.000386822201645
Gc3_375 0 n6 ns375 0 1.84951328068e-05
Gc3_376 0 n6 ns376 0 0.000573520879254
Gc3_377 0 n6 ns377 0 0.00335480781024
Gc3_378 0 n6 ns378 0 0.00124640705995
Gc3_379 0 n6 ns379 0 0.00138917954411
Gc3_380 0 n6 ns380 0 -0.000917502511127
Gc3_381 0 n6 ns381 0 0.0013208013287
Gc3_382 0 n6 ns382 0 0.0025818054778
Gc3_383 0 n6 ns383 0 -0.00614875071515
Gc3_384 0 n6 ns384 0 0.000904394324435
Gc3_385 0 n6 ns385 0 -0.0018607431316
Gc3_386 0 n6 ns386 0 0.00569710243156
Gc3_387 0 n6 ns387 0 -0.00437945528506
Gc3_388 0 n6 ns388 0 -0.00320897043094
Gc3_389 0 n6 ns389 0 0.0207073680994
Gc3_390 0 n6 ns390 0 -0.000329721319082
Gc3_391 0 n6 ns391 0 8.29591946493e-05
Gc3_392 0 n6 ns392 0 -3.25718074814e-05
Gc3_393 0 n6 ns393 0 -0.0126566006478
Gc3_394 0 n6 ns394 0 0.000586997496841
Gc3_395 0 n6 ns395 0 0.000327553614719
Gc3_396 0 n6 ns396 0 0.000240920609566
Gc3_397 0 n6 ns397 0 -2.12322738502e-05
Gc3_398 0 n6 ns398 0 -9.96990202595e-06
Gc3_399 0 n6 ns399 0 -0.000273596129753
Gc3_400 0 n6 ns400 0 2.85380691599e-06
Gc3_401 0 n6 ns401 0 -1.43453324702e-06
Gc3_402 0 n6 ns402 0 4.95037844977e-07
Gc3_403 0 n6 ns403 0 9.44027352426e-06
Gc3_404 0 n6 ns404 0 0.000207248455771
Gc3_405 0 n6 ns405 0 0.00023730907337
Gc3_406 0 n6 ns406 0 -9.86420859385e-05
Gc3_407 0 n6 ns407 0 3.12230118492e-06
Gc3_408 0 n6 ns408 0 1.77772912503e-06
Gc3_409 0 n6 ns409 0 -0.000192483159488
Gc3_410 0 n6 ns410 0 5.47183962957e-05
Gc3_411 0 n6 ns411 0 0.000120098600563
Gc3_412 0 n6 ns412 0 0.000290141003423
Gc3_413 0 n6 ns413 0 6.18550416153e-06
Gc3_414 0 n6 ns414 0 -5.31318542618e-06
Gc3_415 0 n6 ns415 0 -0.000171641058333
Gc3_416 0 n6 ns416 0 0.000289877909632
Gc3_417 0 n6 ns417 0 0.000328237147678
Gc3_418 0 n6 ns418 0 0.000103471738914
Gc3_419 0 n6 ns419 0 -2.09895331638e-05
Gc3_420 0 n6 ns420 0 4.47168728931e-05
Gc3_421 0 n6 ns421 0 -4.43899468011e-05
Gc3_422 0 n6 ns422 0 0.000650293502006
Gc3_423 0 n6 ns423 0 -0.000317707247831
Gc3_424 0 n6 ns424 0 0.000207694523773
Gc3_425 0 n6 ns425 0 0.00172441553884
Gc3_426 0 n6 ns426 0 0.000681501882247
Gc3_427 0 n6 ns427 0 -0.000142087144764
Gc3_428 0 n6 ns428 0 0.000363356470122
Gc3_429 0 n6 ns429 0 -0.000712648182408
Gc3_430 0 n6 ns430 0 -4.23009151186e-05
Gc3_431 0 n6 ns431 0 0.000336183035942
Gc3_432 0 n6 ns432 0 0.000236907864815
Gc3_433 0 n6 ns433 0 0.00121554820999
Gc3_434 0 n6 ns434 0 -0.00412069835299
Gc3_435 0 n6 ns435 0 -0.000131526255853
Gc3_436 0 n6 ns436 0 -0.00114412588298
Gc3_437 0 n6 ns437 0 0.000863824995891
Gc3_438 0 n6 ns438 0 -0.00245891174019
Gc3_439 0 n6 ns439 0 -5.23830089881e-05
Gc3_440 0 n6 ns440 0 0.00126700227254
Gc3_441 0 n6 ns441 0 0.00232120905747
Gc3_442 0 n6 ns442 0 0.00205978124251
Gc3_443 0 n6 ns443 0 0.00321703108478
Gc3_444 0 n6 ns444 0 0.00155704078977
Gc3_445 0 n6 ns445 0 0.00445724973979
Gc3_446 0 n6 ns446 0 0.000608646054085
Gc3_447 0 n6 ns447 0 -9.13339975696e-05
Gc3_448 0 n6 ns448 0 -0.000102759760671
Gd3_1 0 n6 ni1 0 0.0031446494216
Gd3_2 0 n6 ni2 0 -0.00094960557205
Gd3_3 0 n6 ni3 0 -0.00409572811548
Gd3_4 0 n6 ni4 0 0.00503106820494
Gd3_5 0 n6 ni5 0 -0.000178702702493
Gd3_6 0 n6 ni6 0 0.000201935278305
Gd3_7 0 n6 ni7 0 -0.0004692420671
Gd3_8 0 n6 ni8 0 -0.000112621536783
Gc4_1 0 n8 ns1 0 0.0227101318636
Gc4_2 0 n8 ns2 0 0.000253011012983
Gc4_3 0 n8 ns3 0 0.0003135575652
Gc4_4 0 n8 ns4 0 0.000213661932854
Gc4_5 0 n8 ns5 0 -1.14418764808e-05
Gc4_6 0 n8 ns6 0 -1.45606077137e-05
Gc4_7 0 n8 ns7 0 0.000115321861736
Gc4_8 0 n8 ns8 0 -8.80102669003e-05
Gc4_9 0 n8 ns9 0 -4.30865212088e-07
Gc4_10 0 n8 ns10 0 1.16642238771e-08
Gc4_11 0 n8 ns11 0 4.19951658733e-05
Gc4_12 0 n8 ns12 0 8.1893926122e-05
Gc4_13 0 n8 ns13 0 2.28892342917e-06
Gc4_14 0 n8 ns14 0 -0.000149816195682
Gc4_15 0 n8 ns15 0 -2.64522626742e-07
Gc4_16 0 n8 ns16 0 5.06227165593e-07
Gc4_17 0 n8 ns17 0 9.71812185653e-05
Gc4_18 0 n8 ns18 0 -6.63307633139e-05
Gc4_19 0 n8 ns19 0 -0.000161371054954
Gc4_20 0 n8 ns20 0 3.56484092106e-06
Gc4_21 0 n8 ns21 0 -4.59885760393e-06
Gc4_22 0 n8 ns22 0 1.73188021946e-06
Gc4_23 0 n8 ns23 0 1.85812594092e-05
Gc4_24 0 n8 ns24 0 0.000177316878704
Gc4_25 0 n8 ns25 0 0.000122946823996
Gc4_26 0 n8 ns26 0 -0.000129442402521
Gc4_27 0 n8 ns27 0 -3.02354609821e-05
Gc4_28 0 n8 ns28 0 2.20076202884e-05
Gc4_29 0 n8 ns29 0 -0.000202227864763
Gc4_30 0 n8 ns30 0 -0.000199884683367
Gc4_31 0 n8 ns31 0 2.45910322845e-05
Gc4_32 0 n8 ns32 0 -0.000297659889606
Gc4_33 0 n8 ns33 0 -1.9018945464e-06
Gc4_34 0 n8 ns34 0 -0.000474810449561
Gc4_35 0 n8 ns35 0 -4.05733769573e-05
Gc4_36 0 n8 ns36 0 0.000425670236189
Gc4_37 0 n8 ns37 0 1.22304617138e-05
Gc4_38 0 n8 ns38 0 -0.000323475937931
Gc4_39 0 n8 ns39 0 -0.000233078235956
Gc4_40 0 n8 ns40 0 9.21153199121e-05
Gc4_41 0 n8 ns41 0 -0.000926550089983
Gc4_42 0 n8 ns42 0 0.000295376036542
Gc4_43 0 n8 ns43 0 -0.000507825527223
Gc4_44 0 n8 ns44 0 -0.000609505424179
Gc4_45 0 n8 ns45 0 0.00105144782031
Gc4_46 0 n8 ns46 0 -0.000407404285693
Gc4_47 0 n8 ns47 0 0.00108990687288
Gc4_48 0 n8 ns48 0 -0.0015159536295
Gc4_49 0 n8 ns49 0 0.00123153762793
Gc4_50 0 n8 ns50 0 0.000287152042038
Gc4_51 0 n8 ns51 0 -0.000146936614883
Gc4_52 0 n8 ns52 0 -0.000658272265039
Gc4_53 0 n8 ns53 0 -0.000754507342461
Gc4_54 0 n8 ns54 0 -0.000455180540327
Gc4_55 0 n8 ns55 0 1.89354855675e-05
Gc4_56 0 n8 ns56 0 5.15132310081e-05
Gc4_57 0 n8 ns57 0 0.0162264344444
Gc4_58 0 n8 ns58 0 -0.00290422969929
Gc4_59 0 n8 ns59 0 -0.000318652515915
Gc4_60 0 n8 ns60 0 0.00100347340305
Gc4_61 0 n8 ns61 0 2.90756085539e-08
Gc4_62 0 n8 ns62 0 -9.726249304e-06
Gc4_63 0 n8 ns63 0 0.00011516746553
Gc4_64 0 n8 ns64 0 -9.78229580327e-06
Gc4_65 0 n8 ns65 0 -3.20048355044e-06
Gc4_66 0 n8 ns66 0 -2.35903429303e-06
Gc4_67 0 n8 ns67 0 -1.371421395e-05
Gc4_68 0 n8 ns68 0 -0.000156416884585
Gc4_69 0 n8 ns69 0 8.22806970943e-05
Gc4_70 0 n8 ns70 0 -0.000161815741678
Gc4_71 0 n8 ns71 0 -2.51948719634e-06
Gc4_72 0 n8 ns72 0 -7.0599617168e-06
Gc4_73 0 n8 ns73 0 -0.000163901841933
Gc4_74 0 n8 ns74 0 1.91968900249e-05
Gc4_75 0 n8 ns75 0 -0.000152775939133
Gc4_76 0 n8 ns76 0 -8.09308291563e-05
Gc4_77 0 n8 ns77 0 2.01844226893e-05
Gc4_78 0 n8 ns78 0 -9.65579925006e-06
Gc4_79 0 n8 ns79 0 8.76438490263e-05
Gc4_80 0 n8 ns80 0 -0.000192367160387
Gc4_81 0 n8 ns81 0 0.00015993900179
Gc4_82 0 n8 ns82 0 -1.66153561235e-05
Gc4_83 0 n8 ns83 0 4.30532590222e-05
Gc4_84 0 n8 ns84 0 -0.000102198365909
Gc4_85 0 n8 ns85 0 -0.000148627507209
Gc4_86 0 n8 ns86 0 0.000448250021043
Gc4_87 0 n8 ns87 0 0.000158097600541
Gc4_88 0 n8 ns88 0 -9.86573443349e-05
Gc4_89 0 n8 ns89 0 -0.000318064755953
Gc4_90 0 n8 ns90 0 0.000123271675326
Gc4_91 0 n8 ns91 0 -1.38522522114e-05
Gc4_92 0 n8 ns92 0 0.000313161661417
Gc4_93 0 n8 ns93 0 -6.37495707719e-05
Gc4_94 0 n8 ns94 0 -9.04993690184e-05
Gc4_95 0 n8 ns95 0 -0.000303356372425
Gc4_96 0 n8 ns96 0 -3.02018654587e-05
Gc4_97 0 n8 ns97 0 -0.000486258416681
Gc4_98 0 n8 ns98 0 0.000714345713751
Gc4_99 0 n8 ns99 0 -0.000439979387418
Gc4_100 0 n8 ns100 0 -0.000774917800471
Gc4_101 0 n8 ns101 0 0.000871600729612
Gc4_102 0 n8 ns102 0 -6.54687534037e-05
Gc4_103 0 n8 ns103 0 0.00150258661733
Gc4_104 0 n8 ns104 0 -0.00125655883432
Gc4_105 0 n8 ns105 0 0.00114353280163
Gc4_106 0 n8 ns106 0 0.00115299915373
Gc4_107 0 n8 ns107 0 -0.000214333871249
Gc4_108 0 n8 ns108 0 -0.00129387962517
Gc4_109 0 n8 ns109 0 -0.00352639960762
Gc4_110 0 n8 ns110 0 -0.000541182587825
Gc4_111 0 n8 ns111 0 4.33962441703e-05
Gc4_112 0 n8 ns112 0 7.30319719783e-05
Gc4_113 0 n8 ns113 0 -0.00151424382074
Gc4_114 0 n8 ns114 0 -0.000697953534209
Gc4_115 0 n8 ns115 0 0.000556260324936
Gc4_116 0 n8 ns116 0 0.000735343025591
Gc4_117 0 n8 ns117 0 2.36105807147e-05
Gc4_118 0 n8 ns118 0 6.94390764341e-06
Gc4_119 0 n8 ns119 0 0.000196070632629
Gc4_120 0 n8 ns120 0 3.38734595412e-05
Gc4_121 0 n8 ns121 0 -8.99327203021e-07
Gc4_122 0 n8 ns122 0 1.17407168797e-06
Gc4_123 0 n8 ns123 0 6.86910459145e-06
Gc4_124 0 n8 ns124 0 0.000153113528696
Gc4_125 0 n8 ns125 0 0.000257899775244
Gc4_126 0 n8 ns126 0 -0.000132372110605
Gc4_127 0 n8 ns127 0 -1.88042082421e-06
Gc4_128 0 n8 ns128 0 -1.73794841047e-07
Gc4_129 0 n8 ns129 0 0.000163428317231
Gc4_130 0 n8 ns130 0 -2.5950606232e-05
Gc4_131 0 n8 ns131 0 -0.000173244518881
Gc4_132 0 n8 ns132 0 -0.000296671235969
Gc4_133 0 n8 ns133 0 2.41256328885e-06
Gc4_134 0 n8 ns134 0 -6.60850058614e-06
Gc4_135 0 n8 ns135 0 -5.99165954745e-05
Gc4_136 0 n8 ns136 0 0.000194046314625
Gc4_137 0 n8 ns137 0 0.000387890700629
Gc4_138 0 n8 ns138 0 0.000206981282043
Gc4_139 0 n8 ns139 0 -1.41440370322e-05
Gc4_140 0 n8 ns140 0 -4.83692449897e-05
Gc4_141 0 n8 ns141 0 4.20659535106e-05
Gc4_142 0 n8 ns142 0 -0.000267824995
Gc4_143 0 n8 ns143 0 0.000542466937398
Gc4_144 0 n8 ns144 0 -0.000132295020812
Gc4_145 0 n8 ns145 0 0.000739508576982
Gc4_146 0 n8 ns146 0 -5.3911914796e-05
Gc4_147 0 n8 ns147 0 -0.00060925388824
Gc4_148 0 n8 ns148 0 0.000177869535861
Gc4_149 0 n8 ns149 0 0.000594299331422
Gc4_150 0 n8 ns150 0 -0.000193757451454
Gc4_151 0 n8 ns151 0 -0.000211803561125
Gc4_152 0 n8 ns152 0 -0.000250032513984
Gc4_153 0 n8 ns153 0 -0.00114700039649
Gc4_154 0 n8 ns154 0 -0.0010112958595
Gc4_155 0 n8 ns155 0 0.000465179978233
Gc4_156 0 n8 ns156 0 -0.00112170885837
Gc4_157 0 n8 ns157 0 0.00103003046327
Gc4_158 0 n8 ns158 0 0.000651029265827
Gc4_159 0 n8 ns159 0 0.00272654583998
Gc4_160 0 n8 ns160 0 -3.06103345286e-05
Gc4_161 0 n8 ns161 0 0.000626996620388
Gc4_162 0 n8 ns162 0 0.00241232522757
Gc4_163 0 n8 ns163 0 -0.000142919182402
Gc4_164 0 n8 ns164 0 -0.00226438477286
Gc4_165 0 n8 ns165 0 -0.00679025607165
Gc4_166 0 n8 ns166 0 -0.000652343116194
Gc4_167 0 n8 ns167 0 4.34521839444e-05
Gc4_168 0 n8 ns168 0 0.000114964120042
Gc4_169 0 n8 ns169 0 0.0151634279623
Gc4_170 0 n8 ns170 0 0.010234756782
Gc4_171 0 n8 ns171 0 -0.00245737654202
Gc4_172 0 n8 ns172 0 -0.000975525601021
Gc4_173 0 n8 ns173 0 2.24609968187e-05
Gc4_174 0 n8 ns174 0 -1.32323715467e-05
Gc4_175 0 n8 ns175 0 0.000179850489456
Gc4_176 0 n8 ns176 0 -9.18334506042e-06
Gc4_177 0 n8 ns177 0 3.78157162736e-06
Gc4_178 0 n8 ns178 0 1.39514496494e-06
Gc4_179 0 n8 ns179 0 -1.97530172242e-05
Gc4_180 0 n8 ns180 0 -4.98507775305e-05
Gc4_181 0 n8 ns181 0 0.000177924366119
Gc4_182 0 n8 ns182 0 -7.21432584296e-05
Gc4_183 0 n8 ns183 0 3.71721695426e-06
Gc4_184 0 n8 ns184 0 5.1323757819e-06
Gc4_185 0 n8 ns185 0 1.88769517477e-05
Gc4_186 0 n8 ns186 0 2.4742586137e-06
Gc4_187 0 n8 ns187 0 -6.82351952667e-05
Gc4_188 0 n8 ns188 0 -0.000113863923462
Gc4_189 0 n8 ns189 0 -1.29640536682e-05
Gc4_190 0 n8 ns190 0 1.05879453708e-05
Gc4_191 0 n8 ns191 0 -4.59366296775e-05
Gc4_192 0 n8 ns192 0 8.9784875089e-05
Gc4_193 0 n8 ns193 0 0.000111693974003
Gc4_194 0 n8 ns194 0 -6.19522973093e-05
Gc4_195 0 n8 ns195 0 -2.38789561638e-05
Gc4_196 0 n8 ns196 0 5.25691333625e-05
Gc4_197 0 n8 ns197 0 -0.000208448048154
Gc4_198 0 n8 ns198 0 -0.000316947574846
Gc4_199 0 n8 ns199 0 0.000100943393943
Gc4_200 0 n8 ns200 0 -0.000233073367421
Gc4_201 0 n8 ns201 0 6.45060067958e-06
Gc4_202 0 n8 ns202 0 -0.000577616987129
Gc4_203 0 n8 ns203 0 -0.000286565401002
Gc4_204 0 n8 ns204 0 0.000396992956852
Gc4_205 0 n8 ns205 0 2.0905914986e-05
Gc4_206 0 n8 ns206 0 -0.000224338521027
Gc4_207 0 n8 ns207 0 -0.000238467857843
Gc4_208 0 n8 ns208 0 -0.000203364218765
Gc4_209 0 n8 ns209 0 -0.00109570839164
Gc4_210 0 n8 ns210 0 0.000256784476193
Gc4_211 0 n8 ns211 0 0.00034259494099
Gc4_212 0 n8 ns212 0 -0.000989533056065
Gc4_213 0 n8 ns213 0 0.000843707682719
Gc4_214 0 n8 ns214 0 -1.16474537791e-05
Gc4_215 0 n8 ns215 0 0.00305494055246
Gc4_216 0 n8 ns216 0 -0.000487138367901
Gc4_217 0 n8 ns217 0 -0.000123319413932
Gc4_218 0 n8 ns218 0 0.00326997228839
Gc4_219 0 n8 ns219 0 -0.00134672056687
Gc4_220 0 n8 ns220 0 -0.00157170984538
Gc4_221 0 n8 ns221 0 -0.0100645358981
Gc4_222 0 n8 ns222 0 -0.000505654385536
Gc4_223 0 n8 ns223 0 6.29475844042e-05
Gc4_224 0 n8 ns224 0 6.70543164478e-05
Gc4_225 0 n8 ns225 0 -0.000708894526681
Gc4_226 0 n8 ns226 0 -0.000224475827098
Gc4_227 0 n8 ns227 0 0.00025369853231
Gc4_228 0 n8 ns228 0 0.000131827738436
Gc4_229 0 n8 ns229 0 -2.08121250869e-07
Gc4_230 0 n8 ns230 0 1.61934168378e-05
Gc4_231 0 n8 ns231 0 -3.36132187691e-05
Gc4_232 0 n8 ns232 0 7.33014568589e-05
Gc4_233 0 n8 ns233 0 5.54538485213e-08
Gc4_234 0 n8 ns234 0 1.50840203996e-07
Gc4_235 0 n8 ns235 0 6.47128421529e-05
Gc4_236 0 n8 ns236 0 0.000124941788216
Gc4_237 0 n8 ns237 0 -5.22044752347e-05
Gc4_238 0 n8 ns238 0 -9.00405224047e-05
Gc4_239 0 n8 ns239 0 1.68565007363e-08
Gc4_240 0 n8 ns240 0 -1.33182630332e-06
Gc4_241 0 n8 ns241 0 -9.20280336089e-05
Gc4_242 0 n8 ns242 0 9.74245872126e-05
Gc4_243 0 n8 ns243 0 0.000122229637905
Gc4_244 0 n8 ns244 0 -4.03012271727e-05
Gc4_245 0 n8 ns245 0 -6.59933411794e-06
Gc4_246 0 n8 ns246 0 3.316531435e-06
Gc4_247 0 n8 ns247 0 1.31782059434e-05
Gc4_248 0 n8 ns248 0 0.000194952911739
Gc4_249 0 n8 ns249 0 9.62410655955e-05
Gc4_250 0 n8 ns250 0 -0.00020894776529
Gc4_251 0 n8 ns251 0 2.73410916545e-05
Gc4_252 0 n8 ns252 0 -3.77877414338e-05
Gc4_253 0 n8 ns253 0 0.000241459034277
Gc4_254 0 n8 ns254 0 0.000157933508313
Gc4_255 0 n8 ns255 0 2.79452339674e-05
Gc4_256 0 n8 ns256 0 0.000131271368973
Gc4_257 0 n8 ns257 0 0.000111932828728
Gc4_258 0 n8 ns258 0 -0.000695062644553
Gc4_259 0 n8 ns259 0 0.000119479903172
Gc4_260 0 n8 ns260 0 0.000189396695873
Gc4_261 0 n8 ns261 0 1.95644254284e-05
Gc4_262 0 n8 ns262 0 0.000366255634277
Gc4_263 0 n8 ns263 0 0.000188933310156
Gc4_264 0 n8 ns264 0 -0.000143746700816
Gc4_265 0 n8 ns265 0 -0.00110359448234
Gc4_266 0 n8 ns266 0 2.02146992836e-05
Gc4_267 0 n8 ns267 0 -0.00064673487396
Gc4_268 0 n8 ns268 0 -0.000330557653813
Gc4_269 0 n8 ns269 0 -0.00128330334318
Gc4_270 0 n8 ns270 0 0.00017128916257
Gc4_271 0 n8 ns271 0 -0.000536079649145
Gc4_272 0 n8 ns272 0 0.000866501464525
Gc4_273 0 n8 ns273 0 0.00142573956536
Gc4_274 0 n8 ns274 0 6.10479764742e-06
Gc4_275 0 n8 ns275 0 0.0011064066382
Gc4_276 0 n8 ns276 0 -0.000246874555416
Gc4_277 0 n8 ns277 0 0.00104585575934
Gc4_278 0 n8 ns278 0 0.000374733817435
Gc4_279 0 n8 ns279 0 -3.40616999901e-05
Gc4_280 0 n8 ns280 0 -1.74767218818e-05
Gc4_281 0 n8 ns281 0 -0.0029539134103
Gc4_282 0 n8 ns282 0 0.000696611049231
Gc4_283 0 n8 ns283 0 -7.5916833728e-05
Gc4_284 0 n8 ns284 0 -0.000153142199937
Gc4_285 0 n8 ns285 0 -2.51989248371e-06
Gc4_286 0 n8 ns286 0 1.67253380431e-05
Gc4_287 0 n8 ns287 0 -0.000108936621965
Gc4_288 0 n8 ns288 0 3.3906841265e-05
Gc4_289 0 n8 ns289 0 -4.42013475677e-06
Gc4_290 0 n8 ns290 0 -4.11858102997e-06
Gc4_291 0 n8 ns291 0 1.90872022396e-06
Gc4_292 0 n8 ns292 0 -0.000183525099472
Gc4_293 0 n8 ns293 0 6.06579088173e-05
Gc4_294 0 n8 ns294 0 -0.000176032921024
Gc4_295 0 n8 ns295 0 4.35319449641e-06
Gc4_296 0 n8 ns296 0 1.09130789511e-05
Gc4_297 0 n8 ns297 0 0.000198103190356
Gc4_298 0 n8 ns298 0 -2.39923572126e-05
Gc4_299 0 n8 ns299 0 0.000192573930584
Gc4_300 0 n8 ns300 0 4.62870829617e-05
Gc4_301 0 n8 ns301 0 2.57067184171e-05
Gc4_302 0 n8 ns302 0 -1.40082895405e-05
Gc4_303 0 n8 ns303 0 8.3287461971e-05
Gc4_304 0 n8 ns304 0 -0.00030681099672
Gc4_305 0 n8 ns305 0 0.000218415815487
Gc4_306 0 n8 ns306 0 -0.000111322366913
Gc4_307 0 n8 ns307 0 -6.74178321263e-05
Gc4_308 0 n8 ns308 0 9.30386647271e-05
Gc4_309 0 n8 ns309 0 -0.000148106231066
Gc4_310 0 n8 ns310 0 -0.00041413437712
Gc4_311 0 n8 ns311 0 -2.41669154633e-05
Gc4_312 0 n8 ns312 0 0.000592136397415
Gc4_313 0 n8 ns313 0 -0.000450357424941
Gc4_314 0 n8 ns314 0 0.000604687740263
Gc4_315 0 n8 ns315 0 5.48090673032e-05
Gc4_316 0 n8 ns316 0 0.00079587854266
Gc4_317 0 n8 ns317 0 -4.89318681472e-05
Gc4_318 0 n8 ns318 0 4.71458841772e-05
Gc4_319 0 n8 ns319 0 0.000527557007999
Gc4_320 0 n8 ns320 0 -1.84718703836e-05
Gc4_321 0 n8 ns321 0 0.000719672904781
Gc4_322 0 n8 ns322 0 -0.000663440528537
Gc4_323 0 n8 ns323 0 -0.00071047471008
Gc4_324 0 n8 ns324 0 -0.000958691971507
Gc4_325 0 n8 ns325 0 -0.000588365563866
Gc4_326 0 n8 ns326 0 7.4061292149e-05
Gc4_327 0 n8 ns327 0 -0.00097191620275
Gc4_328 0 n8 ns328 0 0.00185802824369
Gc4_329 0 n8 ns329 0 0.0022242031934
Gc4_330 0 n8 ns330 0 0.000745642631063
Gc4_331 0 n8 ns331 0 0.00243377407978
Gc4_332 0 n8 ns332 0 5.45834786387e-05
Gc4_333 0 n8 ns333 0 0.00325281884857
Gc4_334 0 n8 ns334 0 0.000424092745199
Gc4_335 0 n8 ns335 0 -6.74557576297e-05
Gc4_336 0 n8 ns336 0 -2.6533829914e-05
Gc4_337 0 n8 ns337 0 -0.0126635761607
Gc4_338 0 n8 ns338 0 0.000587562607247
Gc4_339 0 n8 ns339 0 0.000327970050067
Gc4_340 0 n8 ns340 0 0.000241245928752
Gc4_341 0 n8 ns341 0 -2.11909104773e-05
Gc4_342 0 n8 ns342 0 -9.97148559081e-06
Gc4_343 0 n8 ns343 0 -0.000273476469671
Gc4_344 0 n8 ns344 0 2.91460202052e-06
Gc4_345 0 n8 ns345 0 -1.42064499814e-06
Gc4_346 0 n8 ns346 0 5.0497214925e-07
Gc4_347 0 n8 ns347 0 9.41336577042e-06
Gc4_348 0 n8 ns348 0 0.000207294295962
Gc4_349 0 n8 ns349 0 0.000237017277886
Gc4_350 0 n8 ns350 0 -9.86084119822e-05
Gc4_351 0 n8 ns351 0 3.11415786365e-06
Gc4_352 0 n8 ns352 0 1.75343462858e-06
Gc4_353 0 n8 ns353 0 -0.000192494158849
Gc4_354 0 n8 ns354 0 5.47645818938e-05
Gc4_355 0 n8 ns355 0 0.000120076598175
Gc4_356 0 n8 ns356 0 0.00028994022435
Gc4_357 0 n8 ns357 0 6.13451445021e-06
Gc4_358 0 n8 ns358 0 -5.29094927658e-06
Gc4_359 0 n8 ns359 0 -0.000171673941687
Gc4_360 0 n8 ns360 0 0.000290001080028
Gc4_361 0 n8 ns361 0 0.000328141610459
Gc4_362 0 n8 ns362 0 0.000103216741285
Gc4_363 0 n8 ns363 0 -2.08703887306e-05
Gc4_364 0 n8 ns364 0 4.4553868163e-05
Gc4_365 0 n8 ns365 0 -4.40987875072e-05
Gc4_366 0 n8 ns366 0 0.000650414073322
Gc4_367 0 n8 ns367 0 -0.000317977401632
Gc4_368 0 n8 ns368 0 0.00020761567266
Gc4_369 0 n8 ns369 0 0.00172389519959
Gc4_370 0 n8 ns370 0 0.000680623946886
Gc4_371 0 n8 ns371 0 -0.000142355202025
Gc4_372 0 n8 ns372 0 0.000363478887129
Gc4_373 0 n8 ns373 0 -0.00071251515981
Gc4_374 0 n8 ns374 0 -4.21514160812e-05
Gc4_375 0 n8 ns375 0 0.000336222462151
Gc4_376 0 n8 ns376 0 0.000236984713848
Gc4_377 0 n8 ns377 0 0.00121533192219
Gc4_378 0 n8 ns378 0 -0.00411994731316
Gc4_379 0 n8 ns379 0 -0.000131468342992
Gc4_380 0 n8 ns380 0 -0.00114414938087
Gc4_381 0 n8 ns381 0 0.000863466853609
Gc4_382 0 n8 ns382 0 -0.00245856274907
Gc4_383 0 n8 ns383 0 -5.26185240399e-05
Gc4_384 0 n8 ns384 0 0.00126710305241
Gc4_385 0 n8 ns385 0 0.00232107796591
Gc4_386 0 n8 ns386 0 0.00205989977433
Gc4_387 0 n8 ns387 0 0.00321714142796
Gc4_388 0 n8 ns388 0 0.00155700597717
Gc4_389 0 n8 ns389 0 0.00445710985616
Gc4_390 0 n8 ns390 0 0.000608694386388
Gc4_391 0 n8 ns391 0 -9.13528499869e-05
Gc4_392 0 n8 ns392 0 -0.000102760511086
Gc4_393 0 n8 ns393 0 -0.00728186158097
Gc4_394 0 n8 ns394 0 -0.000261054130791
Gc4_395 0 n8 ns395 0 -0.000180674102477
Gc4_396 0 n8 ns396 0 -0.000112943319557
Gc4_397 0 n8 ns397 0 -1.7469211333e-05
Gc4_398 0 n8 ns398 0 -3.37318089387e-06
Gc4_399 0 n8 ns399 0 -0.000276117936695
Gc4_400 0 n8 ns400 0 -1.1193723138e-05
Gc4_401 0 n8 ns401 0 4.70813524554e-06
Gc4_402 0 n8 ns402 0 3.53962637651e-06
Gc4_403 0 n8 ns403 0 -2.52655500945e-05
Gc4_404 0 n8 ns404 0 -0.00013740825219
Gc4_405 0 n8 ns405 0 0.000271447491719
Gc4_406 0 n8 ns406 0 -0.000184646970544
Gc4_407 0 n8 ns407 0 -4.60148578928e-06
Gc4_408 0 n8 ns408 0 -1.12467581259e-05
Gc4_409 0 n8 ns409 0 0.00014930657887
Gc4_410 0 n8 ns410 0 -4.92851735604e-05
Gc4_411 0 n8 ns411 0 0.00021102164424
Gc4_412 0 n8 ns412 0 0.000290558350468
Gc4_413 0 n8 ns413 0 -2.73742288894e-05
Gc4_414 0 n8 ns414 0 1.53733793843e-05
Gc4_415 0 n8 ns415 0 -4.42132550362e-06
Gc4_416 0 n8 ns416 0 -0.000231203591868
Gc4_417 0 n8 ns417 0 0.000404388528416
Gc4_418 0 n8 ns418 0 0.000105203209485
Gc4_419 0 n8 ns419 0 5.25300776548e-05
Gc4_420 0 n8 ns420 0 -0.000121145578154
Gc4_421 0 n8 ns421 0 -5.30973755802e-05
Gc4_422 0 n8 ns422 0 -0.000448880188687
Gc4_423 0 n8 ns423 0 -0.000503173807437
Gc4_424 0 n8 ns424 0 8.27211636505e-05
Gc4_425 0 n8 ns425 0 -0.00138548575577
Gc4_426 0 n8 ns426 0 -0.000437845675148
Gc4_427 0 n8 ns427 0 -0.000658863178492
Gc4_428 0 n8 ns428 0 0.000373811611575
Gc4_429 0 n8 ns429 0 0.000339259100866
Gc4_430 0 n8 ns430 0 -2.45652588523e-05
Gc4_431 0 n8 ns431 0 0.000196382669037
Gc4_432 0 n8 ns432 0 0.00032535794698
Gc4_433 0 n8 ns433 0 0.00228124585502
Gc4_434 0 n8 ns434 0 0.00341093346882
Gc4_435 0 n8 ns435 0 0.000636897971166
Gc4_436 0 n8 ns436 0 -0.000933342322679
Gc4_437 0 n8 ns437 0 -1.95607932541e-05
Gc4_438 0 n8 ns438 0 0.00474170405642
Gc4_439 0 n8 ns439 0 -0.00693250320035
Gc4_440 0 n8 ns440 0 0.00196027087989
Gc4_441 0 n8 ns441 0 -0.00179386376687
Gc4_442 0 n8 ns442 0 0.00441396807317
Gc4_443 0 n8 ns443 0 -0.00512712781547
Gc4_444 0 n8 ns444 0 -0.00466717622678
Gc4_445 0 n8 ns445 0 0.0197696618278
Gc4_446 0 n8 ns446 0 -0.000394636055694
Gc4_447 0 n8 ns447 0 9.46215403063e-05
Gc4_448 0 n8 ns448 0 7.0898148958e-05
Gd4_1 0 n8 ni1 0 -0.000949928301852
Gd4_2 0 n8 ni2 0 0.00386358406253
Gd4_3 0 n8 ni3 0 0.00503106662012
Gd4_4 0 n8 ni4 0 -0.00579308485172
Gd4_5 0 n8 ni5 0 0.000203108566201
Gd4_6 0 n8 ni6 0 -0.000467287531536
Gd4_7 0 n8 ni7 0 -0.000111719641059
Gd4_8 0 n8 ni8 0 9.77691500609e-05
Gc5_1 0 n10 ns1 0 -0.00966173118487
Gc5_2 0 n10 ns2 0 0.000617715264017
Gc5_3 0 n10 ns3 0 -0.000189718790319
Gc5_4 0 n10 ns4 0 -0.000279521900908
Gc5_5 0 n10 ns5 0 -2.28942536024e-05
Gc5_6 0 n10 ns6 0 -1.39529295885e-05
Gc5_7 0 n10 ns7 0 -0.000259321336803
Gc5_8 0 n10 ns8 0 -5.45994257144e-05
Gc5_9 0 n10 ns9 0 8.68902320328e-07
Gc5_10 0 n10 ns10 0 -5.04555888124e-07
Gc5_11 0 n10 ns11 0 -8.57745723473e-05
Gc5_12 0 n10 ns12 0 -0.000164894646937
Gc5_13 0 n10 ns13 0 0.000310312038606
Gc5_14 0 n10 ns14 0 -0.000108354182133
Gc5_15 0 n10 ns15 0 -2.02825576136e-06
Gc5_16 0 n10 ns16 0 -2.88029996725e-07
Gc5_17 0 n10 ns17 0 0.000157510986923
Gc5_18 0 n10 ns18 0 -0.000124317391299
Gc5_19 0 n10 ns19 0 0.000114590971595
Gc5_20 0 n10 ns20 0 0.000341523595046
Gc5_21 0 n10 ns21 0 -4.11025691784e-07
Gc5_22 0 n10 ns22 0 5.58709062066e-06
Gc5_23 0 n10 ns23 0 -8.59896475411e-05
Gc5_24 0 n10 ns24 0 -0.000284721383006
Gc5_25 0 n10 ns25 0 0.000325491200056
Gc5_26 0 n10 ns26 0 0.000267354722744
Gc5_27 0 n10 ns27 0 -1.5923595488e-05
Gc5_28 0 n10 ns28 0 -3.9397542984e-05
Gc5_29 0 n10 ns29 0 -0.000305126234043
Gc5_30 0 n10 ns30 0 -0.000371657203451
Gc5_31 0 n10 ns31 0 -0.000524819549201
Gc5_32 0 n10 ns32 0 1.98939370199e-05
Gc5_33 0 n10 ns33 0 -0.000776211341928
Gc5_34 0 n10 ns34 0 0.000590387182642
Gc5_35 0 n10 ns35 0 -0.000659474089078
Gc5_36 0 n10 ns36 0 0.000178372175271
Gc5_37 0 n10 ns37 0 0.000112936944507
Gc5_38 0 n10 ns38 0 -0.000386725924825
Gc5_39 0 n10 ns39 0 1.9585675652e-05
Gc5_40 0 n10 ns40 0 0.000574141165252
Gc5_41 0 n10 ns41 0 0.00335828689104
Gc5_42 0 n10 ns42 0 0.00124133474778
Gc5_43 0 n10 ns43 0 0.00138851197537
Gc5_44 0 n10 ns44 0 -0.000920571592918
Gc5_45 0 n10 ns45 0 0.00132369812636
Gc5_46 0 n10 ns46 0 0.0025813050303
Gc5_47 0 n10 ns47 0 -0.00615029943895
Gc5_48 0 n10 ns48 0 0.000910759465744
Gc5_49 0 n10 ns49 0 -0.00185800796785
Gc5_50 0 n10 ns50 0 0.00569935587707
Gc5_51 0 n10 ns51 0 -0.00438175882636
Gc5_52 0 n10 ns52 0 -0.00320747111898
Gc5_53 0 n10 ns53 0 0.0207123609287
Gc5_54 0 n10 ns54 0 -0.000329575127554
Gc5_55 0 n10 ns55 0 8.31134713519e-05
Gc5_56 0 n10 ns56 0 -3.26484460348e-05
Gc5_57 0 n10 ns57 0 -0.0126554502061
Gc5_58 0 n10 ns58 0 0.000588769965365
Gc5_59 0 n10 ns59 0 0.000327639766297
Gc5_60 0 n10 ns60 0 0.000240251231677
Gc5_61 0 n10 ns61 0 -2.1199543946e-05
Gc5_62 0 n10 ns62 0 -9.9148857968e-06
Gc5_63 0 n10 ns63 0 -0.000273638522034
Gc5_64 0 n10 ns64 0 2.99417358566e-06
Gc5_65 0 n10 ns65 0 -1.42597854921e-06
Gc5_66 0 n10 ns66 0 5.23319458107e-07
Gc5_67 0 n10 ns67 0 9.53028425926e-06
Gc5_68 0 n10 ns68 0 0.000207127838822
Gc5_69 0 n10 ns69 0 0.000237167866135
Gc5_70 0 n10 ns70 0 -9.88891383357e-05
Gc5_71 0 n10 ns71 0 3.12988552484e-06
Gc5_72 0 n10 ns72 0 1.73142152037e-06
Gc5_73 0 n10 ns73 0 -0.000192347736331
Gc5_74 0 n10 ns74 0 5.47383757936e-05
Gc5_75 0 n10 ns75 0 0.000120292853249
Gc5_76 0 n10 ns76 0 0.000290061115799
Gc5_77 0 n10 ns77 0 6.10826120598e-06
Gc5_78 0 n10 ns78 0 -5.30595930246e-06
Gc5_79 0 n10 ns79 0 -0.000171597781531
Gc5_80 0 n10 ns80 0 0.000289904187414
Gc5_81 0 n10 ns81 0 0.000328307769176
Gc5_82 0 n10 ns82 0 0.000102998442536
Gc5_83 0 n10 ns83 0 -2.08724910359e-05
Gc5_84 0 n10 ns84 0 4.45141423022e-05
Gc5_85 0 n10 ns85 0 -4.39904737548e-05
Gc5_86 0 n10 ns86 0 0.000649895609656
Gc5_87 0 n10 ns87 0 -0.00031777944203
Gc5_88 0 n10 ns88 0 0.000208029227763
Gc5_89 0 n10 ns89 0 0.00172349061919
Gc5_90 0 n10 ns90 0 0.00067933575516
Gc5_91 0 n10 ns91 0 -0.000142166872338
Gc5_92 0 n10 ns92 0 0.000363804592729
Gc5_93 0 n10 ns93 0 -0.00071227697736
Gc5_94 0 n10 ns94 0 -4.14702713613e-05
Gc5_95 0 n10 ns95 0 0.000336212856074
Gc5_96 0 n10 ns96 0 0.000236773147297
Gc5_97 0 n10 ns97 0 0.00121258774212
Gc5_98 0 n10 ns98 0 -0.00411907028351
Gc5_99 0 n10 ns99 0 -0.000132192377272
Gc5_100 0 n10 ns100 0 -0.00114372887074
Gc5_101 0 n10 ns101 0 0.000860689728768
Gc5_102 0 n10 ns102 0 -0.00245794908415
Gc5_103 0 n10 ns103 0 -5.32604560186e-05
Gc5_104 0 n10 ns104 0 0.00126582097328
Gc5_105 0 n10 ns105 0 0.00232157442223
Gc5_106 0 n10 ns106 0 0.00205769418782
Gc5_107 0 n10 ns107 0 0.00321778032345
Gc5_108 0 n10 ns108 0 0.00155491550089
Gc5_109 0 n10 ns109 0 0.00445670621953
Gc5_110 0 n10 ns110 0 0.000608524816408
Gc5_111 0 n10 ns111 0 -9.13957743679e-05
Gc5_112 0 n10 ns112 0 -0.000102721789876
Gc5_113 0 n10 ns113 0 0.00410513960189
Gc5_114 0 n10 ns114 0 7.39651644815e-05
Gc5_115 0 n10 ns115 0 -0.000192909791114
Gc5_116 0 n10 ns116 0 -0.000281569400946
Gc5_117 0 n10 ns117 0 1.15492662173e-05
Gc5_118 0 n10 ns118 0 2.80589282623e-05
Gc5_119 0 n10 ns119 0 4.65957079044e-05
Gc5_120 0 n10 ns120 0 3.30218275956e-05
Gc5_121 0 n10 ns121 0 -1.39762250048e-07
Gc5_122 0 n10 ns122 0 -2.32625740368e-07
Gc5_123 0 n10 ns123 0 8.1783859207e-06
Gc5_124 0 n10 ns124 0 -0.000267802150606
Gc5_125 0 n10 ns125 0 -9.08756794559e-05
Gc5_126 0 n10 ns126 0 -0.000114995918407
Gc5_127 0 n10 ns127 0 9.53562468433e-07
Gc5_128 0 n10 ns128 0 1.65877456632e-07
Gc5_129 0 n10 ns129 0 0.000297755066068
Gc5_130 0 n10 ns130 0 -3.40126644089e-05
Gc5_131 0 n10 ns131 0 0.000128552461829
Gc5_132 0 n10 ns132 0 -0.000124974693734
Gc5_133 0 n10 ns133 0 1.84335663807e-07
Gc5_134 0 n10 ns134 0 -3.70048389766e-06
Gc5_135 0 n10 ns135 0 0.000179930290333
Gc5_136 0 n10 ns136 0 -0.000433280092544
Gc5_137 0 n10 ns137 0 2.60080330077e-05
Gc5_138 0 n10 ns138 0 -0.000219770549068
Gc5_139 0 n10 ns139 0 -1.92007513107e-06
Gc5_140 0 n10 ns140 0 1.02553997197e-05
Gc5_141 0 n10 ns141 0 -1.09620153522e-06
Gc5_142 0 n10 ns142 0 -0.000836228597647
Gc5_143 0 n10 ns143 0 0.000157977798758
Gc5_144 0 n10 ns144 0 0.000415009385618
Gc5_145 0 n10 ns145 0 -0.00161092477203
Gc5_146 0 n10 ns146 0 -0.000276257464599
Gc5_147 0 n10 ns147 0 0.000142059356231
Gc5_148 0 n10 ns148 0 0.00054716302741
Gc5_149 0 n10 ns149 0 0.00052589071387
Gc5_150 0 n10 ns150 0 0.00018908719047
Gc5_151 0 n10 ns151 0 0.000372483621195
Gc5_152 0 n10 ns152 0 -0.000195297210923
Gc5_153 0 n10 ns153 0 -0.000740119444705
Gc5_154 0 n10 ns154 0 0.00224474371318
Gc5_155 0 n10 ns155 0 -0.000798348629308
Gc5_156 0 n10 ns156 0 -0.000247462604111
Gc5_157 0 n10 ns157 0 -0.00181778598031
Gc5_158 0 n10 ns158 0 0.00180957927609
Gc5_159 0 n10 ns159 0 -0.00120937884253
Gc5_160 0 n10 ns160 0 0.00117387779498
Gc5_161 0 n10 ns161 0 0.00145364252892
Gc5_162 0 n10 ns162 0 -0.000441616352751
Gc5_163 0 n10 ns163 0 0.00152048735557
Gc5_164 0 n10 ns164 0 -0.000929481847367
Gc5_165 0 n10 ns165 0 0.0017654657725
Gc5_166 0 n10 ns166 0 0.000106014243689
Gc5_167 0 n10 ns167 0 -4.38085740323e-05
Gc5_168 0 n10 ns168 0 2.94830890058e-05
Gc5_169 0 n10 ns169 0 -0.000708846116416
Gc5_170 0 n10 ns170 0 -0.000224480904634
Gc5_171 0 n10 ns171 0 0.000253696571054
Gc5_172 0 n10 ns172 0 0.00013183045723
Gc5_173 0 n10 ns173 0 -2.08036948988e-07
Gc5_174 0 n10 ns174 0 1.61934932536e-05
Gc5_175 0 n10 ns175 0 -3.36133874159e-05
Gc5_176 0 n10 ns176 0 7.33010676962e-05
Gc5_177 0 n10 ns177 0 5.5452095861e-08
Gc5_178 0 n10 ns178 0 1.50835653348e-07
Gc5_179 0 n10 ns179 0 6.47127822743e-05
Gc5_180 0 n10 ns180 0 0.000124941676473
Gc5_181 0 n10 ns181 0 -5.22043197693e-05
Gc5_182 0 n10 ns182 0 -9.00406080742e-05
Gc5_183 0 n10 ns183 0 1.68541230161e-08
Gc5_184 0 n10 ns184 0 -1.33181386065e-06
Gc5_185 0 n10 ns185 0 -9.2028087844e-05
Gc5_186 0 n10 ns186 0 9.74246813493e-05
Gc5_187 0 n10 ns187 0 0.000122229745495
Gc5_188 0 n10 ns188 0 -4.03014391709e-05
Gc5_189 0 n10 ns189 0 -6.59933457689e-06
Gc5_190 0 n10 ns190 0 3.31651642513e-06
Gc5_191 0 n10 ns191 0 1.31787737769e-05
Gc5_192 0 n10 ns192 0 0.000194952292586
Gc5_193 0 n10 ns193 0 9.62415134388e-05
Gc5_194 0 n10 ns194 0 -0.000208947483302
Gc5_195 0 n10 ns195 0 2.73410866932e-05
Gc5_196 0 n10 ns196 0 -3.77876329657e-05
Gc5_197 0 n10 ns197 0 0.000241459106645
Gc5_198 0 n10 ns198 0 0.00015793393701
Gc5_199 0 n10 ns199 0 2.79455237713e-05
Gc5_200 0 n10 ns200 0 0.000131271502126
Gc5_201 0 n10 ns201 0 0.000111928923664
Gc5_202 0 n10 ns202 0 -0.000695062313473
Gc5_203 0 n10 ns203 0 0.000119480994894
Gc5_204 0 n10 ns204 0 0.000189399903169
Gc5_205 0 n10 ns205 0 1.95653506518e-05
Gc5_206 0 n10 ns206 0 0.00036625653239
Gc5_207 0 n10 ns207 0 0.000188933444885
Gc5_208 0 n10 ns208 0 -0.000143746649701
Gc5_209 0 n10 ns209 0 -0.0011035924057
Gc5_210 0 n10 ns210 0 2.02209100133e-05
Gc5_211 0 n10 ns211 0 -0.000646740173943
Gc5_212 0 n10 ns212 0 -0.000330557786299
Gc5_213 0 n10 ns213 0 -0.00128330440882
Gc5_214 0 n10 ns214 0 0.000171296352683
Gc5_215 0 n10 ns215 0 -0.00053608222333
Gc5_216 0 n10 ns216 0 0.000866505355592
Gc5_217 0 n10 ns217 0 0.00142574144803
Gc5_218 0 n10 ns218 0 6.10038557404e-06
Gc5_219 0 n10 ns219 0 0.00110640652754
Gc5_220 0 n10 ns220 0 -0.000246878922
Gc5_221 0 n10 ns221 0 0.00104585752855
Gc5_222 0 n10 ns222 0 0.000374733309088
Gc5_223 0 n10 ns223 0 -3.40616425777e-05
Gc5_224 0 n10 ns224 0 -1.7476478383e-05
Gc5_225 0 n10 ns225 0 0.00373953716142
Gc5_226 0 n10 ns226 0 0.0104330876249
Gc5_227 0 n10 ns227 0 -0.00225046406573
Gc5_228 0 n10 ns228 0 -0.000725222901665
Gc5_229 0 n10 ns229 0 3.25389796732e-05
Gc5_230 0 n10 ns230 0 -4.25635621301e-06
Gc5_231 0 n10 ns231 0 0.000115515365363
Gc5_232 0 n10 ns232 0 3.99809351591e-05
Gc5_233 0 n10 ns233 0 5.39270185124e-07
Gc5_234 0 n10 ns234 0 -1.66622788832e-06
Gc5_235 0 n10 ns235 0 -6.6779084368e-05
Gc5_236 0 n10 ns236 0 -5.06061913437e-05
Gc5_237 0 n10 ns237 0 0.000201359462477
Gc5_238 0 n10 ns238 0 5.4727142193e-06
Gc5_239 0 n10 ns239 0 1.93377929724e-06
Gc5_240 0 n10 ns240 0 -1.82030214386e-06
Gc5_241 0 n10 ns241 0 -8.52140794431e-06
Gc5_242 0 n10 ns242 0 6.60557312833e-05
Gc5_243 0 n10 ns243 0 7.85756668849e-06
Gc5_244 0 n10 ns244 0 -0.000163906284372
Gc5_245 0 n10 ns245 0 4.45961626188e-06
Gc5_246 0 n10 ns246 0 3.7271411431e-06
Gc5_247 0 n10 ns247 0 -0.000102470627417
Gc5_248 0 n10 ns248 0 -1.55415209452e-05
Gc5_249 0 n10 ns249 0 0.000100099074938
Gc5_250 0 n10 ns250 0 8.15950879571e-05
Gc5_251 0 n10 ns251 0 2.45708280342e-05
Gc5_252 0 n10 ns252 0 -4.22371724236e-06
Gc5_253 0 n10 ns253 0 3.16086411828e-05
Gc5_254 0 n10 ns254 0 -0.000155947275121
Gc5_255 0 n10 ns255 0 0.000169978839717
Gc5_256 0 n10 ns256 0 1.70004595324e-05
Gc5_257 0 n10 ns257 0 0.000205850928456
Gc5_258 0 n10 ns258 0 -5.76634647474e-05
Gc5_259 0 n10 ns259 0 -0.000356077691821
Gc5_260 0 n10 ns260 0 4.63890071769e-05
Gc5_261 0 n10 ns261 0 0.00022008983367
Gc5_262 0 n10 ns262 0 3.22895165006e-05
Gc5_263 0 n10 ns263 0 -0.000104796513513
Gc5_264 0 n10 ns264 0 -0.000339996079533
Gc5_265 0 n10 ns265 0 -0.00061706589335
Gc5_266 0 n10 ns266 0 -0.000331799337421
Gc5_267 0 n10 ns267 0 0.000893652795652
Gc5_268 0 n10 ns268 0 -0.000935505207159
Gc5_269 0 n10 ns269 0 0.000397811011368
Gc5_270 0 n10 ns270 0 0.000530630168743
Gc5_271 0 n10 ns271 0 0.0031626001531
Gc5_272 0 n10 ns272 0 0.000392941862708
Gc5_273 0 n10 ns273 0 -0.000466862711079
Gc5_274 0 n10 ns274 0 0.00379793084227
Gc5_275 0 n10 ns275 0 -0.00103687835115
Gc5_276 0 n10 ns276 0 -0.00157097078005
Gc5_277 0 n10 ns277 0 -0.0108288732574
Gc5_278 0 n10 ns278 0 -0.000579251273077
Gc5_279 0 n10 ns279 0 7.61928276784e-05
Gc5_280 0 n10 ns280 0 0.000129184653553
Gc5_281 0 n10 ns281 0 -0.00150285623456
Gc5_282 0 n10 ns282 0 -0.000701783195441
Gc5_283 0 n10 ns283 0 0.000556065738819
Gc5_284 0 n10 ns284 0 0.000735985748933
Gc5_285 0 n10 ns285 0 2.35689713181e-05
Gc5_286 0 n10 ns286 0 6.87438069893e-06
Gc5_287 0 n10 ns287 0 0.000195704108555
Gc5_288 0 n10 ns288 0 3.3763491583e-05
Gc5_289 0 n10 ns289 0 -8.87306063851e-07
Gc5_290 0 n10 ns290 0 1.19085225036e-06
Gc5_291 0 n10 ns291 0 6.84516349173e-06
Gc5_292 0 n10 ns292 0 0.000152720119104
Gc5_293 0 n10 ns293 0 0.000257393028297
Gc5_294 0 n10 ns294 0 -0.000132461065155
Gc5_295 0 n10 ns295 0 -1.8729013795e-06
Gc5_296 0 n10 ns296 0 -1.39252131416e-07
Gc5_297 0 n10 ns297 0 0.000163078121054
Gc5_298 0 n10 ns298 0 -2.59107191603e-05
Gc5_299 0 n10 ns299 0 -0.000173268471304
Gc5_300 0 n10 ns300 0 -0.000296120279968
Gc5_301 0 n10 ns301 0 2.3108078078e-06
Gc5_302 0 n10 ns302 0 -6.55499345195e-06
Gc5_303 0 n10 ns303 0 -5.97346179852e-05
Gc5_304 0 n10 ns304 0 0.000193727865602
Gc5_305 0 n10 ns305 0 0.000387427499852
Gc5_306 0 n10 ns306 0 0.000206228733282
Gc5_307 0 n10 ns307 0 -1.44591335851e-05
Gc5_308 0 n10 ns308 0 -4.76705369981e-05
Gc5_309 0 n10 ns309 0 4.07416974731e-05
Gc5_310 0 n10 ns310 0 -0.000267750036671
Gc5_311 0 n10 ns311 0 0.000541633163976
Gc5_312 0 n10 ns312 0 -0.000133278647017
Gc5_313 0 n10 ns313 0 0.000738144511838
Gc5_314 0 n10 ns314 0 -5.53346319422e-05
Gc5_315 0 n10 ns315 0 -0.00060824352433
Gc5_316 0 n10 ns316 0 0.00017841316581
Gc5_317 0 n10 ns317 0 0.00059330337504
Gc5_318 0 n10 ns318 0 -0.000194168995694
Gc5_319 0 n10 ns319 0 -0.000211478843811
Gc5_320 0 n10 ns320 0 -0.000249537337668
Gc5_321 0 n10 ns321 0 -0.00114733679239
Gc5_322 0 n10 ns322 0 -0.00101003855774
Gc5_323 0 n10 ns323 0 0.000464868895437
Gc5_324 0 n10 ns324 0 -0.00112064905618
Gc5_325 0 n10 ns325 0 0.00102977773907
Gc5_326 0 n10 ns326 0 0.000650729515193
Gc5_327 0 n10 ns327 0 0.0027261370427
Gc5_328 0 n10 ns328 0 -3.00970457073e-05
Gc5_329 0 n10 ns329 0 0.000627178729365
Gc5_330 0 n10 ns330 0 0.00241167119569
Gc5_331 0 n10 ns331 0 -0.000143064408475
Gc5_332 0 n10 ns332 0 -0.00226490260076
Gc5_333 0 n10 ns333 0 -0.0067902337452
Gc5_334 0 n10 ns334 0 -0.000652193811253
Gc5_335 0 n10 ns335 0 4.34328245723e-05
Gc5_336 0 n10 ns336 0 0.000115026288744
Gc5_337 0 n10 ns337 0 0.0317283470933
Gc5_338 0 n10 ns338 0 -0.00566448264868
Gc5_339 0 n10 ns339 0 -0.000893246044298
Gc5_340 0 n10 ns340 0 0.00147129073008
Gc5_341 0 n10 ns341 0 -1.83404873415e-05
Gc5_342 0 n10 ns342 0 -3.06875713692e-05
Gc5_343 0 n10 ns343 0 -1.53120048157e-05
Gc5_344 0 n10 ns344 0 -2.67976729419e-05
Gc5_345 0 n10 ns345 0 2.45824865101e-07
Gc5_346 0 n10 ns346 0 2.19400686064e-07
Gc5_347 0 n10 ns347 0 -2.82635556027e-05
Gc5_348 0 n10 ns348 0 -0.000295173455148
Gc5_349 0 n10 ns349 0 -5.98247907886e-05
Gc5_350 0 n10 ns350 0 -0.000153964052992
Gc5_351 0 n10 ns351 0 -6.28729996181e-07
Gc5_352 0 n10 ns352 0 5.10185189794e-08
Gc5_353 0 n10 ns353 0 -0.000325519152696
Gc5_354 0 n10 ns354 0 4.22868690163e-05
Gc5_355 0 n10 ns355 0 -0.000115136897867
Gc5_356 0 n10 ns356 0 8.44976051612e-05
Gc5_357 0 n10 ns357 0 2.61315031426e-06
Gc5_358 0 n10 ns358 0 -2.36408134814e-06
Gc5_359 0 n10 ns359 0 0.000152178701007
Gc5_360 0 n10 ns360 0 -0.000386914293834
Gc5_361 0 n10 ns361 0 -4.0556098378e-05
Gc5_362 0 n10 ns362 0 -0.000212094032177
Gc5_363 0 n10 ns363 0 1.45524184149e-05
Gc5_364 0 n10 ns364 0 -4.41226141782e-05
Gc5_365 0 n10 ns365 0 -0.000314471808119
Gc5_366 0 n10 ns366 0 0.000685589250093
Gc5_367 0 n10 ns367 0 -0.000142226453185
Gc5_368 0 n10 ns368 0 -0.000165020881631
Gc5_369 0 n10 ns369 0 -0.00114018726059
Gc5_370 0 n10 ns370 0 6.94538282311e-06
Gc5_371 0 n10 ns371 0 0.000374143887164
Gc5_372 0 n10 ns372 0 0.000435283427584
Gc5_373 0 n10 ns373 0 -0.00074108772698
Gc5_374 0 n10 ns374 0 -1.6434380898e-05
Gc5_375 0 n10 ns375 0 -0.000249332611927
Gc5_376 0 n10 ns376 0 5.33263553438e-05
Gc5_377 0 n10 ns377 0 -5.59883870567e-06
Gc5_378 0 n10 ns378 0 0.00264664128961
Gc5_379 0 n10 ns379 0 -0.00104041205127
Gc5_380 0 n10 ns380 0 -0.000249350358385
Gc5_381 0 n10 ns381 0 0.000170432792143
Gc5_382 0 n10 ns382 0 -0.000973806605226
Gc5_383 0 n10 ns383 0 -1.12889990198e-05
Gc5_384 0 n10 ns384 0 -0.00206129440872
Gc5_385 0 n10 ns385 0 0.0010433723841
Gc5_386 0 n10 ns386 0 0.000181110086772
Gc5_387 0 n10 ns387 0 -0.00030562688415
Gc5_388 0 n10 ns388 0 -4.97365599704e-05
Gc5_389 0 n10 ns389 0 -0.000936912668901
Gc5_390 0 n10 ns390 0 -0.000165083615534
Gc5_391 0 n10 ns391 0 5.1045386714e-05
Gc5_392 0 n10 ns392 0 2.63069186387e-05
Gc5_393 0 n10 ns393 0 0.0227365254859
Gc5_394 0 n10 ns394 0 0.00024737892784
Gc5_395 0 n10 ns395 0 0.000313788009964
Gc5_396 0 n10 ns396 0 0.000215631187573
Gc5_397 0 n10 ns397 0 -1.14431610426e-05
Gc5_398 0 n10 ns398 0 -1.45995602269e-05
Gc5_399 0 n10 ns399 0 0.000115106618321
Gc5_400 0 n10 ns400 0 -8.77359054758e-05
Gc5_401 0 n10 ns401 0 -4.32658833746e-07
Gc5_402 0 n10 ns402 0 1.29273002986e-08
Gc5_403 0 n10 ns403 0 4.19293633716e-05
Gc5_404 0 n10 ns404 0 8.14266055514e-05
Gc5_405 0 n10 ns405 0 2.24710528268e-06
Gc5_406 0 n10 ns406 0 -0.000149844189271
Gc5_407 0 n10 ns407 0 -2.7282569846e-07
Gc5_408 0 n10 ns408 0 4.93919710429e-07
Gc5_409 0 n10 ns409 0 9.66567994527e-05
Gc5_410 0 n10 ns410 0 -6.61819423385e-05
Gc5_411 0 n10 ns411 0 -0.000161356456186
Gc5_412 0 n10 ns412 0 3.54523590466e-06
Gc5_413 0 n10 ns413 0 -4.54366300924e-06
Gc5_414 0 n10 ns414 0 1.68703032882e-06
Gc5_415 0 n10 ns415 0 1.85557505587e-05
Gc5_416 0 n10 ns416 0 0.000176601824223
Gc5_417 0 n10 ns417 0 0.000123014889825
Gc5_418 0 n10 ns418 0 -0.000129393777286
Gc5_419 0 n10 ns419 0 -2.99105086544e-05
Gc5_420 0 n10 ns420 0 2.13580530057e-05
Gc5_421 0 n10 ns421 0 -0.000201547309772
Gc5_422 0 n10 ns422 0 -0.000198619833058
Gc5_423 0 n10 ns423 0 2.45219095407e-05
Gc5_424 0 n10 ns424 0 -0.000297053808884
Gc5_425 0 n10 ns425 0 -2.75325393025e-06
Gc5_426 0 n10 ns426 0 -0.00047406613718
Gc5_427 0 n10 ns427 0 -4.06588662316e-05
Gc5_428 0 n10 ns428 0 0.000425780972
Gc5_429 0 n10 ns429 0 1.17410463306e-05
Gc5_430 0 n10 ns430 0 -0.000322934252083
Gc5_431 0 n10 ns431 0 -0.000233358570933
Gc5_432 0 n10 ns432 0 9.15931328387e-05
Gc5_433 0 n10 ns433 0 -0.000925181618168
Gc5_434 0 n10 ns434 0 0.00029788362242
Gc5_435 0 n10 ns435 0 -0.000507791807537
Gc5_436 0 n10 ns436 0 -0.000609889885196
Gc5_437 0 n10 ns437 0 0.00104990363383
Gc5_438 0 n10 ns438 0 -0.000407409139617
Gc5_439 0 n10 ns439 0 0.00108942207085
Gc5_440 0 n10 ns440 0 -0.00151641533951
Gc5_441 0 n10 ns441 0 0.00123084276992
Gc5_442 0 n10 ns442 0 0.000288841712548
Gc5_443 0 n10 ns443 0 -0.000147651942704
Gc5_444 0 n10 ns444 0 -0.000657357614496
Gc5_445 0 n10 ns445 0 -0.000757785539821
Gc5_446 0 n10 ns446 0 -0.000455334084986
Gc5_447 0 n10 ns447 0 1.88771379458e-05
Gc5_448 0 n10 ns448 0 5.13818923513e-05
Gd5_1 0 n10 ni1 0 -0.000469964191059
Gd5_2 0 n10 ni2 0 -0.000114546867779
Gd5_3 0 n10 ni3 0 -0.000178703045241
Gd5_4 0 n10 ni4 0 0.000203109476833
Gd5_5 0 n10 ni5 0 -0.00409478211339
Gd5_6 0 n10 ni6 0 0.00502994506362
Gd5_7 0 n10 ni7 0 0.00314084446859
Gd5_8 0 n10 ni8 0 -0.000942875049348
Gc6_1 0 n12 ns1 0 -0.0126486701595
Gc6_2 0 n12 ns2 0 0.00058592425693
Gc6_3 0 n12 ns3 0 0.000327970348009
Gc6_4 0 n12 ns4 0 0.000240798153268
Gc6_5 0 n12 ns5 0 -2.12051243082e-05
Gc6_6 0 n12 ns6 0 -9.93016756076e-06
Gc6_7 0 n12 ns7 0 -0.000273571451096
Gc6_8 0 n12 ns8 0 3.13950490992e-06
Gc6_9 0 n12 ns9 0 -1.42174054602e-06
Gc6_10 0 n12 ns10 0 5.23048361583e-07
Gc6_11 0 n12 ns11 0 9.52674218418e-06
Gc6_12 0 n12 ns12 0 0.000207241614472
Gc6_13 0 n12 ns13 0 0.000236998940091
Gc6_14 0 n12 ns14 0 -9.88608343428e-05
Gc6_15 0 n12 ns15 0 3.12550410826e-06
Gc6_16 0 n12 ns16 0 1.73435932112e-06
Gc6_17 0 n12 ns17 0 -0.000192407693121
Gc6_18 0 n12 ns18 0 5.47390088525e-05
Gc6_19 0 n12 ns19 0 0.000120412246123
Gc6_20 0 n12 ns20 0 0.000289835738596
Gc6_21 0 n12 ns21 0 6.12391235926e-06
Gc6_22 0 n12 ns22 0 -5.30001742121e-06
Gc6_23 0 n12 ns23 0 -0.000171653178249
Gc6_24 0 n12 ns24 0 0.000290000856016
Gc6_25 0 n12 ns25 0 0.000328163714525
Gc6_26 0 n12 ns26 0 0.000102838165658
Gc6_27 0 n12 ns27 0 -2.09263168651e-05
Gc6_28 0 n12 ns28 0 4.45712631338e-05
Gc6_29 0 n12 ns29 0 -4.44081606595e-05
Gc6_30 0 n12 ns30 0 0.000649983120622
Gc6_31 0 n12 ns31 0 -0.000317639438208
Gc6_32 0 n12 ns32 0 0.000208206394017
Gc6_33 0 n12 ns33 0 0.00172282213216
Gc6_34 0 n12 ns34 0 0.000679350699091
Gc6_35 0 n12 ns35 0 -0.000142081236059
Gc6_36 0 n12 ns36 0 0.000363996046113
Gc6_37 0 n12 ns37 0 -0.000712563803758
Gc6_38 0 n12 ns38 0 -4.17448845772e-05
Gc6_39 0 n12 ns39 0 0.000336359566098
Gc6_40 0 n12 ns40 0 0.000236316825737
Gc6_41 0 n12 ns41 0 0.0012122105021
Gc6_42 0 n12 ns42 0 -0.00411695684065
Gc6_43 0 n12 ns43 0 -0.000132255982964
Gc6_44 0 n12 ns44 0 -0.0011438185518
Gc6_45 0 n12 ns45 0 0.000860041369421
Gc6_46 0 n12 ns46 0 -0.00245879425833
Gc6_47 0 n12 ns47 0 -5.32063059794e-05
Gc6_48 0 n12 ns48 0 0.00126482555628
Gc6_49 0 n12 ns49 0 0.0023214744804
Gc6_50 0 n12 ns50 0 0.00205861251366
Gc6_51 0 n12 ns51 0 0.00321798913498
Gc6_52 0 n12 ns52 0 0.00155578224983
Gc6_53 0 n12 ns53 0 0.00445566222925
Gc6_54 0 n12 ns54 0 0.000608809036688
Gc6_55 0 n12 ns55 0 -9.13844864236e-05
Gc6_56 0 n12 ns56 0 -0.00010285358431
Gc6_57 0 n12 ns57 0 -0.00729018175256
Gc6_58 0 n12 ns58 0 -0.000258427985427
Gc6_59 0 n12 ns59 0 -0.000180799086596
Gc6_60 0 n12 ns60 0 -0.000113503804897
Gc6_61 0 n12 ns61 0 -1.74097302587e-05
Gc6_62 0 n12 ns62 0 -3.32152918811e-06
Gc6_63 0 n12 ns63 0 -0.000275694431839
Gc6_64 0 n12 ns64 0 -1.10141410364e-05
Gc6_65 0 n12 ns65 0 4.71336841484e-06
Gc6_66 0 n12 ns66 0 3.51765367699e-06
Gc6_67 0 n12 ns67 0 -2.53759943266e-05
Gc6_68 0 n12 ns68 0 -0.000137896180755
Gc6_69 0 n12 ns69 0 0.000270808207223
Gc6_70 0 n12 ns70 0 -0.000184682327559
Gc6_71 0 n12 ns71 0 -4.61974897794e-06
Gc6_72 0 n12 ns72 0 -1.12265372741e-05
Gc6_73 0 n12 ns73 0 0.00014981984997
Gc6_74 0 n12 ns74 0 -4.94717992915e-05
Gc6_75 0 n12 ns75 0 0.000211014496529
Gc6_76 0 n12 ns76 0 0.000289872535689
Gc6_77 0 n12 ns77 0 -2.73481457464e-05
Gc6_78 0 n12 ns78 0 1.53901206934e-05
Gc6_79 0 n12 ns79 0 -4.31773789863e-06
Gc6_80 0 n12 ns80 0 -0.00023197674165
Gc6_81 0 n12 ns81 0 0.000403836228828
Gc6_82 0 n12 ns82 0 0.000104618140805
Gc6_83 0 n12 ns83 0 5.25058531718e-05
Gc6_84 0 n12 ns84 0 -0.000121125616736
Gc6_85 0 n12 ns85 0 -5.35634680642e-05
Gc6_86 0 n12 ns86 0 -0.000450250738493
Gc6_87 0 n12 ns87 0 -0.000502070782065
Gc6_88 0 n12 ns88 0 8.26435791026e-05
Gc6_89 0 n12 ns89 0 -0.00138709228503
Gc6_90 0 n12 ns90 0 -0.000436265887166
Gc6_91 0 n12 ns91 0 -0.000657878583924
Gc6_92 0 n12 ns92 0 0.000373086058497
Gc6_93 0 n12 ns93 0 0.000340041072881
Gc6_94 0 n12 ns94 0 -2.57294833895e-05
Gc6_95 0 n12 ns95 0 0.000195901859503
Gc6_96 0 n12 ns96 0 0.000324940645557
Gc6_97 0 n12 ns97 0 0.00228189095733
Gc6_98 0 n12 ns98 0 0.00341304490605
Gc6_99 0 n12 ns99 0 0.00063761739422
Gc6_100 0 n12 ns100 0 -0.000932054361634
Gc6_101 0 n12 ns101 0 -1.75287958432e-05
Gc6_102 0 n12 ns102 0 0.00474193977577
Gc6_103 0 n12 ns103 0 -0.00693096280821
Gc6_104 0 n12 ns104 0 0.00195858305269
Gc6_105 0 n12 ns105 0 -0.00179584659148
Gc6_106 0 n12 ns106 0 0.00441460060752
Gc6_107 0 n12 ns107 0 -0.00512717208205
Gc6_108 0 n12 ns108 0 -0.00466611347812
Gc6_109 0 n12 ns109 0 0.0197683324374
Gc6_110 0 n12 ns110 0 -0.000394757835409
Gc6_111 0 n12 ns111 0 9.4616489505e-05
Gc6_112 0 n12 ns112 0 7.09150175236e-05
Gc6_113 0 n12 ns113 0 -0.000744364087226
Gc6_114 0 n12 ns114 0 -0.000221958475148
Gc6_115 0 n12 ns115 0 0.000254139951579
Gc6_116 0 n12 ns116 0 0.000131764793499
Gc6_117 0 n12 ns117 0 -2.34094071023e-07
Gc6_118 0 n12 ns118 0 1.61557404681e-05
Gc6_119 0 n12 ns119 0 -3.38830576061e-05
Gc6_120 0 n12 ns120 0 7.31724148212e-05
Gc6_121 0 n12 ns121 0 6.05587036079e-08
Gc6_122 0 n12 ns122 0 1.64266715619e-07
Gc6_123 0 n12 ns123 0 6.48774184994e-05
Gc6_124 0 n12 ns124 0 0.000125412901507
Gc6_125 0 n12 ns125 0 -5.18515470895e-05
Gc6_126 0 n12 ns126 0 -8.99369433592e-05
Gc6_127 0 n12 ns127 0 2.10029427615e-08
Gc6_128 0 n12 ns128 0 -1.35466864887e-06
Gc6_129 0 n12 ns129 0 -9.23899058356e-05
Gc6_130 0 n12 ns130 0 9.76942479133e-05
Gc6_131 0 n12 ns131 0 0.000122171916672
Gc6_132 0 n12 ns132 0 -3.97922828585e-05
Gc6_133 0 n12 ns133 0 -6.65164496608e-06
Gc6_134 0 n12 ns134 0 3.32491315128e-06
Gc6_135 0 n12 ns135 0 1.31124594213e-05
Gc6_136 0 n12 ns136 0 0.000195719644485
Gc6_137 0 n12 ns137 0 9.64946786706e-05
Gc6_138 0 n12 ns138 0 -0.000208541181006
Gc6_139 0 n12 ns139 0 2.74963161006e-05
Gc6_140 0 n12 ns140 0 -3.79022749377e-05
Gc6_141 0 n12 ns141 0 0.000242233107283
Gc6_142 0 n12 ns142 0 0.000158984209904
Gc6_143 0 n12 ns143 0 2.71573120787e-05
Gc6_144 0 n12 ns144 0 0.000130631776175
Gc6_145 0 n12 ns145 0 0.000115264988978
Gc6_146 0 n12 ns146 0 -0.000695986262254
Gc6_147 0 n12 ns147 0 0.000118548016978
Gc6_148 0 n12 ns148 0 0.000188397101741
Gc6_149 0 n12 ns149 0 1.89366248432e-05
Gc6_150 0 n12 ns150 0 0.000366010162957
Gc6_151 0 n12 ns151 0 0.000188898662035
Gc6_152 0 n12 ns152 0 -0.000143075864846
Gc6_153 0 n12 ns153 0 -0.00110509678819
Gc6_154 0 n12 ns154 0 1.68291205369e-05
Gc6_155 0 n12 ns155 0 -0.000646019948825
Gc6_156 0 n12 ns156 0 -0.000330912547501
Gc6_157 0 n12 ns157 0 -0.00128294094264
Gc6_158 0 n12 ns158 0 0.000170985018671
Gc6_159 0 n12 ns159 0 -0.000536784276152
Gc6_160 0 n12 ns160 0 0.000867122756758
Gc6_161 0 n12 ns161 0 0.00142302535823
Gc6_162 0 n12 ns162 0 4.27163287951e-06
Gc6_163 0 n12 ns163 0 0.00110440386823
Gc6_164 0 n12 ns164 0 -0.000246125241555
Gc6_165 0 n12 ns165 0 0.00104594246771
Gc6_166 0 n12 ns166 0 0.000374586797553
Gc6_167 0 n12 ns167 0 -3.40889521337e-05
Gc6_168 0 n12 ns168 0 -1.75496313092e-05
Gc6_169 0 n12 ns169 0 -0.00295366322829
Gc6_170 0 n12 ns170 0 0.000696564275762
Gc6_171 0 n12 ns171 0 -7.59294380685e-05
Gc6_172 0 n12 ns172 0 -0.000153144621264
Gc6_173 0 n12 ns173 0 -2.51954382964e-06
Gc6_174 0 n12 ns174 0 1.67256636257e-05
Gc6_175 0 n12 ns175 0 -0.000108937603532
Gc6_176 0 n12 ns176 0 3.39059846431e-05
Gc6_177 0 n12 ns177 0 -4.42016466766e-06
Gc6_178 0 n12 ns178 0 -4.11863144484e-06
Gc6_179 0 n12 ns179 0 1.91017870263e-06
Gc6_180 0 n12 ns180 0 -0.000183525635833
Gc6_181 0 n12 ns181 0 6.0660070919e-05
Gc6_182 0 n12 ns182 0 -0.000176032145241
Gc6_183 0 n12 ns183 0 4.35320470071e-06
Gc6_184 0 n12 ns184 0 1.09132152433e-05
Gc6_185 0 n12 ns185 0 0.000198104387541
Gc6_186 0 n12 ns186 0 -2.39914484232e-05
Gc6_187 0 n12 ns187 0 0.000192576629562
Gc6_188 0 n12 ns188 0 4.62861110102e-05
Gc6_189 0 n12 ns189 0 2.57067405104e-05
Gc6_190 0 n12 ns190 0 -1.40084225718e-05
Gc6_191 0 n12 ns191 0 8.32930528744e-05
Gc6_192 0 n12 ns192 0 -0.000306814822441
Gc6_193 0 n12 ns193 0 0.000218418623579
Gc6_194 0 n12 ns194 0 -0.000111321221357
Gc6_195 0 n12 ns195 0 -6.74178885151e-05
Gc6_196 0 n12 ns196 0 9.3039699529e-05
Gc6_197 0 n12 ns197 0 -0.000148104056865
Gc6_198 0 n12 ns198 0 -0.000414136507413
Gc6_199 0 n12 ns199 0 -2.41670619445e-05
Gc6_200 0 n12 ns200 0 0.000592139039454
Gc6_201 0 n12 ns201 0 -0.0004503725091
Gc6_202 0 n12 ns202 0 0.000604682465123
Gc6_203 0 n12 ns203 0 5.48113285655e-05
Gc6_204 0 n12 ns204 0 0.000795888249517
Gc6_205 0 n12 ns205 0 -4.89322017239e-05
Gc6_206 0 n12 ns206 0 4.71442409334e-05
Gc6_207 0 n12 ns207 0 0.000527561066959
Gc6_208 0 n12 ns208 0 -1.84733554039e-05
Gc6_209 0 n12 ns209 0 0.000719661455711
Gc6_210 0 n12 ns210 0 -0.000663394771539
Gc6_211 0 n12 ns211 0 -0.000710499588721
Gc6_212 0 n12 ns212 0 -0.000958696198967
Gc6_213 0 n12 ns213 0 -0.000588386801703
Gc6_214 0 n12 ns214 0 7.40848245256e-05
Gc6_215 0 n12 ns215 0 -0.000971941695681
Gc6_216 0 n12 ns216 0 0.00185803494127
Gc6_217 0 n12 ns217 0 0.00222422020224
Gc6_218 0 n12 ns218 0 0.00074561585252
Gc6_219 0 n12 ns219 0 0.00243378429129
Gc6_220 0 n12 ns220 0 5.4559218397e-05
Gc6_221 0 n12 ns221 0 0.00325283596836
Gc6_222 0 n12 ns222 0 0.000424091769606
Gc6_223 0 n12 ns223 0 -6.74553899832e-05
Gc6_224 0 n12 ns224 0 -2.65309273779e-05
Gc6_225 0 n12 ns225 0 -0.00150294646391
Gc6_226 0 n12 ns226 0 -0.00070177055124
Gc6_227 0 n12 ns227 0 0.00055606690199
Gc6_228 0 n12 ns228 0 0.000735984373996
Gc6_229 0 n12 ns229 0 2.35689257224e-05
Gc6_230 0 n12 ns230 0 6.87434176619e-06
Gc6_231 0 n12 ns231 0 0.000195704386662
Gc6_232 0 n12 ns232 0 3.37636925967e-05
Gc6_233 0 n12 ns233 0 -8.87300795839e-07
Gc6_234 0 n12 ns234 0 1.19086516056e-06
Gc6_235 0 n12 ns235 0 6.84492305428e-06
Gc6_236 0 n12 ns236 0 0.000152720243621
Gc6_237 0 n12 ns237 0 0.000257392579829
Gc6_238 0 n12 ns238 0 -0.000132461122141
Gc6_239 0 n12 ns239 0 -1.87289725162e-06
Gc6_240 0 n12 ns240 0 -1.39277707152e-07
Gc6_241 0 n12 ns241 0 0.000163077843853
Gc6_242 0 n12 ns242 0 -2.59109896517e-05
Gc6_243 0 n12 ns243 0 -0.000173269214846
Gc6_244 0 n12 ns244 0 -0.000296119884497
Gc6_245 0 n12 ns245 0 2.31081563248e-06
Gc6_246 0 n12 ns246 0 -6.55496872411e-06
Gc6_247 0 n12 ns247 0 -5.97357599136e-05
Gc6_248 0 n12 ns248 0 0.000193728551705
Gc6_249 0 n12 ns249 0 0.000387426475768
Gc6_250 0 n12 ns250 0 0.000206228047659
Gc6_251 0 n12 ns251 0 -1.44591816608e-05
Gc6_252 0 n12 ns252 0 -4.76707085377e-05
Gc6_253 0 n12 ns253 0 4.07417289044e-05
Gc6_254 0 n12 ns254 0 -0.000267750546822
Gc6_255 0 n12 ns255 0 0.000541632818593
Gc6_256 0 n12 ns256 0 -0.000133278855485
Gc6_257 0 n12 ns257 0 0.000738150229409
Gc6_258 0 n12 ns258 0 -5.53334731281e-05
Gc6_259 0 n12 ns259 0 -0.000608243483405
Gc6_260 0 n12 ns260 0 0.000178407324476
Gc6_261 0 n12 ns261 0 0.000593302374576
Gc6_262 0 n12 ns262 0 -0.000194170179028
Gc6_263 0 n12 ns263 0 -0.00021147942328
Gc6_264 0 n12 ns264 0 -0.000249536262505
Gc6_265 0 n12 ns265 0 -0.00114734179781
Gc6_266 0 n12 ns266 0 -0.00101005436042
Gc6_267 0 n12 ns267 0 0.000464879885527
Gc6_268 0 n12 ns268 0 -0.00112064688222
Gc6_269 0 n12 ns269 0 0.00102977879847
Gc6_270 0 n12 ns270 0 0.000650710708279
Gc6_271 0 n12 ns271 0 0.00272614466236
Gc6_272 0 n12 ns272 0 -3.01085615371e-05
Gc6_273 0 n12 ns273 0 0.000627175028039
Gc6_274 0 n12 ns274 0 0.00241168380955
Gc6_275 0 n12 ns275 0 -0.000143061022576
Gc6_276 0 n12 ns276 0 -0.00226489027545
Gc6_277 0 n12 ns277 0 -0.00679023638501
Gc6_278 0 n12 ns278 0 -0.000652191661093
Gc6_279 0 n12 ns279 0 4.34328345039e-05
Gc6_280 0 n12 ns280 0 0.000115025271811
Gc6_281 0 n12 ns281 0 0.0152231986625
Gc6_282 0 n12 ns282 0 0.01023625606
Gc6_283 0 n12 ns283 0 -0.00245791219965
Gc6_284 0 n12 ns284 0 -0.000975460788254
Gc6_285 0 n12 ns285 0 2.2326420267e-05
Gc6_286 0 n12 ns286 0 -1.32319315002e-05
Gc6_287 0 n12 ns287 0 0.00017986503932
Gc6_288 0 n12 ns288 0 -9.61096238669e-06
Gc6_289 0 n12 ns289 0 3.76827601573e-06
Gc6_290 0 n12 ns290 0 1.37127015345e-06
Gc6_291 0 n12 ns291 0 -1.98829165007e-05
Gc6_292 0 n12 ns292 0 -5.02137137805e-05
Gc6_293 0 n12 ns293 0 0.000177368249433
Gc6_294 0 n12 ns294 0 -7.22272248026e-05
Gc6_295 0 n12 ns295 0 3.70532970686e-06
Gc6_296 0 n12 ns296 0 5.07600554703e-06
Gc6_297 0 n12 ns297 0 1.85775465217e-05
Gc6_298 0 n12 ns298 0 2.61177569448e-06
Gc6_299 0 n12 ns299 0 -6.81117861904e-05
Gc6_300 0 n12 ns300 0 -0.000113440102995
Gc6_301 0 n12 ns301 0 -1.2764432522e-05
Gc6_302 0 n12 ns302 0 1.04944687899e-05
Gc6_303 0 n12 ns303 0 -4.59832690585e-05
Gc6_304 0 n12 ns304 0 8.93657449894e-05
Gc6_305 0 n12 ns305 0 0.000111370327803
Gc6_306 0 n12 ns306 0 -6.18707915278e-05
Gc6_307 0 n12 ns307 0 -2.31828982565e-05
Gc6_308 0 n12 ns308 0 5.13004337989e-05
Gc6_309 0 n12 ns309 0 -0.000206130788694
Gc6_310 0 n12 ns310 0 -0.00031499126033
Gc6_311 0 n12 ns311 0 9.98579576705e-05
Gc6_312 0 n12 ns312 0 -0.000231046914436
Gc6_313 0 n12 ns313 0 5.33106530795e-06
Gc6_314 0 n12 ns314 0 -0.000575049387917
Gc6_315 0 n12 ns315 0 -0.000285770130687
Gc6_316 0 n12 ns316 0 0.000395681106947
Gc6_317 0 n12 ns317 0 2.0496203204e-05
Gc6_318 0 n12 ns318 0 -0.000222687726265
Gc6_319 0 n12 ns319 0 -0.000238084029166
Gc6_320 0 n12 ns320 0 -0.000203275440143
Gc6_321 0 n12 ns321 0 -0.00109160061164
Gc6_322 0 n12 ns322 0 0.000257413279092
Gc6_323 0 n12 ns323 0 0.000343109285634
Gc6_324 0 n12 ns324 0 -0.000987881331346
Gc6_325 0 n12 ns325 0 0.000841173044435
Gc6_326 0 n12 ns326 0 -1.16232218362e-05
Gc6_327 0 n12 ns327 0 0.0030520964152
Gc6_328 0 n12 ns328 0 -0.00048536722243
Gc6_329 0 n12 ns329 0 -0.000125843934403
Gc6_330 0 n12 ns330 0 0.00327057352881
Gc6_331 0 n12 ns331 0 -0.00134640940249
Gc6_332 0 n12 ns332 0 -0.00156992129156
Gc6_333 0 n12 ns333 0 -0.0100653132962
Gc6_334 0 n12 ns334 0 -0.000505319601219
Gc6_335 0 n12 ns335 0 6.2905434553e-05
Gc6_336 0 n12 ns336 0 6.68476395111e-05
Gc6_337 0 n12 ns337 0 0.022701760751
Gc6_338 0 n12 ns338 0 0.000252259727838
Gc6_339 0 n12 ns339 0 0.00031506116041
Gc6_340 0 n12 ns340 0 0.00021526314778
Gc6_341 0 n12 ns341 0 -1.14173028547e-05
Gc6_342 0 n12 ns342 0 -1.46024568619e-05
Gc6_343 0 n12 ns343 0 0.000115162602811
Gc6_344 0 n12 ns344 0 -8.75359768045e-05
Gc6_345 0 n12 ns345 0 -4.36825681761e-07
Gc6_346 0 n12 ns346 0 1.86691858299e-08
Gc6_347 0 n12 ns347 0 4.20777667901e-05
Gc6_348 0 n12 ns348 0 8.17893743178e-05
Gc6_349 0 n12 ns349 0 2.60293820366e-06
Gc6_350 0 n12 ns350 0 -0.000149747271963
Gc6_351 0 n12 ns351 0 -2.77444072104e-07
Gc6_352 0 n12 ns352 0 5.07422949469e-07
Gc6_353 0 n12 ns353 0 9.70227093451e-05
Gc6_354 0 n12 ns354 0 -6.62284395082e-05
Gc6_355 0 n12 ns355 0 -0.000161495804646
Gc6_356 0 n12 ns356 0 3.2689754981e-06
Gc6_357 0 n12 ns357 0 -4.54534241282e-06
Gc6_358 0 n12 ns358 0 1.66975108158e-06
Gc6_359 0 n12 ns359 0 1.8412373826e-05
Gc6_360 0 n12 ns360 0 0.000176997173097
Gc6_361 0 n12 ns361 0 0.000123469067189
Gc6_362 0 n12 ns362 0 -0.000129100622172
Gc6_363 0 n12 ns363 0 -2.98857209294e-05
Gc6_364 0 n12 ns364 0 2.13766369738e-05
Gc6_365 0 n12 ns365 0 -0.000200983342025
Gc6_366 0 n12 ns366 0 -0.000199739472576
Gc6_367 0 n12 ns367 0 2.49698922069e-05
Gc6_368 0 n12 ns368 0 -0.000296694577896
Gc6_369 0 n12 ns369 0 -1.33362479621e-06
Gc6_370 0 n12 ns370 0 -0.000473752264702
Gc6_371 0 n12 ns371 0 -4.13740777348e-05
Gc6_372 0 n12 ns372 0 0.000425261607289
Gc6_373 0 n12 ns373 0 1.23835647866e-05
Gc6_374 0 n12 ns374 0 -0.000323271363238
Gc6_375 0 n12 ns375 0 -0.000233252372566
Gc6_376 0 n12 ns376 0 9.12105083538e-05
Gc6_377 0 n12 ns377 0 -0.000925990230101
Gc6_378 0 n12 ns378 0 0.000296161675305
Gc6_379 0 n12 ns379 0 -0.00050686080233
Gc6_380 0 n12 ns380 0 -0.000610324269974
Gc6_381 0 n12 ns381 0 0.00105044604219
Gc6_382 0 n12 ns382 0 -0.000407069124459
Gc6_383 0 n12 ns383 0 0.00109104826258
Gc6_384 0 n12 ns384 0 -0.00151586387256
Gc6_385 0 n12 ns385 0 0.00122914943243
Gc6_386 0 n12 ns386 0 0.000288922041169
Gc6_387 0 n12 ns387 0 -0.000148871183118
Gc6_388 0 n12 ns388 0 -0.00065519090521
Gc6_389 0 n12 ns389 0 -0.000758773357874
Gc6_390 0 n12 ns390 0 -0.000454952512082
Gc6_391 0 n12 ns391 0 1.88437615906e-05
Gc6_392 0 n12 ns392 0 5.12801227128e-05
Gc6_393 0 n12 ns393 0 0.0161651182913
Gc6_394 0 n12 ns394 0 -0.00290362821089
Gc6_395 0 n12 ns395 0 -0.000319131733572
Gc6_396 0 n12 ns396 0 0.00100250051139
Gc6_397 0 n12 ns397 0 3.99984818196e-08
Gc6_398 0 n12 ns398 0 -9.72265561124e-06
Gc6_399 0 n12 ns399 0 0.000114967178648
Gc6_400 0 n12 ns400 0 -9.76712331819e-06
Gc6_401 0 n12 ns401 0 -3.18432138283e-06
Gc6_402 0 n12 ns402 0 -2.35011329715e-06
Gc6_403 0 n12 ns403 0 -1.35669610806e-05
Gc6_404 0 n12 ns404 0 -0.000156161515378
Gc6_405 0 n12 ns405 0 8.2187230939e-05
Gc6_406 0 n12 ns406 0 -0.000161727862212
Gc6_407 0 n12 ns407 0 -2.49893525604e-06
Gc6_408 0 n12 ns408 0 -7.01697403991e-06
Gc6_409 0 n12 ns409 0 -0.000163593363377
Gc6_410 0 n12 ns410 0 1.90199117575e-05
Gc6_411 0 n12 ns411 0 -0.000152498742581
Gc6_412 0 n12 ns412 0 -8.08000425025e-05
Gc6_413 0 n12 ns413 0 2.00095753365e-05
Gc6_414 0 n12 ns414 0 -9.54632110667e-06
Gc6_415 0 n12 ns415 0 8.79361376114e-05
Gc6_416 0 n12 ns416 0 -0.000191934352724
Gc6_417 0 n12 ns417 0 0.000159558152201
Gc6_418 0 n12 ns418 0 -1.6919488742e-05
Gc6_419 0 n12 ns419 0 4.23992372711e-05
Gc6_420 0 n12 ns420 0 -0.000100934185141
Gc6_421 0 n12 ns421 0 -0.000150818914821
Gc6_422 0 n12 ns422 0 0.000446834645969
Gc6_423 0 n12 ns423 0 0.000158376585548
Gc6_424 0 n12 ns424 0 -9.9972148388e-05
Gc6_425 0 n12 ns425 0 -0.000317692272103
Gc6_426 0 n12 ns426 0 0.000121203012724
Gc6_427 0 n12 ns427 0 -1.4154094763e-05
Gc6_428 0 n12 ns428 0 0.000313527596244
Gc6_429 0 n12 ns429 0 -6.38341804687e-05
Gc6_430 0 n12 ns430 0 -9.10017499958e-05
Gc6_431 0 n12 ns431 0 -0.0003027646432
Gc6_432 0 n12 ns432 0 -3.04058859679e-05
Gc6_433 0 n12 ns433 0 -0.000487519140929
Gc6_434 0 n12 ns434 0 0.000714335589184
Gc6_435 0 n12 ns435 0 -0.000439540784628
Gc6_436 0 n12 ns436 0 -0.000774672821594
Gc6_437 0 n12 ns437 0 0.00087204119982
Gc6_438 0 n12 ns438 0 -6.3368462549e-05
Gc6_439 0 n12 ns439 0 0.00150324842178
Gc6_440 0 n12 ns440 0 -0.00125391224777
Gc6_441 0 n12 ns441 0 0.00114268992556
Gc6_442 0 n12 ns442 0 0.00115250167682
Gc6_443 0 n12 ns443 0 -0.000215621343264
Gc6_444 0 n12 ns444 0 -0.00129621561235
Gc6_445 0 n12 ns445 0 -0.00352822410492
Gc6_446 0 n12 ns446 0 -0.000541467372229
Gc6_447 0 n12 ns447 0 4.33082324805e-05
Gc6_448 0 n12 ns448 0 7.31842942451e-05
Gd6_1 0 n12 ni1 0 -0.000111451372926
Gd6_2 0 n12 ni2 0 9.70822724551e-05
Gd6_3 0 n12 ni3 0 0.000201925531561
Gd6_4 0 n12 ni4 0 -0.000467282381193
Gd6_5 0 n12 ni5 0 0.00502994142612
Gd6_6 0 n12 ni6 0 -0.00579595099873
Gd6_7 0 n12 ni7 0 -0.000942618188439
Gd6_8 0 n12 ni8 0 0.0038641771003
Gc7_1 0 n14 ns1 0 0.00409729877302
Gc7_2 0 n14 ns2 0 7.53350207968e-05
Gc7_3 0 n14 ns3 0 -0.000192526721015
Gc7_4 0 n14 ns4 0 -0.000281886813134
Gc7_5 0 n14 ns5 0 1.15191381175e-05
Gc7_6 0 n14 ns6 0 2.80361241674e-05
Gc7_7 0 n14 ns7 0 4.6541776328e-05
Gc7_8 0 n14 ns8 0 3.30192817185e-05
Gc7_9 0 n14 ns9 0 -1.4047813143e-07
Gc7_10 0 n14 ns10 0 -2.33155233171e-07
Gc7_11 0 n14 ns11 0 8.36585251869e-06
Gc7_12 0 n14 ns12 0 -0.000267058416161
Gc7_13 0 n14 ns13 0 -9.07103304197e-05
Gc7_14 0 n14 ns14 0 -0.00011472320116
Gc7_15 0 n14 ns15 0 9.53176753731e-07
Gc7_16 0 n14 ns16 0 1.66913717674e-07
Gc7_17 0 n14 ns17 0 0.00029706504609
Gc7_18 0 n14 ns18 0 -3.37958637397e-05
Gc7_19 0 n14 ns19 0 0.000128456510867
Gc7_20 0 n14 ns20 0 -0.000124799650118
Gc7_21 0 n14 ns21 0 1.80543195857e-07
Gc7_22 0 n14 ns22 0 -3.69317217867e-06
Gc7_23 0 n14 ns23 0 0.000179773654959
Gc7_24 0 n14 ns24 0 -0.000432063201539
Gc7_25 0 n14 ns25 0 2.5976286332e-05
Gc7_26 0 n14 ns26 0 -0.000219573433001
Gc7_27 0 n14 ns27 0 -1.92916180755e-06
Gc7_28 0 n14 ns28 0 1.0220954658e-05
Gc7_29 0 n14 ns29 0 -1.04610737513e-06
Gc7_30 0 n14 ns30 0 -0.00083492980557
Gc7_31 0 n14 ns31 0 0.000157715642983
Gc7_32 0 n14 ns32 0 0.000414545850657
Gc7_33 0 n14 ns33 0 -0.00160917929242
Gc7_34 0 n14 ns34 0 -0.00027610671218
Gc7_35 0 n14 ns35 0 0.000142009928039
Gc7_36 0 n14 ns36 0 0.000546320780642
Gc7_37 0 n14 ns37 0 0.000525647918974
Gc7_38 0 n14 ns38 0 0.000188863488387
Gc7_39 0 n14 ns39 0 0.000372141013406
Gc7_40 0 n14 ns40 0 -0.0001949854207
Gc7_41 0 n14 ns41 0 -0.00074016905017
Gc7_42 0 n14 ns42 0 0.00224253014739
Gc7_43 0 n14 ns43 0 -0.000798005398459
Gc7_44 0 n14 ns44 0 -0.000246909051312
Gc7_45 0 n14 ns45 0 -0.0018166089551
Gc7_46 0 n14 ns46 0 0.00180810673359
Gc7_47 0 n14 ns47 0 -0.00120877287295
Gc7_48 0 n14 ns48 0 0.00117320895151
Gc7_49 0 n14 ns49 0 0.00145331033361
Gc7_50 0 n14 ns50 0 -0.000441791127069
Gc7_51 0 n14 ns51 0 0.00152084020735
Gc7_52 0 n14 ns52 0 -0.000928293725829
Gc7_53 0 n14 ns53 0 0.00176739926573
Gc7_54 0 n14 ns54 0 0.000105948396154
Gc7_55 0 n14 ns55 0 -4.37789020684e-05
Gc7_56 0 n14 ns56 0 2.94043022357e-05
Gc7_57 0 n14 ns57 0 -0.000734084775673
Gc7_58 0 n14 ns58 0 -0.000221627834149
Gc7_59 0 n14 ns59 0 0.000253496886367
Gc7_60 0 n14 ns60 0 0.000131180482792
Gc7_61 0 n14 ns61 0 -2.20824952352e-07
Gc7_62 0 n14 ns62 0 1.61373781732e-05
Gc7_63 0 n14 ns63 0 -3.38400534828e-05
Gc7_64 0 n14 ns64 0 7.30229681963e-05
Gc7_65 0 n14 ns65 0 5.17511749454e-08
Gc7_66 0 n14 ns66 0 1.5725961548e-07
Gc7_67 0 n14 ns67 0 6.4650164125e-05
Gc7_68 0 n14 ns68 0 0.000124841291013
Gc7_69 0 n14 ns69 0 -5.17915376801e-05
Gc7_70 0 n14 ns70 0 -8.98811367407e-05
Gc7_71 0 n14 ns71 0 2.52186912434e-08
Gc7_72 0 n14 ns72 0 -1.33791462198e-06
Gc7_73 0 n14 ns73 0 -9.18623304514e-05
Gc7_74 0 n14 ns74 0 9.73567448841e-05
Gc7_75 0 n14 ns75 0 0.000122058170976
Gc7_76 0 n14 ns76 0 -3.9769954774e-05
Gc7_77 0 n14 ns77 0 -6.60400417682e-06
Gc7_78 0 n14 ns78 0 3.304172397e-06
Gc7_79 0 n14 ns79 0 1.31278870371e-05
Gc7_80 0 n14 ns80 0 0.000194725804006
Gc7_81 0 n14 ns81 0 9.64031632289e-05
Gc7_82 0 n14 ns82 0 -0.000208345521633
Gc7_83 0 n14 ns83 0 2.73715660916e-05
Gc7_84 0 n14 ns84 0 -3.77294312407e-05
Gc7_85 0 n14 ns85 0 0.000241752176852
Gc7_86 0 n14 ns86 0 0.000157883291545
Gc7_87 0 n14 ns87 0 2.75563786291e-05
Gc7_88 0 n14 ns88 0 0.000130809741906
Gc7_89 0 n14 ns89 0 0.000114251516371
Gc7_90 0 n14 ns90 0 -0.000695419845633
Gc7_91 0 n14 ns91 0 0.000119014538529
Gc7_92 0 n14 ns92 0 0.000188871141219
Gc7_93 0 n14 ns93 0 1.90603962347e-05
Gc7_94 0 n14 ns94 0 0.00036636367151
Gc7_95 0 n14 ns95 0 0.00018870312711
Gc7_96 0 n14 ns96 0 -0.000143157972957
Gc7_97 0 n14 ns97 0 -0.00110329828315
Gc7_98 0 n14 ns98 0 1.65855720304e-05
Gc7_99 0 n14 ns99 0 -0.000646285245197
Gc7_100 0 n14 ns100 0 -0.000330620402875
Gc7_101 0 n14 ns101 0 -0.00128197382538
Gc7_102 0 n14 ns102 0 0.000170971424536
Gc7_103 0 n14 ns103 0 -0.000536345057895
Gc7_104 0 n14 ns104 0 0.000867317529899
Gc7_105 0 n14 ns105 0 0.00142265704064
Gc7_106 0 n14 ns106 0 4.43866079477e-06
Gc7_107 0 n14 ns107 0 0.00110384936945
Gc7_108 0 n14 ns108 0 -0.000245417395624
Gc7_109 0 n14 ns109 0 0.00104634444745
Gc7_110 0 n14 ns110 0 0.000374512385767
Gc7_111 0 n14 ns111 0 -3.41198070151e-05
Gc7_112 0 n14 ns112 0 -1.76169773239e-05
Gc7_113 0 n14 ns113 0 -0.00964333201632
Gc7_114 0 n14 ns114 0 0.000616989496973
Gc7_115 0 n14 ns115 0 -0.000189964392306
Gc7_116 0 n14 ns116 0 -0.000279533904327
Gc7_117 0 n14 ns117 0 -2.28295054824e-05
Gc7_118 0 n14 ns118 0 -1.39628739495e-05
Gc7_119 0 n14 ns119 0 -0.000258674349355
Gc7_120 0 n14 ns120 0 -5.47102764986e-05
Gc7_121 0 n14 ns121 0 8.72759738021e-07
Gc7_122 0 n14 ns122 0 -5.04046507266e-07
Gc7_123 0 n14 ns123 0 -8.58859269333e-05
Gc7_124 0 n14 ns124 0 -0.000165106604082
Gc7_125 0 n14 ns125 0 0.000309708695007
Gc7_126 0 n14 ns126 0 -0.000107831648789
Gc7_127 0 n14 ns127 0 -2.03113457818e-06
Gc7_128 0 n14 ns128 0 -2.94452446583e-07
Gc7_129 0 n14 ns129 0 0.000157747186676
Gc7_130 0 n14 ns130 0 -0.000124461816191
Gc7_131 0 n14 ns131 0 0.000114040404854
Gc7_132 0 n14 ns132 0 0.000340895966555
Gc7_133 0 n14 ns133 0 -4.24926733864e-07
Gc7_134 0 n14 ns134 0 5.58895687072e-06
Gc7_135 0 n14 ns135 0 -8.58529658047e-05
Gc7_136 0 n14 ns136 0 -0.000285082423901
Gc7_137 0 n14 ns137 0 0.000324508565211
Gc7_138 0 n14 ns138 0 0.000267276089156
Gc7_139 0 n14 ns139 0 -1.58872091079e-05
Gc7_140 0 n14 ns140 0 -3.94181836912e-05
Gc7_141 0 n14 ns141 0 -0.000305108344907
Gc7_142 0 n14 ns142 0 -0.000372558636748
Gc7_143 0 n14 ns143 0 -0.000523914373349
Gc7_144 0 n14 ns144 0 1.91831673303e-05
Gc7_145 0 n14 ns145 0 -0.000778194051347
Gc7_146 0 n14 ns146 0 0.000589706563861
Gc7_147 0 n14 ns147 0 -0.000658673892282
Gc7_148 0 n14 ns148 0 0.000177079878632
Gc7_149 0 n14 ns149 0 0.000114066053242
Gc7_150 0 n14 ns150 0 -0.000386822539966
Gc7_151 0 n14 ns151 0 1.84950187272e-05
Gc7_152 0 n14 ns152 0 0.000573521055956
Gc7_153 0 n14 ns153 0 0.0033548073038
Gc7_154 0 n14 ns154 0 0.00124640203707
Gc7_155 0 n14 ns155 0 0.00138918150266
Gc7_156 0 n14 ns156 0 -0.000917501794193
Gc7_157 0 n14 ns157 0 0.00132080463256
Gc7_158 0 n14 ns158 0 0.00258180223106
Gc7_159 0 n14 ns159 0 -0.00614874740679
Gc7_160 0 n14 ns160 0 0.000904393115748
Gc7_161 0 n14 ns161 0 -0.00186074466976
Gc7_162 0 n14 ns162 0 0.00569710367468
Gc7_163 0 n14 ns163 0 -0.00437945756311
Gc7_164 0 n14 ns164 0 -0.00320896886433
Gc7_165 0 n14 ns165 0 0.020707365795
Gc7_166 0 n14 ns166 0 -0.00032972112301
Gc7_167 0 n14 ns167 0 8.29591794433e-05
Gc7_168 0 n14 ns168 0 -3.25720369945e-05
Gc7_169 0 n14 ns169 0 -0.0126635783834
Gc7_170 0 n14 ns170 0 0.000587561737418
Gc7_171 0 n14 ns171 0 0.000327971432596
Gc7_172 0 n14 ns172 0 0.000241244344429
Gc7_173 0 n14 ns173 0 -2.11909084987e-05
Gc7_174 0 n14 ns174 0 -9.97152489888e-06
Gc7_175 0 n14 ns175 0 -0.000273476569886
Gc7_176 0 n14 ns176 0 2.91483760064e-06
Gc7_177 0 n14 ns177 0 -1.42064845044e-06
Gc7_178 0 n14 ns178 0 5.04970388263e-07
Gc7_179 0 n14 ns179 0 9.41354773316e-06
Gc7_180 0 n14 ns180 0 0.000207294366025
Gc7_181 0 n14 ns181 0 0.000237017332928
Gc7_182 0 n14 ns182 0 -9.86082565869e-05
Gc7_183 0 n14 ns183 0 3.11416110348e-06
Gc7_184 0 n14 ns184 0 1.75343764025e-06
Gc7_185 0 n14 ns185 0 -0.000192494011794
Gc7_186 0 n14 ns186 0 5.47645895897e-05
Gc7_187 0 n14 ns187 0 0.000120076740517
Gc7_188 0 n14 ns188 0 0.000289940269136
Gc7_189 0 n14 ns189 0 6.13451720533e-06
Gc7_190 0 n14 ns190 0 -5.29095652959e-06
Gc7_191 0 n14 ns191 0 -0.000171673820884
Gc7_192 0 n14 ns192 0 0.00029000100962
Gc7_193 0 n14 ns193 0 0.000328141709996
Gc7_194 0 n14 ns194 0 0.000103216647027
Gc7_195 0 n14 ns195 0 -2.08703399755e-05
Gc7_196 0 n14 ns196 0 4.45539207176e-05
Gc7_197 0 n14 ns197 0 -4.40986569518e-05
Gc7_198 0 n14 ns198 0 0.000650413689495
Gc7_199 0 n14 ns199 0 -0.000317977441382
Gc7_200 0 n14 ns200 0 0.000207615621083
Gc7_201 0 n14 ns201 0 0.00172389583789
Gc7_202 0 n14 ns202 0 0.000680623669568
Gc7_203 0 n14 ns203 0 -0.000142355280653
Gc7_204 0 n14 ns204 0 0.000363478757628
Gc7_205 0 n14 ns205 0 -0.000712514493856
Gc7_206 0 n14 ns206 0 -4.2151146355e-05
Gc7_207 0 n14 ns207 0 0.000336222504853
Gc7_208 0 n14 ns208 0 0.000236985839373
Gc7_209 0 n14 ns209 0 0.00121533104919
Gc7_210 0 n14 ns210 0 -0.00411995084001
Gc7_211 0 n14 ns211 0 -0.000131468826306
Gc7_212 0 n14 ns212 0 -0.00114414918418
Gc7_213 0 n14 ns213 0 0.000863469221301
Gc7_214 0 n14 ns214 0 -0.00245856364246
Gc7_215 0 n14 ns215 0 -5.26172362301e-05
Gc7_216 0 n14 ns216 0 0.00126710335098
Gc7_217 0 n14 ns217 0 0.00232107738286
Gc7_218 0 n14 ns218 0 0.00205989854887
Gc7_219 0 n14 ns219 0 0.00321713859693
Gc7_220 0 n14 ns220 0 0.00155700531156
Gc7_221 0 n14 ns221 0 0.00445710765253
Gc7_222 0 n14 ns222 0 0.000608694639353
Gc7_223 0 n14 ns223 0 -9.13527911948e-05
Gc7_224 0 n14 ns224 0 -0.000102760549479
Gc7_225 0 n14 ns225 0 0.0317282955165
Gc7_226 0 n14 ns226 0 -0.00566447737038
Gc7_227 0 n14 ns227 0 -0.000893245166735
Gc7_228 0 n14 ns228 0 0.00147129047193
Gc7_229 0 n14 ns229 0 -1.83405045113e-05
Gc7_230 0 n14 ns230 0 -3.06876115535e-05
Gc7_231 0 n14 ns231 0 -1.53120845832e-05
Gc7_232 0 n14 ns232 0 -2.67975407382e-05
Gc7_233 0 n14 ns233 0 2.4582708374e-07
Gc7_234 0 n14 ns234 0 2.1940258525e-07
Gc7_235 0 n14 ns235 0 -2.82635739116e-05
Gc7_236 0 n14 ns236 0 -0.000295173336632
Gc7_237 0 n14 ns237 0 -5.98249102712e-05
Gc7_238 0 n14 ns238 0 -0.000153964024671
Gc7_239 0 n14 ns239 0 -6.28729060486e-07
Gc7_240 0 n14 ns240 0 5.10132328773e-08
Gc7_241 0 n14 ns241 0 -0.000325519066991
Gc7_242 0 n14 ns242 0 4.22868549077e-05
Gc7_243 0 n14 ns243 0 -0.000115136942213
Gc7_244 0 n14 ns244 0 8.44977232639e-05
Gc7_245 0 n14 ns245 0 2.61315041841e-06
Gc7_246 0 n14 ns246 0 -2.36407238506e-06
Gc7_247 0 n14 ns247 0 0.0001521783737
Gc7_248 0 n14 ns248 0 -0.000386913834488
Gc7_249 0 n14 ns249 0 -4.0556292882e-05
Gc7_250 0 n14 ns250 0 -0.000212094121986
Gc7_251 0 n14 ns251 0 1.45524354547e-05
Gc7_252 0 n14 ns252 0 -4.41226591691e-05
Gc7_253 0 n14 ns253 0 -0.000314471948757
Gc7_254 0 n14 ns254 0 0.000685588869307
Gc7_255 0 n14 ns255 0 -0.00014222650386
Gc7_256 0 n14 ns256 0 -0.000165020852341
Gc7_257 0 n14 ns257 0 -0.00114018572299
Gc7_258 0 n14 ns258 0 6.94459988251e-06
Gc7_259 0 n14 ns259 0 0.000374142971522
Gc7_260 0 n14 ns260 0 0.000435282726558
Gc7_261 0 n14 ns261 0 -0.000741087865494
Gc7_262 0 n14 ns262 0 -1.64344638723e-05
Gc7_263 0 n14 ns263 0 -0.000249332638546
Gc7_264 0 n14 ns264 0 5.33267521564e-05
Gc7_265 0 n14 ns265 0 -5.60008971605e-06
Gc7_266 0 n14 ns266 0 0.00264663770534
Gc7_267 0 n14 ns267 0 -0.00104040976647
Gc7_268 0 n14 ns268 0 -0.000249350926534
Gc7_269 0 n14 ns269 0 0.000170433481224
Gc7_270 0 n14 ns270 0 -0.000973809271011
Gc7_271 0 n14 ns271 0 -1.12877034703e-05
Gc7_272 0 n14 ns272 0 -0.00206129516234
Gc7_273 0 n14 ns273 0 0.001043370777
Gc7_274 0 n14 ns274 0 0.000181112218451
Gc7_275 0 n14 ns275 0 -0.00030562840906
Gc7_276 0 n14 ns276 0 -4.97347320635e-05
Gc7_277 0 n14 ns277 0 -0.000936915534456
Gc7_278 0 n14 ns278 0 -0.000165082976165
Gc7_279 0 n14 ns279 0 5.10454717881e-05
Gc7_280 0 n14 ns280 0 2.63067862338e-05
Gc7_281 0 n14 ns281 0 0.0227016405955
Gc7_282 0 n14 ns282 0 0.000252278817551
Gc7_283 0 n14 ns283 0 0.000315065288138
Gc7_284 0 n14 ns284 0 0.000215265346213
Gc7_285 0 n14 ns285 0 -1.14173793651e-05
Gc7_286 0 n14 ns286 0 -1.46025690153e-05
Gc7_287 0 n14 ns287 0 0.000115162705045
Gc7_288 0 n14 ns288 0 -8.75355871731e-05
Gc7_289 0 n14 ns289 0 -4.36813401824e-07
Gc7_290 0 n14 ns290 0 1.86853984513e-08
Gc7_291 0 n14 ns291 0 4.20773281141e-05
Gc7_292 0 n14 ns292 0 8.17894883384e-05
Gc7_293 0 n14 ns293 0 2.6022281167e-06
Gc7_294 0 n14 ns294 0 -0.000149747658187
Gc7_295 0 n14 ns295 0 -2.77458679425e-07
Gc7_296 0 n14 ns296 0 5.07372672677e-07
Gc7_297 0 n14 ns297 0 9.70224931543e-05
Gc7_298 0 n14 ns298 0 -6.62286342478e-05
Gc7_299 0 n14 ns299 0 -0.000161496240599
Gc7_300 0 n14 ns300 0 3.2691315335e-06
Gc7_301 0 n14 ns301 0 -4.54535916963e-06
Gc7_302 0 n14 ns302 0 1.66980389679e-06
Gc7_303 0 n14 ns303 0 1.84105688632e-05
Gc7_304 0 n14 ns304 0 0.000176998764168
Gc7_305 0 n14 ns305 0 0.000123468697542
Gc7_306 0 n14 ns306 0 -0.000129100806713
Gc7_307 0 n14 ns307 0 -2.98855476991e-05
Gc7_308 0 n14 ns308 0 2.1376220731e-05
Gc7_309 0 n14 ns309 0 -0.00020098455727
Gc7_310 0 n14 ns310 0 -0.000199739023974
Gc7_311 0 n14 ns311 0 2.49698928833e-05
Gc7_312 0 n14 ns312 0 -0.000296695266485
Gc7_313 0 n14 ns313 0 -1.32784801689e-06
Gc7_314 0 n14 ns314 0 -0.000473754568345
Gc7_315 0 n14 ns315 0 -4.13784190211e-05
Gc7_316 0 n14 ns316 0 0.000425260827789
Gc7_317 0 n14 ns317 0 1.23830601849e-05
Gc7_318 0 n14 ns318 0 -0.000323270561268
Gc7_319 0 n14 ns319 0 -0.000233253149562
Gc7_320 0 n14 ns320 0 9.12104168157e-05
Gc7_321 0 n14 ns321 0 -0.000925993055698
Gc7_322 0 n14 ns322 0 0.000296150696139
Gc7_323 0 n14 ns323 0 -0.000506853084971
Gc7_324 0 n14 ns324 0 -0.000610331433908
Gc7_325 0 n14 ns325 0 0.00105044986015
Gc7_326 0 n14 ns326 0 -0.000407070899523
Gc7_327 0 n14 ns327 0 0.00109105418391
Gc7_328 0 n14 ns328 0 -0.00151586446566
Gc7_329 0 n14 ns329 0 0.00122914216183
Gc7_330 0 n14 ns330 0 0.00028892790536
Gc7_331 0 n14 ns331 0 -0.000148889140699
Gc7_332 0 n14 ns332 0 -0.000655184519409
Gc7_333 0 n14 ns333 0 -0.000758791312406
Gc7_334 0 n14 ns334 0 -0.000454951288346
Gc7_335 0 n14 ns335 0 1.88436947587e-05
Gc7_336 0 n14 ns336 0 5.12790787259e-05
Gc7_337 0 n14 ns337 0 0.00376369480684
Gc7_338 0 n14 ns338 0 0.010443251303
Gc7_339 0 n14 ns339 0 -0.00225046599154
Gc7_340 0 n14 ns340 0 -0.000727619630339
Gc7_341 0 n14 ns341 0 3.24445550403e-05
Gc7_342 0 n14 ns342 0 -4.21003885363e-06
Gc7_343 0 n14 ns343 0 0.000114922422112
Gc7_344 0 n14 ns344 0 3.94583341177e-05
Gc7_345 0 n14 ns345 0 5.3850805591e-07
Gc7_346 0 n14 ns346 0 -1.66386055279e-06
Gc7_347 0 n14 ns347 0 -6.67538063912e-05
Gc7_348 0 n14 ns348 0 -5.05808864204e-05
Gc7_349 0 n14 ns349 0 0.000200440035362
Gc7_350 0 n14 ns350 0 5.84775647585e-06
Gc7_351 0 n14 ns351 0 1.92703317225e-06
Gc7_352 0 n14 ns352 0 -1.81534617732e-06
Gc7_353 0 n14 ns353 0 -8.47732318802e-06
Gc7_354 0 n14 ns354 0 6.59506018925e-05
Gc7_355 0 n14 ns355 0 8.33172004527e-06
Gc7_356 0 n14 ns356 0 -0.000163057989016
Gc7_357 0 n14 ns357 0 4.44659446715e-06
Gc7_358 0 n14 ns358 0 3.71337669046e-06
Gc7_359 0 n14 ns359 0 -0.000102397810431
Gc7_360 0 n14 ns360 0 -1.53047610856e-05
Gc7_361 0 n14 ns361 0 9.90481091533e-05
Gc7_362 0 n14 ns362 0 8.12601077878e-05
Gc7_363 0 n14 ns363 0 2.45365892015e-05
Gc7_364 0 n14 ns364 0 -4.26200728394e-06
Gc7_365 0 n14 ns365 0 3.16810289766e-05
Gc7_366 0 n14 ns366 0 -0.000155917135341
Gc7_367 0 n14 ns367 0 0.000168946186247
Gc7_368 0 n14 ns368 0 1.77332046734e-05
Gc7_369 0 n14 ns369 0 0.000205135075661
Gc7_370 0 n14 ns370 0 -5.73914463131e-05
Gc7_371 0 n14 ns371 0 -0.000354973360542
Gc7_372 0 n14 ns372 0 4.52729477254e-05
Gc7_373 0 n14 ns373 0 0.000219052503597
Gc7_374 0 n14 ns374 0 3.28100159534e-05
Gc7_375 0 n14 ns375 0 -0.000103828028446
Gc7_376 0 n14 ns376 0 -0.000339501760431
Gc7_377 0 n14 ns377 0 -0.000614944340065
Gc7_378 0 n14 ns378 0 -0.000331170291144
Gc7_379 0 n14 ns379 0 0.000894201116708
Gc7_380 0 n14 ns380 0 -0.000932697316655
Gc7_381 0 n14 ns381 0 0.000395519690311
Gc7_382 0 n14 ns382 0 0.000529947167568
Gc7_383 0 n14 ns383 0 0.00315972285249
Gc7_384 0 n14 ns384 0 0.000395650060232
Gc7_385 0 n14 ns385 0 -0.000469925132721
Gc7_386 0 n14 ns386 0 0.00379829938977
Gc7_387 0 n14 ns387 0 -0.00103662041012
Gc7_388 0 n14 ns388 0 -0.00156901567406
Gc7_389 0 n14 ns389 0 -0.0108287479204
Gc7_390 0 n14 ns390 0 -0.000578740040604
Gc7_391 0 n14 ns391 0 7.6016597986e-05
Gc7_392 0 n14 ns392 0 0.000129056273913
Gc7_393 0 n14 ns393 0 -0.00153562165934
Gc7_394 0 n14 ns394 0 -0.000706063357609
Gc7_395 0 n14 ns395 0 0.000553834865141
Gc7_396 0 n14 ns396 0 0.0007361129312
Gc7_397 0 n14 ns397 0 2.36001630153e-05
Gc7_398 0 n14 ns398 0 6.90481361042e-06
Gc7_399 0 n14 ns399 0 0.000195113315036
Gc7_400 0 n14 ns400 0 3.39365186451e-05
Gc7_401 0 n14 ns401 0 -8.8331119012e-07
Gc7_402 0 n14 ns402 0 1.17926572787e-06
Gc7_403 0 n14 ns403 0 6.73219896109e-06
Gc7_404 0 n14 ns404 0 0.000152196715301
Gc7_405 0 n14 ns405 0 0.000257245164709
Gc7_406 0 n14 ns406 0 -0.000132006697751
Gc7_407 0 n14 ns407 0 -1.85956399944e-06
Gc7_408 0 n14 ns408 0 -1.47864200372e-07
Gc7_409 0 n14 ns409 0 0.000162435070583
Gc7_410 0 n14 ns410 0 -2.57191639092e-05
Gc7_411 0 n14 ns411 0 -0.000172775204202
Gc7_412 0 n14 ns412 0 -0.000295999866179
Gc7_413 0 n14 ns413 0 2.32250746167e-06
Gc7_414 0 n14 ns414 0 -6.52658273913e-06
Gc7_415 0 n14 ns415 0 -5.95193290676e-05
Gc7_416 0 n14 ns416 0 0.000192800654251
Gc7_417 0 n14 ns417 0 0.000386943512546
Gc7_418 0 n14 ns418 0 0.000206440457623
Gc7_419 0 n14 ns419 0 -1.43821129327e-05
Gc7_420 0 n14 ns420 0 -4.75456912141e-05
Gc7_421 0 n14 ns421 0 4.06518861654e-05
Gc7_422 0 n14 ns422 0 -0.000266512025246
Gc7_423 0 n14 ns423 0 0.000541317123764
Gc7_424 0 n14 ns424 0 -0.000133025371367
Gc7_425 0 n14 ns425 0 0.000737184494363
Gc7_426 0 n14 ns426 0 -5.44873991098e-05
Gc7_427 0 n14 ns427 0 -0.000607941797061
Gc7_428 0 n14 ns428 0 0.000177899602442
Gc7_429 0 n14 ns429 0 0.000593059262668
Gc7_430 0 n14 ns430 0 -0.000193633985942
Gc7_431 0 n14 ns431 0 -0.00021127374439
Gc7_432 0 n14 ns432 0 -0.00024970923639
Gc7_433 0 n14 ns433 0 -0.00114652958518
Gc7_434 0 n14 ns434 0 -0.00100999883403
Gc7_435 0 n14 ns435 0 0.000465401394019
Gc7_436 0 n14 ns436 0 -0.00112037839062
Gc7_437 0 n14 ns437 0 0.00102935680698
Gc7_438 0 n14 ns438 0 0.000651224307164
Gc7_439 0 n14 ns439 0 0.00272583650489
Gc7_440 0 n14 ns440 0 -2.90603041711e-05
Gc7_441 0 n14 ns441 0 0.000626685448127
Gc7_442 0 n14 ns442 0 0.00241203563899
Gc7_443 0 n14 ns443 0 -0.000142373002445
Gc7_444 0 n14 ns444 0 -0.00226532296184
Gc7_445 0 n14 ns445 0 -0.00679027279509
Gc7_446 0 n14 ns446 0 -0.000652365528532
Gc7_447 0 n14 ns447 0 4.34311047487e-05
Gc7_448 0 n14 ns448 0 0.000115106190959
Gd7_1 0 n14 ni1 0 -0.000180797774504
Gd7_2 0 n14 ni2 0 0.000200900219406
Gd7_3 0 n14 ni3 0 -0.000469242499437
Gd7_4 0 n14 ni4 0 -0.000111719103939
Gd7_5 0 n14 ni5 0 0.00314084433507
Gd7_6 0 n14 ni6 0 -0.000942616600776
Gd7_7 0 n14 ni7 0 -0.00410537796466
Gd7_8 0 n14 ni8 0 0.00503269662615
Gc8_1 0 n16 ns1 0 -0.000712931426221
Gc8_2 0 n16 ns2 0 -0.000223358260137
Gc8_3 0 n16 ns3 0 0.000253242670963
Gc8_4 0 n16 ns4 0 0.000131395692981
Gc8_5 0 n16 ns5 0 -2.17049179807e-07
Gc8_6 0 n16 ns6 0 1.61885631188e-05
Gc8_7 0 n16 ns7 0 -3.36215853981e-05
Gc8_8 0 n16 ns8 0 7.3184917099e-05
Gc8_9 0 n16 ns9 0 5.29569681822e-08
Gc8_10 0 n16 ns10 0 1.50543995445e-07
Gc8_11 0 n16 ns11 0 6.45796432919e-05
Gc8_12 0 n16 ns12 0 0.000124457261616
Gc8_13 0 n16 ns13 0 -5.2077929954e-05
Gc8_14 0 n16 ns14 0 -9.00032664717e-05
Gc8_15 0 n16 ns15 0 1.98073985269e-08
Gc8_16 0 n16 ns16 0 -1.33386152891e-06
Gc8_17 0 n16 ns17 0 -9.15320784861e-05
Gc8_18 0 n16 ns18 0 9.72016659897e-05
Gc8_19 0 n16 ns19 0 0.000122148480348
Gc8_20 0 n16 ns20 0 -4.01992033887e-05
Gc8_21 0 n16 ns21 0 -6.61082787787e-06
Gc8_22 0 n16 ns22 0 3.30653707811e-06
Gc8_23 0 n16 ns23 0 1.33372018208e-05
Gc8_24 0 n16 ns24 0 0.000194130193479
Gc8_25 0 n16 ns25 0 9.61872289792e-05
Gc8_26 0 n16 ns26 0 -0.000208595127842
Gc8_27 0 n16 ns27 0 2.74013357683e-05
Gc8_28 0 n16 ns28 0 -3.77953547965e-05
Gc8_29 0 n16 ns29 0 0.000241617504665
Gc8_30 0 n16 ns30 0 0.000157219625825
Gc8_31 0 n16 ns31 0 2.80096800266e-05
Gc8_32 0 n16 ns32 0 0.000131199935019
Gc8_33 0 n16 ns33 0 0.00011152323175
Gc8_34 0 n16 ns34 0 -0.000695226825541
Gc8_35 0 n16 ns35 0 0.00011932066391
Gc8_36 0 n16 ns36 0 0.000189589302567
Gc8_37 0 n16 ns37 0 1.96332232126e-05
Gc8_38 0 n16 ns38 0 0.000366493493125
Gc8_39 0 n16 ns39 0 0.000188975343354
Gc8_40 0 n16 ns40 0 -0.000143574421276
Gc8_41 0 n16 ns41 0 -0.00110363672461
Gc8_42 0 n16 ns42 0 2.04379577608e-05
Gc8_43 0 n16 ns43 0 -0.000646685099737
Gc8_44 0 n16 ns44 0 -0.00033088533168
Gc8_45 0 n16 ns45 0 -0.00128365323436
Gc8_46 0 n16 ns46 0 0.000172293431458
Gc8_47 0 n16 ns47 0 -0.000536367277008
Gc8_48 0 n16 ns48 0 0.000866856702471
Gc8_49 0 n16 ns49 0 0.00142600986769
Gc8_50 0 n16 ns50 0 5.91965389743e-06
Gc8_51 0 n16 ns51 0 0.00110633029078
Gc8_52 0 n16 ns52 0 -0.000247843609871
Gc8_53 0 n16 ns53 0 0.00104576654594
Gc8_54 0 n16 ns54 0 0.000374662247355
Gc8_55 0 n16 ns55 0 -3.40301503826e-05
Gc8_56 0 n16 ns56 0 -1.74253712166e-05
Gc8_57 0 n16 ns57 0 -0.00295379921318
Gc8_58 0 n16 ns58 0 0.000693701074803
Gc8_59 0 n16 ns59 0 -7.51046749846e-05
Gc8_60 0 n16 ns60 0 -0.000152000279319
Gc8_61 0 n16 ns61 0 -2.52961221842e-06
Gc8_62 0 n16 ns62 0 1.66989830265e-05
Gc8_63 0 n16 ns63 0 -0.000108906125952
Gc8_64 0 n16 ns64 0 3.40413580267e-05
Gc8_65 0 n16 ns65 0 -4.40632241701e-06
Gc8_66 0 n16 ns66 0 -4.11234597108e-06
Gc8_67 0 n16 ns67 0 2.00277808649e-06
Gc8_68 0 n16 ns68 0 -0.000182877514127
Gc8_69 0 n16 ns69 0 6.05374153059e-05
Gc8_70 0 n16 ns70 0 -0.000175913019101
Gc8_71 0 n16 ns71 0 4.34129025032e-06
Gc8_72 0 n16 ns72 0 1.08969848294e-05
Gc8_73 0 n16 ns73 0 0.000197481098818
Gc8_74 0 n16 ns74 0 -2.37865591135e-05
Gc8_75 0 n16 ns75 0 0.000192540710448
Gc8_76 0 n16 ns76 0 4.62278374664e-05
Gc8_77 0 n16 ns77 0 2.56829293479e-05
Gc8_78 0 n16 ns78 0 -1.39805222891e-05
Gc8_79 0 n16 ns79 0 8.3077673431e-05
Gc8_80 0 n16 ns80 0 -0.000305734867443
Gc8_81 0 n16 ns81 0 0.000218304794125
Gc8_82 0 n16 ns82 0 -0.000111485568055
Gc8_83 0 n16 ns83 0 -6.73763848359e-05
Gc8_84 0 n16 ns84 0 9.28989097248e-05
Gc8_85 0 n16 ns85 0 -0.000148415445401
Gc8_86 0 n16 ns86 0 -0.000412880142606
Gc8_87 0 n16 ns87 0 -2.44106930994e-05
Gc8_88 0 n16 ns88 0 0.000591866484077
Gc8_89 0 n16 ns89 0 -0.000450190065809
Gc8_90 0 n16 ns90 0 0.000604158455617
Gc8_91 0 n16 ns91 0 5.45609173712e-05
Gc8_92 0 n16 ns92 0 0.000795719444954
Gc8_93 0 n16 ns93 0 -4.9462142295e-05
Gc8_94 0 n16 ns94 0 4.71600308924e-05
Gc8_95 0 n16 ns95 0 0.00052735536975
Gc8_96 0 n16 ns96 0 -1.86236439959e-05
Gc8_97 0 n16 ns97 0 0.000719755677199
Gc8_98 0 n16 ns98 0 -0.000662017711303
Gc8_99 0 n16 ns99 0 -0.000710393857711
Gc8_100 0 n16 ns100 0 -0.000958718854031
Gc8_101 0 n16 ns101 0 -0.000589180403344
Gc8_102 0 n16 ns102 0 7.36928077478e-05
Gc8_103 0 n16 ns103 0 -0.000972448683581
Gc8_104 0 n16 ns104 0 0.00185748353621
Gc8_105 0 n16 ns105 0 0.00222410390496
Gc8_106 0 n16 ns106 0 0.000745962276767
Gc8_107 0 n16 ns107 0 0.00243420023168
Gc8_108 0 n16 ns108 0 5.46325994636e-05
Gc8_109 0 n16 ns109 0 0.00325226534575
Gc8_110 0 n16 ns110 0 0.000424213144134
Gc8_111 0 n16 ns111 0 -6.74321543781e-05
Gc8_112 0 n16 ns112 0 -2.66543724534e-05
Gc8_113 0 n16 ns113 0 -0.0126566620133
Gc8_114 0 n16 ns114 0 0.000587002691496
Gc8_115 0 n16 ns115 0 0.000327554015667
Gc8_116 0 n16 ns116 0 0.000240919951928
Gc8_117 0 n16 ns117 0 -2.12322861238e-05
Gc8_118 0 n16 ns118 0 -9.9698777653e-06
Gc8_119 0 n16 ns119 0 -0.00027359599998
Gc8_120 0 n16 ns120 0 2.85370785676e-06
Gc8_121 0 n16 ns121 0 -1.43453275293e-06
Gc8_122 0 n16 ns122 0 4.95045030185e-07
Gc8_123 0 n16 ns123 0 9.44016142384e-06
Gc8_124 0 n16 ns124 0 0.000207248489219
Gc8_125 0 n16 ns125 0 0.000237308943219
Gc8_126 0 n16 ns126 0 -9.86421628301e-05
Gc8_127 0 n16 ns127 0 3.12230367492e-06
Gc8_128 0 n16 ns128 0 1.7777229601e-06
Gc8_129 0 n16 ns129 0 -0.000192483238813
Gc8_130 0 n16 ns130 0 5.47183974521e-05
Gc8_131 0 n16 ns131 0 0.000120098392374
Gc8_132 0 n16 ns132 0 0.000290141063039
Gc8_133 0 n16 ns133 0 6.18549554561e-06
Gc8_134 0 n16 ns134 0 -5.31317410707e-06
Gc8_135 0 n16 ns135 0 -0.000171641566014
Gc8_136 0 n16 ns136 0 0.000289878027493
Gc8_137 0 n16 ns137 0 0.000328237175726
Gc8_138 0 n16 ns138 0 0.000103471524851
Gc8_139 0 n16 ns139 0 -2.0989515539e-05
Gc8_140 0 n16 ns140 0 4.47168687562e-05
Gc8_141 0 n16 ns141 0 -4.43893501085e-05
Gc8_142 0 n16 ns142 0 0.000650293516069
Gc8_143 0 n16 ns143 0 -0.000317707573997
Gc8_144 0 n16 ns144 0 0.000207694089279
Gc8_145 0 n16 ns145 0 0.00172441835097
Gc8_146 0 n16 ns146 0 0.000681503495561
Gc8_147 0 n16 ns147 0 -0.000142086045049
Gc8_148 0 n16 ns148 0 0.000363354159327
Gc8_149 0 n16 ns149 0 -0.000712647674417
Gc8_150 0 n16 ns150 0 -4.23014757039e-05
Gc8_151 0 n16 ns151 0 0.000336182394663
Gc8_152 0 n16 ns152 0 0.000236908266167
Gc8_153 0 n16 ns153 0 0.00121555011268
Gc8_154 0 n16 ns154 0 -0.00412070795032
Gc8_155 0 n16 ns155 0 -0.000131523276367
Gc8_156 0 n16 ns156 0 -0.0011441239822
Gc8_157 0 n16 ns157 0 0.000863829952996
Gc8_158 0 n16 ns158 0 -0.00245891518196
Gc8_159 0 n16 ns159 0 -5.237848081e-05
Gc8_160 0 n16 ns160 0 0.00126700180796
Gc8_161 0 n16 ns161 0 0.00232120769108
Gc8_162 0 n16 ns162 0 0.00205978310597
Gc8_163 0 n16 ns163 0 0.00321703088527
Gc8_164 0 n16 ns164 0 0.001557041932
Gc8_165 0 n16 ns165 0 0.0044572499043
Gc8_166 0 n16 ns166 0 0.000608645905592
Gc8_167 0 n16 ns167 0 -9.13340247774e-05
Gc8_168 0 n16 ns168 0 -0.000102759872809
Gc8_169 0 n16 ns169 0 -0.0072818810926
Gc8_170 0 n16 ns170 0 -0.00026105177859
Gc8_171 0 n16 ns171 0 -0.000180675953113
Gc8_172 0 n16 ns172 0 -0.00011294149314
Gc8_173 0 n16 ns173 0 -1.74691721534e-05
Gc8_174 0 n16 ns174 0 -3.37310504821e-06
Gc8_175 0 n16 ns175 0 -0.000276117966537
Gc8_176 0 n16 ns176 0 -1.1194070098e-05
Gc8_177 0 n16 ns177 0 4.70813091458e-06
Gc8_178 0 n16 ns178 0 3.53962872535e-06
Gc8_179 0 n16 ns179 0 -2.52656006038e-05
Gc8_180 0 n16 ns180 0 -0.000137408284039
Gc8_181 0 n16 ns181 0 0.000271447600205
Gc8_182 0 n16 ns182 0 -0.000184647018821
Gc8_183 0 n16 ns183 0 -4.60148420083e-06
Gc8_184 0 n16 ns184 0 -1.12467492166e-05
Gc8_185 0 n16 ns185 0 0.000149306481355
Gc8_186 0 n16 ns186 0 -4.92851373839e-05
Gc8_187 0 n16 ns187 0 0.000211021653201
Gc8_188 0 n16 ns188 0 0.000290558220336
Gc8_189 0 n16 ns189 0 -2.73742338546e-05
Gc8_190 0 n16 ns190 0 1.53733677676e-05
Gc8_191 0 n16 ns191 0 -4.42099733636e-06
Gc8_192 0 n16 ns192 0 -0.000231203889782
Gc8_193 0 n16 ns193 0 0.000404388726274
Gc8_194 0 n16 ns194 0 0.000105203404013
Gc8_195 0 n16 ns195 0 5.25300165355e-05
Gc8_196 0 n16 ns196 0 -0.000121145550111
Gc8_197 0 n16 ns197 0 -5.30974320418e-05
Gc8_198 0 n16 ns198 0 -0.000448879800343
Gc8_199 0 n16 ns199 0 -0.000503173278692
Gc8_200 0 n16 ns200 0 8.27212187135e-05
Gc8_201 0 n16 ns201 0 -0.00138548797413
Gc8_202 0 n16 ns202 0 -0.000437845262534
Gc8_203 0 n16 ns203 0 -0.000658862302423
Gc8_204 0 n16 ns204 0 0.000373814586846
Gc8_205 0 n16 ns205 0 0.000339259899971
Gc8_206 0 n16 ns206 0 -2.45639922601e-05
Gc8_207 0 n16 ns207 0 0.000196382155464
Gc8_208 0 n16 ns208 0 0.000325358626371
Gc8_209 0 n16 ns209 0 0.00228124993807
Gc8_210 0 n16 ns210 0 0.00341093218385
Gc8_211 0 n16 ns211 0 0.000636895565195
Gc8_212 0 n16 ns212 0 -0.000933342838952
Gc8_213 0 n16 ns213 0 -1.95595816228e-05
Gc8_214 0 n16 ns214 0 0.00474170560164
Gc8_215 0 n16 ns215 0 -0.00693250401552
Gc8_216 0 n16 ns216 0 0.00196027237683
Gc8_217 0 n16 ns217 0 -0.00179386347399
Gc8_218 0 n16 ns218 0 0.00441396679507
Gc8_219 0 n16 ns219 0 -0.00512712888688
Gc8_220 0 n16 ns220 0 -0.0046671774312
Gc8_221 0 n16 ns221 0 0.0197696627967
Gc8_222 0 n16 ns222 0 -0.000394635414651
Gc8_223 0 n16 ns223 0 9.46216350685e-05
Gc8_224 0 n16 ns224 0 7.08981930218e-05
Gc8_225 0 n16 ns225 0 0.0227365214075
Gc8_226 0 n16 ns226 0 0.000247378320382
Gc8_227 0 n16 ns227 0 0.000313788744131
Gc8_228 0 n16 ns228 0 0.000215630048132
Gc8_229 0 n16 ns229 0 -1.14431823593e-05
Gc8_230 0 n16 ns230 0 -1.45995894223e-05
Gc8_231 0 n16 ns231 0 0.000115106637709
Gc8_232 0 n16 ns232 0 -8.77357744424e-05
Gc8_233 0 n16 ns233 0 -4.32657780366e-07
Gc8_234 0 n16 ns234 0 1.29293228568e-08
Gc8_235 0 n16 ns235 0 4.19293569849e-05
Gc8_236 0 n16 ns236 0 8.14266777137e-05
Gc8_237 0 n16 ns237 0 2.24701742898e-06
Gc8_238 0 n16 ns238 0 -0.000149844149455
Gc8_239 0 n16 ns239 0 -2.72824980403e-07
Gc8_240 0 n16 ns240 0 4.9391635236e-07
Gc8_241 0 n16 ns241 0 9.66569157172e-05
Gc8_242 0 n16 ns242 0 -6.61819271759e-05
Gc8_243 0 n16 ns243 0 -0.000161356398651
Gc8_244 0 n16 ns244 0 3.54533308095e-06
Gc8_245 0 n16 ns245 0 -4.54366231885e-06
Gc8_246 0 n16 ns246 0 1.68703472485e-06
Gc8_247 0 n16 ns247 0 1.85555338018e-05
Gc8_248 0 n16 ns248 0 0.00017660208973
Gc8_249 0 n16 ns249 0 0.000123014767639
Gc8_250 0 n16 ns250 0 -0.000129393962373
Gc8_251 0 n16 ns251 0 -2.99104632235e-05
Gc8_252 0 n16 ns252 0 2.13579707124e-05
Gc8_253 0 n16 ns253 0 -0.000201547424284
Gc8_254 0 n16 ns254 0 -0.000198620196603
Gc8_255 0 n16 ns255 0 2.45217562501e-05
Gc8_256 0 n16 ns256 0 -0.000297053824282
Gc8_257 0 n16 ns257 0 -2.75147429941e-06
Gc8_258 0 n16 ns258 0 -0.000474067807276
Gc8_259 0 n16 ns259 0 -4.0660463757e-05
Gc8_260 0 n16 ns260 0 0.000425780462988
Gc8_261 0 n16 ns261 0 1.17405433533e-05
Gc8_262 0 n16 ns262 0 -0.00032293412736
Gc8_263 0 n16 ns263 0 -0.000233358808442
Gc8_264 0 n16 ns264 0 9.15934153485e-05
Gc8_265 0 n16 ns265 0 -0.000925182504986
Gc8_266 0 n16 ns266 0 0.00029787947525
Gc8_267 0 n16 ns267 0 -0.000507788254183
Gc8_268 0 n16 ns268 0 -0.000609890295118
Gc8_269 0 n16 ns269 0 0.00104990269462
Gc8_270 0 n16 ns270 0 -0.000407413213655
Gc8_271 0 n16 ns271 0 0.00108942210754
Gc8_272 0 n16 ns272 0 -0.0015164172412
Gc8_273 0 n16 ns273 0 0.00123083947997
Gc8_274 0 n16 ns274 0 0.00028884407828
Gc8_275 0 n16 ns275 0 -0.000147656578384
Gc8_276 0 n16 ns276 0 -0.000657355022901
Gc8_277 0 n16 ns277 0 -0.000757790881066
Gc8_278 0 n16 ns278 0 -0.000455333631425
Gc8_279 0 n16 ns279 0 1.88773037387e-05
Gc8_280 0 n16 ns280 0 5.13816408162e-05
Gc8_281 0 n16 ns281 0 0.0161650918141
Gc8_282 0 n16 ns282 0 -0.00290362729975
Gc8_283 0 n16 ns283 0 -0.000319130087495
Gc8_284 0 n16 ns284 0 0.00100250096451
Gc8_285 0 n16 ns285 0 4.00041896348e-08
Gc8_286 0 n16 ns286 0 -9.72270391619e-06
Gc8_287 0 n16 ns287 0 0.000114966999602
Gc8_288 0 n16 ns288 0 -9.76686798829e-06
Gc8_289 0 n16 ns289 0 -3.18432208732e-06
Gc8_290 0 n16 ns290 0 -2.35010145354e-06
Gc8_291 0 n16 ns291 0 -1.35670141801e-05
Gc8_292 0 n16 ns292 0 -0.000156161425566
Gc8_293 0 n16 ns293 0 8.21871206096e-05
Gc8_294 0 n16 ns294 0 -0.00016172793601
Gc8_295 0 n16 ns295 0 -2.49894773185e-06
Gc8_296 0 n16 ns296 0 -7.01697253243e-06
Gc8_297 0 n16 ns297 0 -0.000163593151404
Gc8_298 0 n16 ns298 0 1.90201102899e-05
Gc8_299 0 n16 ns299 0 -0.000152498428013
Gc8_300 0 n16 ns300 0 -8.08000598635e-05
Gc8_301 0 n16 ns301 0 2.00095671095e-05
Gc8_302 0 n16 ns302 0 -9.54630651434e-06
Gc8_303 0 n16 ns303 0 8.79358961304e-05
Gc8_304 0 n16 ns304 0 -0.000191934085154
Gc8_305 0 n16 ns305 0 0.000159558626521
Gc8_306 0 n16 ns306 0 -1.69195207374e-05
Gc8_307 0 n16 ns307 0 4.23993324417e-05
Gc8_308 0 n16 ns308 0 -0.000100934272113
Gc8_309 0 n16 ns309 0 -0.000150818776524
Gc8_310 0 n16 ns310 0 0.000446834485076
Gc8_311 0 n16 ns311 0 0.000158376407244
Gc8_312 0 n16 ns312 0 -9.99722830273e-05
Gc8_313 0 n16 ns313 0 -0.000317690731157
Gc8_314 0 n16 ns314 0 0.000121201417921
Gc8_315 0 n16 ns315 0 -1.41554714899e-05
Gc8_316 0 n16 ns316 0 0.000313529367133
Gc8_317 0 n16 ns317 0 -6.38325016644e-05
Gc8_318 0 n16 ns318 0 -9.10021048353e-05
Gc8_319 0 n16 ns319 0 -0.000302764318602
Gc8_320 0 n16 ns320 0 -3.04048861126e-05
Gc8_321 0 n16 ns321 0 -0.000487522424806
Gc8_322 0 n16 ns322 0 0.000714327604533
Gc8_323 0 n16 ns323 0 -0.000439537708625
Gc8_324 0 n16 ns324 0 -0.000774678346804
Gc8_325 0 n16 ns325 0 0.00087204511857
Gc8_326 0 n16 ns326 0 -6.33653961069e-05
Gc8_327 0 n16 ns327 0 0.00150325257659
Gc8_328 0 n16 ns328 0 -0.00125391135665
Gc8_329 0 n16 ns329 0 0.00114268843959
Gc8_330 0 n16 ns330 0 0.00115250479168
Gc8_331 0 n16 ns331 0 -0.000215626493978
Gc8_332 0 n16 ns332 0 -0.00129621488256
Gc8_333 0 n16 ns333 0 -0.00352822860981
Gc8_334 0 n16 ns334 0 -0.000541468982342
Gc8_335 0 n16 ns335 0 4.33081647765e-05
Gc8_336 0 n16 ns336 0 7.31844871493e-05
Gc8_337 0 n16 ns337 0 -0.00153561164918
Gc8_338 0 n16 ns338 0 -0.000706063632338
Gc8_339 0 n16 ns339 0 0.000553833915496
Gc8_340 0 n16 ns340 0 0.00073611314981
Gc8_341 0 n16 ns341 0 2.36001574532e-05
Gc8_342 0 n16 ns342 0 6.90485503821e-06
Gc8_343 0 n16 ns343 0 0.000195113456392
Gc8_344 0 n16 ns344 0 3.39363807131e-05
Gc8_345 0 n16 ns345 0 -8.83311857631e-07
Gc8_346 0 n16 ns346 0 1.17926841616e-06
Gc8_347 0 n16 ns347 0 6.73216368296e-06
Gc8_348 0 n16 ns348 0 0.000152196678249
Gc8_349 0 n16 ns349 0 0.000257245220337
Gc8_350 0 n16 ns350 0 -0.000132006714398
Gc8_351 0 n16 ns351 0 -1.85956649497e-06
Gc8_352 0 n16 ns352 0 -1.47861762853e-07
Gc8_353 0 n16 ns353 0 0.000162435010881
Gc8_354 0 n16 ns354 0 -2.57191981301e-05
Gc8_355 0 n16 ns355 0 -0.00017277520197
Gc8_356 0 n16 ns356 0 -0.000295999944648
Gc8_357 0 n16 ns357 0 2.32250381805e-06
Gc8_358 0 n16 ns358 0 -6.5265852893e-06
Gc8_359 0 n16 ns359 0 -5.95192654013e-05
Gc8_360 0 n16 ns360 0 0.000192800638168
Gc8_361 0 n16 ns361 0 0.000386943490607
Gc8_362 0 n16 ns362 0 0.000206440601093
Gc8_363 0 n16 ns363 0 -1.43821431293e-05
Gc8_364 0 n16 ns364 0 -4.75457147666e-05
Gc8_365 0 n16 ns365 0 4.0651755033e-05
Gc8_366 0 n16 ns366 0 -0.000266511741187
Gc8_367 0 n16 ns367 0 0.000541317213097
Gc8_368 0 n16 ns368 0 -0.000133025306993
Gc8_369 0 n16 ns369 0 0.000737183990166
Gc8_370 0 n16 ns370 0 -5.4487401363e-05
Gc8_371 0 n16 ns371 0 -0.000607941962424
Gc8_372 0 n16 ns372 0 0.000177900024529
Gc8_373 0 n16 ns373 0 0.000593058868568
Gc8_374 0 n16 ns374 0 -0.000193633689299
Gc8_375 0 n16 ns375 0 -0.000211274156264
Gc8_376 0 n16 ns376 0 -0.000249709589021
Gc8_377 0 n16 ns377 0 -0.00114652818762
Gc8_378 0 n16 ns378 0 -0.00100999903253
Gc8_379 0 n16 ns379 0 0.000465402612647
Gc8_380 0 n16 ns380 0 -0.00112037929413
Gc8_381 0 n16 ns381 0 0.00102935589661
Gc8_382 0 n16 ns382 0 0.000651223981341
Gc8_383 0 n16 ns383 0 0.00272583673419
Gc8_384 0 n16 ns384 0 -2.90610026469e-05
Gc8_385 0 n16 ns385 0 0.00062668462751
Gc8_386 0 n16 ns386 0 0.00241203669733
Gc8_387 0 n16 ns387 0 -0.00014237489682
Gc8_388 0 n16 ns388 0 -0.00226532127631
Gc8_389 0 n16 ns389 0 -0.00679027441178
Gc8_390 0 n16 ns390 0 -0.000652365321145
Gc8_391 0 n16 ns391 0 4.34311436712e-05
Gc8_392 0 n16 ns392 0 0.000115106007717
Gc8_393 0 n16 ns393 0 0.0152292354101
Gc8_394 0 n16 ns394 0 0.010242371916
Gc8_395 0 n16 ns395 0 -0.00245576054964
Gc8_396 0 n16 ns396 0 -0.000976302730069
Gc8_397 0 n16 ns397 0 2.23858149761e-05
Gc8_398 0 n16 ns398 0 -1.32071903009e-05
Gc8_399 0 n16 ns399 0 0.000180041490108
Gc8_400 0 n16 ns400 0 -9.56987349682e-06
Gc8_401 0 n16 ns401 0 3.75458178223e-06
Gc8_402 0 n16 ns402 0 1.38112564851e-06
Gc8_403 0 n16 ns403 0 -1.977246105e-05
Gc8_404 0 n16 ns404 0 -4.93547597954e-05
Gc8_405 0 n16 ns405 0 0.000177817780296
Gc8_406 0 n16 ns406 0 -7.21962930361e-05
Gc8_407 0 n16 ns407 0 3.68500317495e-06
Gc8_408 0 n16 ns408 0 5.07567971731e-06
Gc8_409 0 n16 ns409 0 1.94928775904e-05
Gc8_410 0 n16 ns410 0 2.38402430828e-06
Gc8_411 0 n16 ns411 0 -6.82391353871e-05
Gc8_412 0 n16 ns412 0 -0.000114026327413
Gc8_413 0 n16 ns413 0 -1.27633295874e-05
Gc8_414 0 n16 ns414 0 1.04538317619e-05
Gc8_415 0 n16 ns415 0 -4.62831366788e-05
Gc8_416 0 n16 ns416 0 9.05473436554e-05
Gc8_417 0 n16 ns417 0 0.000112091405771
Gc8_418 0 n16 ns418 0 -6.13027868498e-05
Gc8_419 0 n16 ns419 0 -2.32270033229e-05
Gc8_420 0 n16 ns420 0 5.11592834533e-05
Gc8_421 0 n16 ns421 0 -0.000205799399779
Gc8_422 0 n16 ns422 0 -0.000316686512197
Gc8_423 0 n16 ns423 0 0.000101025756779
Gc8_424 0 n16 ns424 0 -0.000231052287892
Gc8_425 0 n16 ns425 0 7.12669489114e-06
Gc8_426 0 n16 ns426 0 -0.000575654825555
Gc8_427 0 n16 ns427 0 -0.000286877323753
Gc8_428 0 n16 ns428 0 0.00039617336701
Gc8_429 0 n16 ns429 0 2.15370879504e-05
Gc8_430 0 n16 ns430 0 -0.000223661870213
Gc8_431 0 n16 ns431 0 -0.000238668057355
Gc8_432 0 n16 ns432 0 -0.000203439453578
Gc8_433 0 n16 ns433 0 -0.00109466625691
Gc8_434 0 n16 ns434 0 0.000256091634326
Gc8_435 0 n16 ns435 0 0.000342586765356
Gc8_436 0 n16 ns436 0 -0.000989948742085
Gc8_437 0 n16 ns437 0 0.00084295096225
Gc8_438 0 n16 ns438 0 -1.27235721377e-05
Gc8_439 0 n16 ns439 0 0.00305422806197
Gc8_440 0 n16 ns440 0 -0.000488796213562
Gc8_441 0 n16 ns441 0 -0.000123652557955
Gc8_442 0 n16 ns442 0 0.00327015801057
Gc8_443 0 n16 ns443 0 -0.00134740247786
Gc8_444 0 n16 ns444 0 -0.00156952902344
Gc8_445 0 n16 ns445 0 -0.0100647142319
Gc8_446 0 n16 ns446 0 -0.000505677820917
Gc8_447 0 n16 ns447 0 6.29080302293e-05
Gc8_448 0 n16 ns448 0 6.68306271e-05
Gd8_1 0 n16 ni1 0 0.000202728832348
Gd8_2 0 n16 ni2 0 -0.000463497343493
Gd8_3 0 n16 ni3 0 -0.000112621890281
Gd8_4 0 n16 ni4 0 9.77695158038e-05
Gd8_5 0 n16 ni5 0 -0.000942875307866
Gd8_6 0 n16 ni6 0 0.00386417962443
Gd8_7 0 n16 ni7 0 0.00503269664391
Gd8_8 0 n16 ni8 0 -0.00579818317536
.ends m4linesveryHighFreq_HFSS_100mil_fws
