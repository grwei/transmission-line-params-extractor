* begin ansoft header
* node 1 Diff1
* node 2 Comm1
* node 3 trace_p_1_T1
* node 4 trace_n_1_T1
* node 5 Diff2
* node 6 Comm2
* node 7 trace_p_1_T2
* node 8 trace_n_1_T2
* 
* created by ElectronicsDesktop
* end ansoft header

.subckt m4lines_HFSS_lfws 1 2 3 4 5 6 7 8 
v5_1 5 9 dc 0.0
v6_2 6 10 dc 0.0
v7_3 7 11 dc 0.0
v8_4 8 12 dc 0.0
rl1_5to1 9 13 3835.3354425521
ls1_5to1 13 1 234.38199300545n
rs2_5to1 9 14 0.045833372916536
ls2_5to1 14 1 2.1215070299218n
rl1_6to2 10 15 3500.0117127773
ls1_6to2 15 2 231.45957130715n
rs2_6to2 10 16 0.046414385774099
ls2_6to2 16 2 2.1074169538709n
rl1_7to3 11 17 4310.7987941295
ls1_7to3 17 3 237.479062293n
rs2_7to3 11 18 0.045433748286339
ls2_7to3 18 3 2.1224558692175n
rl1_8to4 12 19 3551.1037170345
ls1_8to4 19 4 231.59202743085n
rs2_8to4 12 20 0.046388645670636
ls2_8to4 20 4 2.106954193598n
rc1_1to0 1 21 1e-05
cs1_1to0 21 0 0.051848691793394p
rp_1to0 1 0 103376.12245141
rc1_5to0 5 22 1e-05
cs1_5to0 22 0 0.051182998384235p
rp_5to0 5 0 102306.63005705
rc1_2to0 2 23 1e-05
cs1_2to0 23 0 0.080266896914659p
rp_2to0 2 0 111221.07360796
rc1_6to0 6 24 1e-05
cs1_6to0 24 0 0.07981233438926p
rp_6to0 6 0 115445.73322451
rc1_3to0 3 25 1e-05
cs1_3to0 25 0 0.049364606183987p
rp_3to0 3 0 102287.96150766
rc1_7to0 7 26 1e-05
cs1_7to0 26 0 0.048759294971844p
rp_7to0 7 0 104006.12269259
rc1_4to0 4 27 1e-05
cs1_4to0 27 0 0.028734848403042p
rp_4to0 4 0 113143.93592502
rc1_8to0 8 28 1e-05
cs1_8to0 28 0 0.028291393055291p
rp_8to0 8 0 113448.17667139
f5to1_6to2b1 15 2 v5_1 0.0071197563183946
f5to1_6to2b2 16 2 v5_1 -0.3638884550589
f6to2_5to1b1 13 1 v6_2 0.0072539370697742
f6to2_5to1b2 14 1 v6_2 -0.36150394671169
f5to1_7to3b1 17 3 v5_1 0.001371700769288
f5to1_7to3b2 18 3 v5_1 -0.060495256504794
f7to3_5to1b1 13 1 v7_3 0.0013244669012531
f7to3_5to1b2 14 1 v7_3 -0.060514636880718
f5to1_8to4b1 19 4 v5_1 0.0026524105244988
f5to1_8to4b2 20 4 v5_1 -0.11125821644144
f8to4_5to1b1 13 1 v8_4 0.0027016973874664
f8to4_5to1b2 14 1 v8_4 -0.11050615624767
f6to2_7to3b1 17 3 v6_2 0.0028425237434578
f6to2_7to3b2 18 3 v6_2 -0.11047901374462
f7to3_6to2b1 15 2 v7_3 0.0026600452861052
f7to3_6to2b2 16 2 v7_3 -0.11123704712977
f6to2_8to4b1 19 4 v6_2 0.0069850136190426
f6to2_8to4b2 20 4 v6_2 -0.22546969225303
f8to4_6to2b1 15 2 v8_4 0.0069360925450015
f8to4_6to2b2 16 2 v8_4 -0.22541304041666
f7to3_8to4b1 19 4 v7_3 0.0071444254646874
f7to3_8to4b2 20 4 v7_3 -0.36408123832714
f8to4_7to3b1 17 3 v8_4 0.0074959363885776
f8to4_7to3b2 18 3 v8_4 -0.36148652477251
cm_1to29 1 29 0.10732380005767p
cm_5to29 5 29 0.10732380005767p
cm_29to2 29 2 0.10732380005767p
cm_29to6 29 6 0.10732380005767p
cm_1to30 1 30 0.10732380005767p
cm_5to30 5 30 0.10732380005767p
cm_30to3 30 3 0.10732380005767p
cm_30to7 30 7 0.10732380005767p
cm_1to31 1 31 0.10732380005767p
cm_5to31 5 31 0.10732380005767p
cm_31to4 31 4 0.10732380005767p
cm_31to8 31 8 0.10732380005767p
cm_2to32 2 32 0.0042043094643768p
cm_6to32 6 32 0.0042043094643768p
cm_32to3 32 3 0.0042043094643768p
cm_32to7 32 7 0.0042043094643768p
cm_2to33 2 33 0.0042043094643768p
cm_6to33 6 33 0.0042043094643768p
cm_33to4 33 4 0.0042043094643768p
cm_33to8 33 8 0.0042043094643768p
cm_3to34 3 34 0.1073449840084p
cm_7to34 7 34 0.1073449840084p
cm_34to4 34 4 0.1073449840084p
cm_34to8 34 8 0.1073449840084p
.ends m4lines_HFSS_lfws

