* begin ansoft header
* node 1 Diff1
* node 2 Comm1
* node 3 trace_p_1_T1
* node 4 trace_n_1_T1
* node 5 Diff2
* node 6 Comm2
* node 7 trace_p_1_T2
* node 8 trace_n_1_T2
* 
* created by ElectronicsDesktop
* end ansoft header

.subckt m4lines_veryHighFreq_lfws 1 2 3 4 5 6 7 8 
v5_1 5 9 dc 0.0
v6_2 6 10 dc 0.0
v7_3 7 11 dc 0.0
v8_4 8 12 dc 0.0
rl1_5to1 9 13 0.09983015052918
ls1_5to1 13 1 1.0874380320888n
rl1_6to2 10 14 0.1013583226084
ls1_6to2 14 2 1.0786916204276n
rl1_7to3 11 15 0.10018608179236
ls1_7to3 15 3 1.0872197412239n
rl1_8to4 12 16 0.1012183218269
ls1_8to4 16 4 1.0787539957967n
rc1_1to0 1 17 1e-05
cs1_1to0 17 0 0.00058473468156642p
rp_1to0 1 0 46921.599621906
rc1_5to0 5 18 1e-05
cs1_5to0 18 0 0.00050064481975569p
rp_5to0 5 0 47451.238437414
rc1_2to0 2 19 1e-05
cs1_2to0 19 0 0.040559496873679p
rp_2to0 2 0 52225.813923077
rc1_6to0 6 20 1e-05
cs1_6to0 20 0 0.040486254665818p
rp_6to0 6 0 52966.953536199
rc1_3to0 3 21 1e-05
cs1_3to0 21 0 0.025577859334706p
rp_3to0 3 0 46837.465603273
rc1_7to0 7 22 1e-05
cs1_7to0 22 0 0.025492081212892p
rp_7to0 7 0 47588.136216363
rc1_4to0 4 23 1e-05
cs1_4to0 23 0 0.015562424004516p
rp_4to0 4 0 52103.572685355
rc1_8to0 8 24 1e-05
cs1_8to0 24 0 0.015500686630428p
rp_8to0 8 0 53011.303069945
cm_1to25 1 25 0.051921464308808p
cm_5to25 5 25 0.051921464308808p
cm_25to2 25 2 0.051921464308808p
cm_25to6 25 6 0.051921464308808p
cm_1to26 1 26 0.051921464308808p
cm_5to26 5 26 0.051921464308808p
cm_26to3 26 3 0.051921464308808p
cm_26to7 26 7 0.051921464308808p
cm_1to27 1 27 0.051921464308808p
cm_5to27 5 27 0.051921464308808p
cm_27to4 27 4 0.051921464308808p
cm_27to8 27 8 0.051921464308808p
cm_2to28 2 28 0.0019120486183093p
cm_6to28 6 28 0.0019120486183093p
cm_28to3 28 3 0.0019120486183093p
cm_28to7 28 7 0.0019120486183093p
cm_2to29 2 29 0.0019120486183093p
cm_6to29 6 29 0.0019120486183093p
cm_29to4 29 4 0.0019120486183093p
cm_29to8 29 8 0.0019120486183093p
cm_3to30 3 30 0.051916353373613p
cm_7to30 7 30 0.051916353373613p
cm_30to4 30 4 0.051916353373613p
cm_30to8 30 8 0.051916353373613p
.ends m4lines_veryHighFreq_lfws

