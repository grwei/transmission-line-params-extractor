* BEGIN ANSOFT HEADER
* node 1    trace_p_0_T1
* node 2    trace_n_0_T1
* node 3    trace_p_1_T1
* node 4    trace_n_1_T1
* node 5    trace_p_0_T2
* node 6    trace_n_0_T2
* node 7    trace_p_1_T2
* node 8    trace_n_1_T2
*   Format: HSPICE
*   Topckt: m4lines_port_fws
*     Date: Sat Jun 06 09:41:15 2020
*    Notes: Frequency range: 0 to 7e+10 Hz, 701 points
*         : Maximum number of poles: 10000
*         : S-Matrix fitting error tolerance: 0.001
*         : Causality check tolerance: auto
*         : Passivity enforcement: on (by iterated fitting)
*         : Causality enforcement: off
*         : Fitting method: FastFit
*         : Matrix fitting: By entire matrix (required by FastFit)
*         : Ensure Z-parameter accuracy: on
*         : Relative error control: off
*         : Common ground option: on
*         : Final fitting error: 0.00473093
*         : Final model order: 104
* END ANSOFT HEADER

.subckt m4lines_port_fws 1 2 3 4 5 6 7 8
Vam1 1 n2 dc 0
Rport1 n2 0 50 noise=0
Vam2 2 n4 dc 0
Rport2 n4 0 50 noise=0
Vam3 3 n6 dc 0
Rport3 n6 0 50 noise=0
Vam4 4 n8 dc 0
Rport4 n8 0 50 noise=0
Vam5 5 n10 dc 0
Rport5 n10 0 50 noise=0
Vam6 6 n12 dc 0
Rport6 n12 0 50 noise=0
Vam7 7 n14 dc 0
Rport7 n14 0 50 noise=0
Vam8 8 n16 dc 0
Rport8 n16 0 50 noise=0

Fi1 0 ni1 Vam1 50
Gi1 0 ni1 1 0 1
Rt1 ni1 0 1 noise=0
Fi2 0 ni2 Vam2 50
Gi2 0 ni2 2 0 1
Rt2 ni2 0 1 noise=0
Fi3 0 ni3 Vam3 50
Gi3 0 ni3 3 0 1
Rt3 ni3 0 1 noise=0
Fi4 0 ni4 Vam4 50
Gi4 0 ni4 4 0 1
Rt4 ni4 0 1 noise=0
Fi5 0 ni5 Vam5 50
Gi5 0 ni5 5 0 1
Rt5 ni5 0 1 noise=0
Fi6 0 ni6 Vam6 50
Gi6 0 ni6 6 0 1
Rt6 ni6 0 1 noise=0
Fi7 0 ni7 Vam7 50
Gi7 0 ni7 7 0 1
Rt7 ni7 0 1 noise=0
Fi8 0 ni8 Vam8 50
Gi8 0 ni8 8 0 1
Rt8 ni8 0 1 noise=0

Ca1 ns1 0 1e-12
Ca2 ns2 0 1e-12
Ra1 ns1 0 3.94856876484 noise=0
Ra2 ns2 0 3.94856876484 noise=0
Ga1 ns1 0 ns2 0 -2.15302669132
Ga2 ns2 0 ns1 0 2.15302669132
Ca3 ns3 0 1e-12
Ca4 ns4 0 1e-12
Ra3 ns3 0 15.0340813991 noise=0
Ra4 ns4 0 15.0340813991 noise=0
Ga3 ns3 0 ns4 0 -1.15977236587
Ga4 ns4 0 ns3 0 1.15977236587
Ca5 ns5 0 1e-12
Ca6 ns6 0 1e-12
Ra5 ns5 0 1.57905702417 noise=0
Ra6 ns6 0 1.57905702417 noise=0
Ga5 ns5 0 ns6 0 -0.228371344881
Ga6 ns6 0 ns5 0 0.228371344881
Ca7 ns7 0 1e-12
Ca8 ns8 0 1e-12
Ra7 ns7 0 6.93869622444 noise=0
Ra8 ns8 0 6.93869622444 noise=0
Ga7 ns7 0 ns8 0 -0.166818924494
Ga8 ns8 0 ns7 0 0.166818924494
Ca9 ns9 0 1e-12
Ca10 ns10 0 1e-12
Ra9 ns9 0 105.254899829 noise=0
Ra10 ns10 0 105.254899829 noise=0
Ga9 ns9 0 ns10 0 -0.00215881551475
Ga10 ns10 0 ns9 0 0.00215881551475
Ca11 ns11 0 1e-12
Ra11 ns11 0 1278.30041043 noise=0
Ca12 ns12 0 1e-12
Ra12 ns12 0 33983.3277547 noise=0
Ca13 ns13 0 1e-12
Ra13 ns13 0 23276.0424715 noise=0
Ca14 ns14 0 1e-12
Ca15 ns15 0 1e-12
Ra14 ns14 0 3.94856876484 noise=0
Ra15 ns15 0 3.94856876484 noise=0
Ga14 ns14 0 ns15 0 -2.15302669132
Ga15 ns15 0 ns14 0 2.15302669132
Ca16 ns16 0 1e-12
Ca17 ns17 0 1e-12
Ra16 ns16 0 15.0340813991 noise=0
Ra17 ns17 0 15.0340813991 noise=0
Ga16 ns16 0 ns17 0 -1.15977236587
Ga17 ns17 0 ns16 0 1.15977236587
Ca18 ns18 0 1e-12
Ca19 ns19 0 1e-12
Ra18 ns18 0 1.57905702417 noise=0
Ra19 ns19 0 1.57905702417 noise=0
Ga18 ns18 0 ns19 0 -0.228371344881
Ga19 ns19 0 ns18 0 0.228371344881
Ca20 ns20 0 1e-12
Ca21 ns21 0 1e-12
Ra20 ns20 0 6.93869622444 noise=0
Ra21 ns21 0 6.93869622444 noise=0
Ga20 ns20 0 ns21 0 -0.166818924494
Ga21 ns21 0 ns20 0 0.166818924494
Ca22 ns22 0 1e-12
Ca23 ns23 0 1e-12
Ra22 ns22 0 105.254899829 noise=0
Ra23 ns23 0 105.254899829 noise=0
Ga22 ns22 0 ns23 0 -0.00215881551475
Ga23 ns23 0 ns22 0 0.00215881551475
Ca24 ns24 0 1e-12
Ra24 ns24 0 1278.30041043 noise=0
Ca25 ns25 0 1e-12
Ra25 ns25 0 33983.3277547 noise=0
Ca26 ns26 0 1e-12
Ra26 ns26 0 23276.0424715 noise=0
Ca27 ns27 0 1e-12
Ca28 ns28 0 1e-12
Ra27 ns27 0 3.94856876484 noise=0
Ra28 ns28 0 3.94856876484 noise=0
Ga27 ns27 0 ns28 0 -2.15302669132
Ga28 ns28 0 ns27 0 2.15302669132
Ca29 ns29 0 1e-12
Ca30 ns30 0 1e-12
Ra29 ns29 0 15.0340813991 noise=0
Ra30 ns30 0 15.0340813991 noise=0
Ga29 ns29 0 ns30 0 -1.15977236587
Ga30 ns30 0 ns29 0 1.15977236587
Ca31 ns31 0 1e-12
Ca32 ns32 0 1e-12
Ra31 ns31 0 1.57905702417 noise=0
Ra32 ns32 0 1.57905702417 noise=0
Ga31 ns31 0 ns32 0 -0.228371344881
Ga32 ns32 0 ns31 0 0.228371344881
Ca33 ns33 0 1e-12
Ca34 ns34 0 1e-12
Ra33 ns33 0 6.93869622444 noise=0
Ra34 ns34 0 6.93869622444 noise=0
Ga33 ns33 0 ns34 0 -0.166818924494
Ga34 ns34 0 ns33 0 0.166818924494
Ca35 ns35 0 1e-12
Ca36 ns36 0 1e-12
Ra35 ns35 0 105.254899829 noise=0
Ra36 ns36 0 105.254899829 noise=0
Ga35 ns35 0 ns36 0 -0.00215881551475
Ga36 ns36 0 ns35 0 0.00215881551475
Ca37 ns37 0 1e-12
Ra37 ns37 0 1278.30041043 noise=0
Ca38 ns38 0 1e-12
Ra38 ns38 0 33983.3277547 noise=0
Ca39 ns39 0 1e-12
Ra39 ns39 0 23276.0424715 noise=0
Ca40 ns40 0 1e-12
Ca41 ns41 0 1e-12
Ra40 ns40 0 3.94856876484 noise=0
Ra41 ns41 0 3.94856876484 noise=0
Ga40 ns40 0 ns41 0 -2.15302669132
Ga41 ns41 0 ns40 0 2.15302669132
Ca42 ns42 0 1e-12
Ca43 ns43 0 1e-12
Ra42 ns42 0 15.0340813991 noise=0
Ra43 ns43 0 15.0340813991 noise=0
Ga42 ns42 0 ns43 0 -1.15977236587
Ga43 ns43 0 ns42 0 1.15977236587
Ca44 ns44 0 1e-12
Ca45 ns45 0 1e-12
Ra44 ns44 0 1.57905702417 noise=0
Ra45 ns45 0 1.57905702417 noise=0
Ga44 ns44 0 ns45 0 -0.228371344881
Ga45 ns45 0 ns44 0 0.228371344881
Ca46 ns46 0 1e-12
Ca47 ns47 0 1e-12
Ra46 ns46 0 6.93869622444 noise=0
Ra47 ns47 0 6.93869622444 noise=0
Ga46 ns46 0 ns47 0 -0.166818924494
Ga47 ns47 0 ns46 0 0.166818924494
Ca48 ns48 0 1e-12
Ca49 ns49 0 1e-12
Ra48 ns48 0 105.254899829 noise=0
Ra49 ns49 0 105.254899829 noise=0
Ga48 ns48 0 ns49 0 -0.00215881551475
Ga49 ns49 0 ns48 0 0.00215881551475
Ca50 ns50 0 1e-12
Ra50 ns50 0 1278.30041043 noise=0
Ca51 ns51 0 1e-12
Ra51 ns51 0 33983.3277547 noise=0
Ca52 ns52 0 1e-12
Ra52 ns52 0 23276.0424715 noise=0
Ca53 ns53 0 1e-12
Ca54 ns54 0 1e-12
Ra53 ns53 0 3.94856876484 noise=0
Ra54 ns54 0 3.94856876484 noise=0
Ga53 ns53 0 ns54 0 -2.15302669132
Ga54 ns54 0 ns53 0 2.15302669132
Ca55 ns55 0 1e-12
Ca56 ns56 0 1e-12
Ra55 ns55 0 15.0340813991 noise=0
Ra56 ns56 0 15.0340813991 noise=0
Ga55 ns55 0 ns56 0 -1.15977236587
Ga56 ns56 0 ns55 0 1.15977236587
Ca57 ns57 0 1e-12
Ca58 ns58 0 1e-12
Ra57 ns57 0 1.57905702417 noise=0
Ra58 ns58 0 1.57905702417 noise=0
Ga57 ns57 0 ns58 0 -0.228371344881
Ga58 ns58 0 ns57 0 0.228371344881
Ca59 ns59 0 1e-12
Ca60 ns60 0 1e-12
Ra59 ns59 0 6.93869622444 noise=0
Ra60 ns60 0 6.93869622444 noise=0
Ga59 ns59 0 ns60 0 -0.166818924494
Ga60 ns60 0 ns59 0 0.166818924494
Ca61 ns61 0 1e-12
Ca62 ns62 0 1e-12
Ra61 ns61 0 105.254899829 noise=0
Ra62 ns62 0 105.254899829 noise=0
Ga61 ns61 0 ns62 0 -0.00215881551475
Ga62 ns62 0 ns61 0 0.00215881551475
Ca63 ns63 0 1e-12
Ra63 ns63 0 1278.30041043 noise=0
Ca64 ns64 0 1e-12
Ra64 ns64 0 33983.3277547 noise=0
Ca65 ns65 0 1e-12
Ra65 ns65 0 23276.0424715 noise=0
Ca66 ns66 0 1e-12
Ca67 ns67 0 1e-12
Ra66 ns66 0 3.94856876484 noise=0
Ra67 ns67 0 3.94856876484 noise=0
Ga66 ns66 0 ns67 0 -2.15302669132
Ga67 ns67 0 ns66 0 2.15302669132
Ca68 ns68 0 1e-12
Ca69 ns69 0 1e-12
Ra68 ns68 0 15.0340813991 noise=0
Ra69 ns69 0 15.0340813991 noise=0
Ga68 ns68 0 ns69 0 -1.15977236587
Ga69 ns69 0 ns68 0 1.15977236587
Ca70 ns70 0 1e-12
Ca71 ns71 0 1e-12
Ra70 ns70 0 1.57905702417 noise=0
Ra71 ns71 0 1.57905702417 noise=0
Ga70 ns70 0 ns71 0 -0.228371344881
Ga71 ns71 0 ns70 0 0.228371344881
Ca72 ns72 0 1e-12
Ca73 ns73 0 1e-12
Ra72 ns72 0 6.93869622444 noise=0
Ra73 ns73 0 6.93869622444 noise=0
Ga72 ns72 0 ns73 0 -0.166818924494
Ga73 ns73 0 ns72 0 0.166818924494
Ca74 ns74 0 1e-12
Ca75 ns75 0 1e-12
Ra74 ns74 0 105.254899829 noise=0
Ra75 ns75 0 105.254899829 noise=0
Ga74 ns74 0 ns75 0 -0.00215881551475
Ga75 ns75 0 ns74 0 0.00215881551475
Ca76 ns76 0 1e-12
Ra76 ns76 0 1278.30041043 noise=0
Ca77 ns77 0 1e-12
Ra77 ns77 0 33983.3277547 noise=0
Ca78 ns78 0 1e-12
Ra78 ns78 0 23276.0424715 noise=0
Ca79 ns79 0 1e-12
Ca80 ns80 0 1e-12
Ra79 ns79 0 3.94856876484 noise=0
Ra80 ns80 0 3.94856876484 noise=0
Ga79 ns79 0 ns80 0 -2.15302669132
Ga80 ns80 0 ns79 0 2.15302669132
Ca81 ns81 0 1e-12
Ca82 ns82 0 1e-12
Ra81 ns81 0 15.0340813991 noise=0
Ra82 ns82 0 15.0340813991 noise=0
Ga81 ns81 0 ns82 0 -1.15977236587
Ga82 ns82 0 ns81 0 1.15977236587
Ca83 ns83 0 1e-12
Ca84 ns84 0 1e-12
Ra83 ns83 0 1.57905702417 noise=0
Ra84 ns84 0 1.57905702417 noise=0
Ga83 ns83 0 ns84 0 -0.228371344881
Ga84 ns84 0 ns83 0 0.228371344881
Ca85 ns85 0 1e-12
Ca86 ns86 0 1e-12
Ra85 ns85 0 6.93869622444 noise=0
Ra86 ns86 0 6.93869622444 noise=0
Ga85 ns85 0 ns86 0 -0.166818924494
Ga86 ns86 0 ns85 0 0.166818924494
Ca87 ns87 0 1e-12
Ca88 ns88 0 1e-12
Ra87 ns87 0 105.254899829 noise=0
Ra88 ns88 0 105.254899829 noise=0
Ga87 ns87 0 ns88 0 -0.00215881551475
Ga88 ns88 0 ns87 0 0.00215881551475
Ca89 ns89 0 1e-12
Ra89 ns89 0 1278.30041043 noise=0
Ca90 ns90 0 1e-12
Ra90 ns90 0 33983.3277547 noise=0
Ca91 ns91 0 1e-12
Ra91 ns91 0 23276.0424715 noise=0
Ca92 ns92 0 1e-12
Ca93 ns93 0 1e-12
Ra92 ns92 0 3.94856876484 noise=0
Ra93 ns93 0 3.94856876484 noise=0
Ga92 ns92 0 ns93 0 -2.15302669132
Ga93 ns93 0 ns92 0 2.15302669132
Ca94 ns94 0 1e-12
Ca95 ns95 0 1e-12
Ra94 ns94 0 15.0340813991 noise=0
Ra95 ns95 0 15.0340813991 noise=0
Ga94 ns94 0 ns95 0 -1.15977236587
Ga95 ns95 0 ns94 0 1.15977236587
Ca96 ns96 0 1e-12
Ca97 ns97 0 1e-12
Ra96 ns96 0 1.57905702417 noise=0
Ra97 ns97 0 1.57905702417 noise=0
Ga96 ns96 0 ns97 0 -0.228371344881
Ga97 ns97 0 ns96 0 0.228371344881
Ca98 ns98 0 1e-12
Ca99 ns99 0 1e-12
Ra98 ns98 0 6.93869622444 noise=0
Ra99 ns99 0 6.93869622444 noise=0
Ga98 ns98 0 ns99 0 -0.166818924494
Ga99 ns99 0 ns98 0 0.166818924494
Ca100 ns100 0 1e-12
Ca101 ns101 0 1e-12
Ra100 ns100 0 105.254899829 noise=0
Ra101 ns101 0 105.254899829 noise=0
Ga100 ns100 0 ns101 0 -0.00215881551475
Ga101 ns101 0 ns100 0 0.00215881551475
Ca102 ns102 0 1e-12
Ra102 ns102 0 1278.30041043 noise=0
Ca103 ns103 0 1e-12
Ra103 ns103 0 33983.3277547 noise=0
Ca104 ns104 0 1e-12
Ra104 ns104 0 23276.0424715 noise=0

Gb1_1 ns1 0 ni1 0 2.18281673738
Gb3_1 ns3 0 ni1 0 1.16358718058
Gb5_1 ns5 0 ni1 0 0.715642657222
Gb7_1 ns7 0 ni1 0 0.291327405282
Gb9_1 ns9 0 ni1 0 0.00999128417038
Gb11_1 ns11 0 ni1 0 0.000782288726372
Gb12_1 ns12 0 ni1 0 2.9426194139e-05
Gb13_1 ns13 0 ni1 0 4.29626299757e-05
Gb14_2 ns14 0 ni2 0 2.18281673738
Gb16_2 ns16 0 ni2 0 1.16358718058
Gb18_2 ns18 0 ni2 0 0.715642657222
Gb20_2 ns20 0 ni2 0 0.291327405282
Gb22_2 ns22 0 ni2 0 0.00999128417038
Gb24_2 ns24 0 ni2 0 0.000782288726372
Gb25_2 ns25 0 ni2 0 2.9426194139e-05
Gb26_2 ns26 0 ni2 0 4.29626299757e-05
Gb27_3 ns27 0 ni3 0 2.18281673738
Gb29_3 ns29 0 ni3 0 1.16358718058
Gb31_3 ns31 0 ni3 0 0.715642657222
Gb33_3 ns33 0 ni3 0 0.291327405282
Gb35_3 ns35 0 ni3 0 0.00999128417038
Gb37_3 ns37 0 ni3 0 0.000782288726372
Gb38_3 ns38 0 ni3 0 2.9426194139e-05
Gb39_3 ns39 0 ni3 0 4.29626299757e-05
Gb40_4 ns40 0 ni4 0 2.18281673738
Gb42_4 ns42 0 ni4 0 1.16358718058
Gb44_4 ns44 0 ni4 0 0.715642657222
Gb46_4 ns46 0 ni4 0 0.291327405282
Gb48_4 ns48 0 ni4 0 0.00999128417038
Gb50_4 ns50 0 ni4 0 0.000782288726372
Gb51_4 ns51 0 ni4 0 2.9426194139e-05
Gb52_4 ns52 0 ni4 0 4.29626299757e-05
Gb53_5 ns53 0 ni5 0 2.18281673738
Gb55_5 ns55 0 ni5 0 1.16358718058
Gb57_5 ns57 0 ni5 0 0.715642657222
Gb59_5 ns59 0 ni5 0 0.291327405282
Gb61_5 ns61 0 ni5 0 0.00999128417038
Gb63_5 ns63 0 ni5 0 0.000782288726372
Gb64_5 ns64 0 ni5 0 2.9426194139e-05
Gb65_5 ns65 0 ni5 0 4.29626299757e-05
Gb66_6 ns66 0 ni6 0 2.18281673738
Gb68_6 ns68 0 ni6 0 1.16358718058
Gb70_6 ns70 0 ni6 0 0.715642657222
Gb72_6 ns72 0 ni6 0 0.291327405282
Gb74_6 ns74 0 ni6 0 0.00999128417038
Gb76_6 ns76 0 ni6 0 0.000782288726372
Gb77_6 ns77 0 ni6 0 2.9426194139e-05
Gb78_6 ns78 0 ni6 0 4.29626299757e-05
Gb79_7 ns79 0 ni7 0 2.18281673738
Gb81_7 ns81 0 ni7 0 1.16358718058
Gb83_7 ns83 0 ni7 0 0.715642657222
Gb85_7 ns85 0 ni7 0 0.291327405282
Gb87_7 ns87 0 ni7 0 0.00999128417038
Gb89_7 ns89 0 ni7 0 0.000782288726372
Gb90_7 ns90 0 ni7 0 2.9426194139e-05
Gb91_7 ns91 0 ni7 0 4.29626299757e-05
Gb92_8 ns92 0 ni8 0 2.18281673738
Gb94_8 ns94 0 ni8 0 1.16358718058
Gb96_8 ns96 0 ni8 0 0.715642657222
Gb98_8 ns98 0 ni8 0 0.291327405282
Gb100_8 ns100 0 ni8 0 0.00999128417038
Gb102_8 ns102 0 ni8 0 0.000782288726372
Gb103_8 ns103 0 ni8 0 2.9426194139e-05
Gb104_8 ns104 0 ni8 0 4.29626299757e-05

Gc1_1 0 n2 ns1 0 0.00142908116134
Gc1_2 0 n2 ns2 0 0.0022905132688
Gc1_3 0 n2 ns3 0 0.000112455606693
Gc1_4 0 n2 ns4 0 0.0016564851108
Gc1_5 0 n2 ns5 0 -0.000560756694312
Gc1_6 0 n2 ns6 0 -0.00364601948029
Gc1_7 0 n2 ns7 0 -0.000141354140526
Gc1_8 0 n2 ns8 0 0.000158637408551
Gc1_9 0 n2 ns9 0 7.95596836179e-05
Gc1_10 0 n2 ns10 0 0.000140997228753
Gc1_11 0 n2 ns11 0 4.14341393047e-05
Gc1_12 0 n2 ns12 0 -0.00155949874459
Gc1_13 0 n2 ns13 0 -0.000552351274449
Gc1_14 0 n2 ns14 0 0.000460678773102
Gc1_15 0 n2 ns15 0 0.000722310903946
Gc1_16 0 n2 ns16 0 6.2468769393e-05
Gc1_17 0 n2 ns17 0 0.000473677597114
Gc1_18 0 n2 ns18 0 -0.0014635964679
Gc1_19 0 n2 ns19 0 -0.00349880635773
Gc1_20 0 n2 ns20 0 -9.25504629169e-05
Gc1_21 0 n2 ns21 0 0.000137382289662
Gc1_22 0 n2 ns22 0 -2.71215137064e-05
Gc1_23 0 n2 ns23 0 -0.000230495608075
Gc1_24 0 n2 ns24 0 -3.23071877914e-06
Gc1_25 0 n2 ns25 0 0.000699337402706
Gc1_26 0 n2 ns26 0 -6.73853434182e-06
Gc1_27 0 n2 ns27 0 1.27608207765e-07
Gc1_28 0 n2 ns28 0 -2.19326656994e-05
Gc1_29 0 n2 ns29 0 8.73381953777e-06
Gc1_30 0 n2 ns30 0 -9.04684507887e-05
Gc1_31 0 n2 ns31 0 2.51159785081e-05
Gc1_32 0 n2 ns32 0 -0.000236035831447
Gc1_33 0 n2 ns33 0 -0.000122847599685
Gc1_34 0 n2 ns34 0 -1.91054997556e-05
Gc1_35 0 n2 ns35 0 -1.32977690873e-05
Gc1_36 0 n2 ns36 0 -2.61574101869e-05
Gc1_37 0 n2 ns37 0 -6.39664123488e-06
Gc1_38 0 n2 ns38 0 3.19896234991e-05
Gc1_39 0 n2 ns39 0 1.29656244228e-05
Gc1_40 0 n2 ns40 0 8.77224188209e-07
Gc1_41 0 n2 ns41 0 -1.89544899371e-05
Gc1_42 0 n2 ns42 0 1.5864566019e-05
Gc1_43 0 n2 ns43 0 -6.76305394117e-05
Gc1_44 0 n2 ns44 0 -0.000396446796065
Gc1_45 0 n2 ns45 0 -0.000669114664956
Gc1_46 0 n2 ns46 0 -4.1430638989e-05
Gc1_47 0 n2 ns47 0 -3.81842347673e-05
Gc1_48 0 n2 ns48 0 -1.1594242694e-06
Gc1_49 0 n2 ns49 0 -1.29567694664e-05
Gc1_50 0 n2 ns50 0 3.55493987626e-06
Gc1_51 0 n2 ns51 0 5.29263364952e-05
Gc1_52 0 n2 ns52 0 2.73400442002e-05
Gd1_1 0 n2 ni1 0 -0.000318840485699
Gd1_2 0 n2 ni2 0 0.00155079635812
Gd1_3 0 n2 ni3 0 0.00031217807293
Gd1_4 0 n2 ni4 0 0.000378821848244
Gc2_1 0 n4 ns1 0 0.000460678773104
Gc2_2 0 n4 ns2 0 0.000722310903949
Gc2_3 0 n4 ns3 0 6.2468769393e-05
Gc2_4 0 n4 ns4 0 0.000473677597116
Gc2_5 0 n4 ns5 0 -0.0014635964679
Gc2_6 0 n4 ns6 0 -0.00349880635772
Gc2_7 0 n4 ns7 0 -9.25504629171e-05
Gc2_8 0 n4 ns8 0 0.000137382289662
Gc2_9 0 n4 ns9 0 -2.71215137066e-05
Gc2_10 0 n4 ns10 0 -0.000230495608076
Gc2_11 0 n4 ns11 0 -3.23071877922e-06
Gc2_12 0 n4 ns12 0 0.000699337402708
Gc2_13 0 n4 ns13 0 -6.7385343407e-06
Gc2_14 0 n4 ns14 0 0.000391932179398
Gc2_15 0 n4 ns15 0 0.000553692705588
Gc2_16 0 n4 ns16 0 9.40269584415e-05
Gc2_17 0 n4 ns17 0 0.000373181185777
Gc2_18 0 n4 ns18 0 -0.00143380958801
Gc2_19 0 n4 ns19 0 -0.00374107828263
Gc2_20 0 n4 ns20 0 -0.000132666895209
Gc2_21 0 n4 ns21 0 0.00013622568566
Gc2_22 0 n4 ns22 0 7.60454397694e-05
Gc2_23 0 n4 ns23 0 0.000134230823901
Gc2_24 0 n4 ns24 0 3.62553772766e-05
Gc2_25 0 n4 ns25 0 -0.00150025341666
Gc2_26 0 n4 ns26 0 -0.000709850438285
Gc2_27 0 n4 ns27 0 -5.27467593374e-06
Gc2_28 0 n4 ns28 0 -3.00632972555e-05
Gc2_29 0 n4 ns29 0 1.59270237533e-05
Gc2_30 0 n4 ns30 0 -7.72816514678e-05
Gc2_31 0 n4 ns31 0 -0.000408032275591
Gc2_32 0 n4 ns32 0 -0.000681169942292
Gc2_33 0 n4 ns33 0 -4.12047858561e-05
Gc2_34 0 n4 ns34 0 -3.73414995513e-05
Gc2_35 0 n4 ns35 0 -1.4160041418e-06
Gc2_36 0 n4 ns36 0 -1.40157996613e-05
Gc2_37 0 n4 ns37 0 3.42421863686e-06
Gc2_38 0 n4 ns38 0 5.43051980909e-05
Gc2_39 0 n4 ns39 0 2.62321805886e-05
Gc2_40 0 n4 ns40 0 0.000596263656179
Gc2_41 0 n4 ns41 0 0.000976197202738
Gc2_42 0 n4 ns42 0 4.5147570942e-05
Gc2_43 0 n4 ns43 0 0.00069415807517
Gc2_44 0 n4 ns44 0 -0.000359760418821
Gc2_45 0 n4 ns45 0 -0.00162028756761
Gc2_46 0 n4 ns46 0 -5.67988174773e-05
Gc2_47 0 n4 ns47 0 7.00648970754e-05
Gc2_48 0 n4 ns48 0 -2.35340035969e-06
Gc2_49 0 n4 ns49 0 -7.11803008347e-05
Gc2_50 0 n4 ns50 0 2.54917273766e-06
Gc2_51 0 n4 ns51 0 0.000221805669356
Gc2_52 0 n4 ns52 0 1.39712782548e-05
Gd2_1 0 n4 ni1 0 0.00155079635812
Gd2_2 0 n4 ni2 0 0.00152966184128
Gd2_3 0 n4 ni3 0 0.000390900306215
Gd2_4 0 n4 ni4 0 0.000132027691434
Gc3_1 0 n6 ns1 0 1.27608207868e-07
Gc3_2 0 n6 ns2 0 -2.19326656993e-05
Gc3_3 0 n6 ns3 0 8.73381953779e-06
Gc3_4 0 n6 ns4 0 -9.04684507887e-05
Gc3_5 0 n6 ns5 0 2.5115978508e-05
Gc3_6 0 n6 ns6 0 -0.000236035831447
Gc3_7 0 n6 ns7 0 -0.000122847599685
Gc3_8 0 n6 ns8 0 -1.91054997556e-05
Gc3_9 0 n6 ns9 0 -1.32977690873e-05
Gc3_10 0 n6 ns10 0 -2.6157410187e-05
Gc3_11 0 n6 ns11 0 -6.39664123489e-06
Gc3_12 0 n6 ns12 0 3.19896234992e-05
Gc3_13 0 n6 ns13 0 1.29656244228e-05
Gc3_14 0 n6 ns14 0 -5.27467593377e-06
Gc3_15 0 n6 ns15 0 -3.00632972555e-05
Gc3_16 0 n6 ns16 0 1.59270237533e-05
Gc3_17 0 n6 ns17 0 -7.72816514677e-05
Gc3_18 0 n6 ns18 0 -0.000408032275591
Gc3_19 0 n6 ns19 0 -0.000681169942292
Gc3_20 0 n6 ns20 0 -4.12047858561e-05
Gc3_21 0 n6 ns21 0 -3.73414995513e-05
Gc3_22 0 n6 ns22 0 -1.4160041418e-06
Gc3_23 0 n6 ns23 0 -1.40157996613e-05
Gc3_24 0 n6 ns24 0 3.42421863686e-06
Gc3_25 0 n6 ns25 0 5.43051980909e-05
Gc3_26 0 n6 ns26 0 2.62321805886e-05
Gc3_27 0 n6 ns27 0 0.00144994570026
Gc3_28 0 n6 ns28 0 0.00232349159503
Gc3_29 0 n6 ns29 0 0.000113463552268
Gc3_30 0 n6 ns30 0 0.00167654198341
Gc3_31 0 n6 ns31 0 -0.000548387013357
Gc3_32 0 n6 ns32 0 -0.00365396180048
Gc3_33 0 n6 ns33 0 -0.000141542506546
Gc3_34 0 n6 ns34 0 0.000160057934679
Gc3_35 0 n6 ns35 0 7.88198494583e-05
Gc3_36 0 n6 ns36 0 0.000138721785731
Gc3_37 0 n6 ns37 0 4.12614353032e-05
Gc3_38 0 n6 ns38 0 -0.00156156266205
Gc3_39 0 n6 ns39 0 -0.000547671429107
Gc3_40 0 n6 ns40 0 0.000452174365459
Gc3_41 0 n6 ns41 0 0.000706907480471
Gc3_42 0 n6 ns42 0 6.32136528224e-05
Gc3_43 0 n6 ns43 0 0.000459458903986
Gc3_44 0 n6 ns44 0 -0.00147935421517
Gc3_45 0 n6 ns45 0 -0.0035236273904
Gc3_46 0 n6 ns46 0 -9.49489811671e-05
Gc3_47 0 n6 ns47 0 0.00013875550719
Gc3_48 0 n6 ns48 0 -2.81286376733e-05
Gc3_49 0 n6 ns49 0 -0.000234245401501
Gc3_50 0 n6 ns50 0 -3.67414702326e-06
Gc3_51 0 n6 ns51 0 0.000706918743806
Gc3_52 0 n6 ns52 0 -7.28686185714e-06
Gd3_1 0 n6 ni1 0 0.00031217807293
Gd3_2 0 n6 ni2 0 0.000390900306215
Gd3_3 0 n6 ni3 0 -0.000367670605914
Gd3_4 0 n6 ni4 0 0.00157883341718
Gc4_1 0 n8 ns1 0 8.77224188028e-07
Gc4_2 0 n8 ns2 0 -1.89544899374e-05
Gc4_3 0 n8 ns3 0 1.5864566019e-05
Gc4_4 0 n8 ns4 0 -6.76305394118e-05
Gc4_5 0 n8 ns5 0 -0.000396446796065
Gc4_6 0 n8 ns6 0 -0.000669114664956
Gc4_7 0 n8 ns7 0 -4.14306389889e-05
Gc4_8 0 n8 ns8 0 -3.81842347673e-05
Gc4_9 0 n8 ns9 0 -1.15942426939e-06
Gc4_10 0 n8 ns10 0 -1.29567694664e-05
Gc4_11 0 n8 ns11 0 3.55493987627e-06
Gc4_12 0 n8 ns12 0 5.2926336495e-05
Gc4_13 0 n8 ns13 0 2.73400442001e-05
Gc4_14 0 n8 ns14 0 0.000596263656178
Gc4_15 0 n8 ns15 0 0.000976197202737
Gc4_16 0 n8 ns16 0 4.5147570942e-05
Gc4_17 0 n8 ns17 0 0.000694158075169
Gc4_18 0 n8 ns18 0 -0.000359760418821
Gc4_19 0 n8 ns19 0 -0.00162028756761
Gc4_20 0 n8 ns20 0 -5.67988174773e-05
Gc4_21 0 n8 ns21 0 7.00648970753e-05
Gc4_22 0 n8 ns22 0 -2.35340035965e-06
Gc4_23 0 n8 ns23 0 -7.11803008346e-05
Gc4_24 0 n8 ns24 0 2.54917273768e-06
Gc4_25 0 n8 ns25 0 0.000221805669355
Gc4_26 0 n8 ns26 0 1.39712782545e-05
Gc4_27 0 n8 ns27 0 0.000452174365458
Gc4_28 0 n8 ns28 0 0.000706907480468
Gc4_29 0 n8 ns29 0 6.32136528225e-05
Gc4_30 0 n8 ns30 0 0.000459458903984
Gc4_31 0 n8 ns31 0 -0.00147935421517
Gc4_32 0 n8 ns32 0 -0.0035236273904
Gc4_33 0 n8 ns33 0 -9.49489811669e-05
Gc4_34 0 n8 ns34 0 0.00013875550719
Gc4_35 0 n8 ns35 0 -2.81286376732e-05
Gc4_36 0 n8 ns36 0 -0.000234245401501
Gc4_37 0 n8 ns37 0 -3.6741470232e-06
Gc4_38 0 n8 ns38 0 0.000706918743803
Gc4_39 0 n8 ns39 0 -7.28686185809e-06
Gc4_40 0 n8 ns40 0 0.000394111116324
Gc4_41 0 n8 ns41 0 0.000556786785427
Gc4_42 0 n8 ns42 0 9.47206494839e-05
Gc4_43 0 n8 ns43 0 0.000374793721417
Gc4_44 0 n8 ns44 0 -0.00143765336387
Gc4_45 0 n8 ns45 0 -0.00374783371063
Gc4_46 0 n8 ns46 0 -0.0001315816592
Gc4_47 0 n8 ns47 0 0.000135911834894
Gc4_48 0 n8 ns48 0 7.62068495299e-05
Gc4_49 0 n8 ns49 0 0.000134695615131
Gc4_50 0 n8 ns50 0 3.64439012873e-05
Gc4_51 0 n8 ns51 0 -0.0015070076413
Gc4_52 0 n8 ns52 0 -0.000710021944524
Gd4_1 0 n8 ni1 0 0.000378821848244
Gd4_2 0 n8 ni2 0 0.000132027691435
Gd4_3 0 n8 ni3 0 0.00157883341718
Gd4_4 0 n8 ni4 0 0.00151868695176
Gc5_53 0 n10 ns53 0 0.0014503478784
Gc5_54 0 n10 ns54 0 0.00231852238807
Gc5_55 0 n10 ns55 0 0.000115129784089
Gc5_56 0 n10 ns56 0 0.00166100110303
Gc5_57 0 n10 ns57 0 -0.00057567224741
Gc5_58 0 n10 ns58 0 -0.00371149057077
Gc5_59 0 n10 ns59 0 -0.000144720161698
Gc5_60 0 n10 ns60 0 0.000163297708185
Gc5_61 0 n10 ns61 0 7.73059844458e-05
Gc5_62 0 n10 ns62 0 0.000134130877019
Gc5_63 0 n10 ns63 0 4.06164675499e-05
Gc5_64 0 n10 ns64 0 -0.00156371254318
Gc5_65 0 n10 ns65 0 -0.00054771870641
Gc5_66 0 n10 ns66 0 0.000474926753124
Gc5_67 0 n10 ns67 0 0.000741927677524
Gc5_68 0 n10 ns68 0 6.55830754716e-05
Gc5_69 0 n10 ns69 0 0.00047913219028
Gc5_70 0 n10 ns70 0 -0.00147500822441
Gc5_71 0 n10 ns71 0 -0.00354597921792
Gc5_72 0 n10 ns72 0 -9.44378649205e-05
Gc5_73 0 n10 ns73 0 0.000140528300831
Gc5_74 0 n10 ns74 0 -2.8311959023e-05
Gc5_75 0 n10 ns75 0 -0.000234206016483
Gc5_76 0 n10 ns76 0 -3.69875276906e-06
Gc5_77 0 n10 ns77 0 0.000696389219673
Gc5_78 0 n10 ns78 0 -4.62921696222e-06
Gc5_79 0 n10 ns79 0 -2.29514471368e-06
Gc5_80 0 n10 ns80 0 -2.77530201331e-05
Gc5_81 0 n10 ns81 0 9.3031863334e-06
Gc5_82 0 n10 ns82 0 -9.82787155188e-05
Gc5_83 0 n10 ns83 0 3.44917460449e-06
Gc5_84 0 n10 ns84 0 -0.000261726390453
Gc5_85 0 n10 ns85 0 -0.000121197204833
Gc5_86 0 n10 ns86 0 -1.9466700696e-05
Gc5_87 0 n10 ns87 0 -1.29658839357e-05
Gc5_88 0 n10 ns88 0 -2.51069710757e-05
Gc5_89 0 n10 ns89 0 -6.16034299039e-06
Gc5_90 0 n10 ns90 0 3.11073737759e-05
Gc5_91 0 n10 ns91 0 1.34579731369e-05
Gc5_92 0 n10 ns92 0 7.63371248757e-06
Gc5_93 0 n10 ns93 0 -1.03386931621e-05
Gc5_94 0 n10 ns94 0 1.70118546675e-05
Gc5_95 0 n10 ns95 0 -6.69174069355e-05
Gc5_96 0 n10 ns96 0 -0.00041133510426
Gc5_97 0 n10 ns97 0 -0.000698733322723
Gc5_98 0 n10 ns98 0 -4.05792279847e-05
Gc5_99 0 n10 ns99 0 -3.71465337128e-05
Gc5_100 0 n10 ns100 0 -1.23189660534e-06
Gc5_101 0 n10 ns101 0 -1.30982242138e-05
Gc5_102 0 n10 ns102 0 3.5342796233e-06
Gc5_103 0 n10 ns103 0 5.13641247967e-05
Gc5_104 0 n10 ns104 0 2.84462664288e-05
Gd5_5 0 n10 ni5 0 -0.000367506116176
Gd5_6 0 n10 ni6 0 0.00152366847592
Gd5_7 0 n10 ni7 0 0.000315138206101
Gd5_8 0 n10 ni8 0 0.000365460831507
Gc6_53 0 n12 ns53 0 0.000474926753123
Gc6_54 0 n12 ns54 0 0.000741927677522
Gc6_55 0 n12 ns55 0 6.55830754716e-05
Gc6_56 0 n12 ns56 0 0.000479132190278
Gc6_57 0 n12 ns57 0 -0.00147500822441
Gc6_58 0 n12 ns58 0 -0.00354597921792
Gc6_59 0 n12 ns59 0 -9.44378649204e-05
Gc6_60 0 n12 ns60 0 0.000140528300831
Gc6_61 0 n12 ns61 0 -2.83119590229e-05
Gc6_62 0 n12 ns62 0 -0.000234206016483
Gc6_63 0 n12 ns63 0 -3.69875276901e-06
Gc6_64 0 n12 ns64 0 0.000696389219671
Gc6_65 0 n12 ns65 0 -4.62921696299e-06
Gc6_66 0 n12 ns66 0 0.000395528997379
Gc6_67 0 n12 ns67 0 0.000557551835303
Gc6_68 0 n12 ns68 0 9.65773296643e-05
Gc6_69 0 n12 ns69 0 0.000371180623308
Gc6_70 0 n12 ns70 0 -0.00144866742984
Gc6_71 0 n12 ns71 0 -0.00377969574137
Gc6_72 0 n12 ns72 0 -0.000135017941545
Gc6_73 0 n12 ns73 0 0.00013762810402
Gc6_74 0 n12 ns74 0 7.54295769786e-05
Gc6_75 0 n12 ns75 0 0.000132136181885
Gc6_76 0 n12 ns76 0 3.60022481713e-05
Gc6_77 0 n12 ns77 0 -0.00149996179362
Gc6_78 0 n12 ns78 0 -0.000709750454606
Gc6_79 0 n12 ns79 0 -2.78056574248e-06
Gc6_80 0 n12 ns80 0 -2.57935407088e-05
Gc6_81 0 n12 ns81 0 1.64583240608e-05
Gc6_82 0 n12 ns82 0 -7.42110039877e-05
Gc6_83 0 n12 ns83 0 -0.000404974649941
Gc6_84 0 n12 ns84 0 -0.000678408061432
Gc6_85 0 n12 ns85 0 -4.10889402543e-05
Gc6_86 0 n12 ns86 0 -3.7447001912e-05
Gc6_87 0 n12 ns87 0 -1.14599772015e-06
Gc6_88 0 n12 ns88 0 -1.27455947247e-05
Gc6_89 0 n12 ns89 0 3.45914346117e-06
Gc6_90 0 n12 ns90 0 5.35493792521e-05
Gc6_91 0 n12 ns91 0 2.63367125031e-05
Gc6_92 0 n12 ns92 0 0.000592652286888
Gc6_93 0 n12 ns93 0 0.000968960244026
Gc6_94 0 n12 ns94 0 4.59426853158e-05
Gc6_95 0 n12 ns95 0 0.000686193579921
Gc6_96 0 n12 ns96 0 -0.000371918092218
Gc6_97 0 n12 ns97 0 -0.00163531086767
Gc6_98 0 n12 ns98 0 -5.66934403148e-05
Gc6_99 0 n12 ns99 0 7.0540258634e-05
Gc6_100 0 n12 ns100 0 -2.40540694012e-06
Gc6_101 0 n12 ns101 0 -7.11082409398e-05
Gc6_102 0 n12 ns102 0 2.45823275746e-06
Gc6_103 0 n12 ns103 0 0.000222025945237
Gc6_104 0 n12 ns104 0 1.33820096123e-05
Gd6_5 0 n12 ni5 0 0.00152366847592
Gd6_6 0 n12 ni6 0 0.00153419193007
Gd6_7 0 n12 ni7 0 0.000385794457698
Gd6_8 0 n12 ni8 0 0.000138868871671
Gc7_53 0 n14 ns53 0 -2.29514471376e-06
Gc7_54 0 n14 ns54 0 -2.77530201332e-05
Gc7_55 0 n14 ns55 0 9.3031863334e-06
Gc7_56 0 n14 ns56 0 -9.82787155188e-05
Gc7_57 0 n14 ns57 0 3.44917460443e-06
Gc7_58 0 n14 ns58 0 -0.000261726390453
Gc7_59 0 n14 ns59 0 -0.000121197204833
Gc7_60 0 n14 ns60 0 -1.9466700696e-05
Gc7_61 0 n14 ns61 0 -1.29658839357e-05
Gc7_62 0 n14 ns62 0 -2.51069710756e-05
Gc7_63 0 n14 ns63 0 -6.16034299038e-06
Gc7_64 0 n14 ns64 0 3.11073737758e-05
Gc7_65 0 n14 ns65 0 1.34579731369e-05
Gc7_66 0 n14 ns66 0 -2.78056574232e-06
Gc7_67 0 n14 ns67 0 -2.57935407086e-05
Gc7_68 0 n14 ns68 0 1.64583240607e-05
Gc7_69 0 n14 ns69 0 -7.42110039876e-05
Gc7_70 0 n14 ns70 0 -0.000404974649941
Gc7_71 0 n14 ns71 0 -0.000678408061432
Gc7_72 0 n14 ns72 0 -4.10889402543e-05
Gc7_73 0 n14 ns73 0 -3.7447001912e-05
Gc7_74 0 n14 ns74 0 -1.14599772016e-06
Gc7_75 0 n14 ns75 0 -1.27455947248e-05
Gc7_76 0 n14 ns76 0 3.45914346116e-06
Gc7_77 0 n14 ns77 0 5.35493792523e-05
Gc7_78 0 n14 ns78 0 2.63367125032e-05
Gc7_79 0 n14 ns79 0 0.00142516887178
Gc7_80 0 n14 ns80 0 0.00228570015596
Gc7_81 0 n14 ns81 0 0.000111985332131
Gc7_82 0 n14 ns82 0 0.00165652964641
Gc7_83 0 n14 ns83 0 -0.000555093088213
Gc7_84 0 n14 ns84 0 -0.00362324974229
Gc7_85 0 n14 ns85 0 -0.000138830654793
Gc7_86 0 n14 ns86 0 0.000157703340721
Gc7_87 0 n14 ns87 0 8.03133507718e-05
Gc7_88 0 n14 ns88 0 0.000143740600683
Gc7_89 0 n14 ns89 0 4.16532195795e-05
Gc7_90 0 n14 ns90 0 -0.00155850277643
Gc7_91 0 n14 ns91 0 -0.000552664830265
Gc7_92 0 n14 ns92 0 0.000464549364354
Gc7_93 0 n14 ns93 0 0.000729546096376
Gc7_94 0 n14 ns94 0 6.21067673478e-05
Gc7_95 0 n14 ns95 0 0.000479841897054
Gc7_96 0 n14 ns96 0 -0.0014489874963
Gc7_97 0 n14 ns97 0 -0.00348468595749
Gc7_98 0 n14 ns98 0 -9.46704884364e-05
Gc7_99 0 n14 ns99 0 0.000137424118057
Gc7_100 0 n14 ns100 0 -2.71491985409e-05
Gc7_101 0 n14 ns101 0 -0.000230063851563
Gc7_102 0 n14 ns102 0 -3.39590745056e-06
Gc7_103 0 n14 ns103 0 0.000702757308051
Gc7_104 0 n14 ns104 0 -6.26638663213e-06
Gd7_5 0 n14 ni5 0 0.000315138206101
Gd7_6 0 n14 ni6 0 0.000385794457697
Gd7_7 0 n14 ni7 0 -0.000318659757872
Gd7_8 0 n14 ni8 0 0.00155013910939
Gc8_53 0 n16 ns53 0 7.63371248733e-06
Gc8_54 0 n16 ns54 0 -1.03386931625e-05
Gc8_55 0 n16 ns55 0 1.70118546675e-05
Gc8_56 0 n16 ns56 0 -6.69174069358e-05
Gc8_57 0 n16 ns57 0 -0.00041133510426
Gc8_58 0 n16 ns58 0 -0.000698733322723
Gc8_59 0 n16 ns59 0 -4.05792279847e-05
Gc8_60 0 n16 ns60 0 -3.71465337128e-05
Gc8_61 0 n16 ns61 0 -1.23189660533e-06
Gc8_62 0 n16 ns62 0 -1.30982242137e-05
Gc8_63 0 n16 ns63 0 3.53427962331e-06
Gc8_64 0 n16 ns64 0 5.13641247963e-05
Gc8_65 0 n16 ns65 0 2.84462664286e-05
Gc8_66 0 n16 ns66 0 0.000592652286889
Gc8_67 0 n16 ns67 0 0.000968960244026
Gc8_68 0 n16 ns68 0 4.59426853158e-05
Gc8_69 0 n16 ns69 0 0.000686193579921
Gc8_70 0 n16 ns70 0 -0.000371918092218
Gc8_71 0 n16 ns71 0 -0.00163531086767
Gc8_72 0 n16 ns72 0 -5.66934403148e-05
Gc8_73 0 n16 ns73 0 7.0540258634e-05
Gc8_74 0 n16 ns74 0 -2.40540694015e-06
Gc8_75 0 n16 ns75 0 -7.11082409399e-05
Gc8_76 0 n16 ns76 0 2.45823275745e-06
Gc8_77 0 n16 ns77 0 0.000222025945238
Gc8_78 0 n16 ns78 0 1.33820096125e-05
Gc8_79 0 n16 ns79 0 0.000464549364354
Gc8_80 0 n16 ns80 0 0.000729546096376
Gc8_81 0 n16 ns81 0 6.21067673478e-05
Gc8_82 0 n16 ns82 0 0.000479841897053
Gc8_83 0 n16 ns83 0 -0.00144898749631
Gc8_84 0 n16 ns84 0 -0.00348468595749
Gc8_85 0 n16 ns85 0 -9.46704884364e-05
Gc8_86 0 n16 ns86 0 0.000137424118057
Gc8_87 0 n16 ns87 0 -2.71491985409e-05
Gc8_88 0 n16 ns88 0 -0.000230063851563
Gc8_89 0 n16 ns89 0 -3.39590745055e-06
Gc8_90 0 n16 ns90 0 0.00070275730805
Gc8_91 0 n16 ns91 0 -6.26638663231e-06
Gc8_92 0 n16 ns92 0 0.00038436134727
Gc8_93 0 n16 ns93 0 0.000540080325188
Gc8_94 0 n16 ns94 0 9.40293709717e-05
Gc8_95 0 n16 ns95 0 0.000361879809206
Gc8_96 0 n16 ns96 0 -0.00145456747916
Gc8_97 0 n16 ns97 0 -0.00376077843219
Gc8_98 0 n16 ns98 0 -0.00013088120037
Gc8_99 0 n16 ns99 0 0.000136341125514
Gc8_100 0 n16 ns100 0 7.60751465728e-05
Gc8_101 0 n16 ns101 0 0.000133935567018
Gc8_102 0 n16 ns102 0 3.63488558216e-05
Gc8_103 0 n16 ns103 0 -0.00149986958399
Gc8_104 0 n16 ns104 0 -0.000710410648662
Gd8_5 0 n16 ni5 0 0.000365460831508
Gd8_6 0 n16 ni6 0 0.000138868871671
Gd8_7 0 n16 ni7 0 0.00155013910939
Gd8_8 0 n16 ni8 0 0.00154102322751
.ends m4lines_port_fws
