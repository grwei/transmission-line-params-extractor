* BEGIN ANSOFT HEADER
* node 1    1:trace_p_0_T1_A
* node 2    1:trace_n_0_T1_A
* node 3    1:trace_n_1_T1_A
* node 4    1:trace_p_1_T1_A
* node 5    Ground_A
* node 6    1:trace_p_0_T1_B
* node 7    1:trace_n_0_T1_B
* node 8    1:trace_n_1_T1_B
* node 9    1:trace_p_1_T1_B
* node 10   Ground_B
*  Project: 4lines_veryHighFreq
*   Design: 2-diff-pairs
*   Length: 5
*   Format: HSPICE
*  Creator: Ansoft HFSS
*     Date: Sat Jun 06 18:38:17 2020
* END ANSOFT HEADER

.subckt ckt_m4lines_veryHighFreq_W 1 2 3 4 inref 5 6 7 8 outref length=2.54M

.model m4lines_veryHighFreq_W_1 W MODELTYPE=table N=4
+ RMODEL=r_m4lines_veryHighFreq_W_1 LMODEL=l_m4lines_veryHighFreq_W_1
+ GMODEL=g_m4lines_veryHighFreq_W_1 CMODEL=c_m4lines_veryHighFreq_W_1

* Example usage:
W1 1 2 3 4 inref 5 6 7 8 outref N=4 L=length TABLEMODEL=m4lines_veryHighFreq_W_1

.model r_m4lines_veryHighFreq_W_1 sp N=4 SPACING=nonuniform VALTYPE=real
+ INTERPOLATION=spline
+ DATA = 600
+ 0           
+        6.261736242051261
+       0.6684715379461887
+        6.377864916833254
+       0.2826728878941096
+       0.8559903459373164
+        6.374345933058062
+       0.1201295641379421
+       0.2811319884149726
+       0.6661056209785412
+         6.27437506597599
+ 6e+08       
+        17.16602021463065
+        1.581718391472655
+        17.51036311303858
+       0.6614412203087239
+        2.254836236598286
+         17.4912630450617
+       0.2420325169879826
+        0.656980418127239
+        1.581752083724183
+        17.22949207405247
+ 1.1e+09     
+        23.59351460335346
+        1.970831241751713
+         24.1048480387836
+       0.8006082533660617
+        3.026161731564372
+        24.07819871982417
+       0.2088873961887264
+       0.7955773917357565
+        1.973891104446969
+        23.69328765132619
+ 1.6e+09     
+         29.3175635182098
+        2.330345152429206
+        30.04640119176534
+       0.7945607007167228
+        3.614970840830058
+        30.01294884621569
+      -0.1444487808025694
+       0.7930774588734827
+        2.334779943959239
+         29.4570691053138
+ 2.1e+09     
+        34.38590372235392
+        2.867247744533854
+        35.18649325133151
+       0.9004364561810362
+        4.084624582322306
+        35.15336384534071
+      -0.3546848150431027
+       0.8993795543263321
+        2.871994828126375
+        34.54833362784322
+ 2.6e+09     
+         38.5423097625984
+        3.251967345894116
+        39.33381652721985
+          1.0246614425912
+        4.381617080110924
+        39.30567974687667
+      -0.4069411399700977
+        1.021628527039997
+        3.256197181878748
+        38.71549024004252
+ 3.1e+09     
+        41.98329072612757
+        3.496943600316263
+        42.75196559479232
+        1.167668088314755
+        4.623337350489276
+        42.73123299909383
+      -0.3051732854717014
+          1.1611095431772
+        3.500334573822903
+        42.16051774632864
+ 3.6e+09     
+        44.98480461622582
+        3.705083061670372
+        45.75991763249516
+        1.357871665938491
+        4.970202610793359
+        45.74773837577082
+     -0.06902803846415684
+        1.346839684456547
+        3.707723854678363
+        45.16297178006421
+ 4.1e+09     
+        47.77060417996347
+        3.970678248928344
+        48.60319766503232
+        1.622968582583021
+        5.555703602264881
+        48.60014948317339
+       0.2729093325795016
+        1.606945869805822
+         3.97290837802092
+         47.9486190052937
+ 4.6e+09     
+        50.48805316123251
+        4.347922586067769
+        51.42821882890364
+        1.972006533392416
+        6.410117421277009
+        51.43463906274915
+       0.6864648008413685
+        1.950817321075046
+        4.350158459043644
+        50.66585302493288
+ 5.1e+09     
+        53.21761305360312
+        4.844094100232534
+        54.28757388820721
+         2.38405084195086
+        7.401184135373949
+        54.30366893524681
+        1.133107514525441
+        2.357819184881632
+        4.846623526176458
+        53.39556241423573
+ 5.6e+09     
+        55.98953585659228
+        5.426262984315174
+         57.1704947232607
+         2.81879786545518
+        8.305981399047335
+        57.19633413554457
+        1.573481978323348
+        2.787934431801826
+         5.42900240150755
+        56.16802989539996
+ 6.1e+09     
+        58.80014737472479
+        6.037086363955919
+        60.05083024360616
+        3.246770311825928
+        9.003489498970186
+        60.08629777308323
+        1.974063246222053
+        3.211979891053165
+        6.039352298894379
+        58.97934545680759
+ 6.6e+09     
+        61.62513424930499
+        6.610723592592122
+        62.91223222025369
+        3.661737390807022
+        9.549503096523232
+         62.9570080518913
+        2.311753600704219
+        3.624036255328011
+        6.611170979304896
+        61.80482282238584
+ 7.1e+09     
+        64.43105227460738
+         7.08971862949311
+        65.74197940329421
+        4.066440350057811
+        10.07068536310605
+        65.79564245178429
+        2.575697142606129
+        4.027160466984707
+        7.086691479540798
+        64.61068587942748
+ 7.6e+09     
+        67.18805748996546
+        7.452027265532099
+        68.52585611428609
+         4.46152081681047
+        10.65866198686495
+        68.58815679728761
+        2.771720542477905
+        4.422239521330206
+        7.444458381772193
+        67.36700211332473
+ 8.1e+09     
+        69.88294395838609
+        7.743816671447835
+        71.25658467517061
+         4.85167755667857
+        11.34689455225178
+        71.32777475270993
+        2.932002846082346
+        4.813917344987765
+        7.732269519070353
+        70.06078327861394
+ 8.6e+09     
+        72.52639027340503
+        8.095806706621955
+        73.94343083153043
+        5.263061523029681
+         12.1306976368427
+        74.02432254353928
+        3.129043772044632
+        5.227489187487424
+        8.082534058857787
+        72.70293492292826
+ 9.1e+09     
+        75.14809742255692
+         8.70076393759506
+        76.61051427987179
+        5.765637728069409
+        12.99140484641196
+        76.70199898037887
+        3.493177375720148
+        5.730512646355473
+         8.68785939020713
+        75.32280026808829
+ 9.6e+09     
+        77.78131902974312
+        9.756234062009833
+        79.28354254967662
+        6.498100801299851
+        13.91400026527981
+        79.38579007492103
+        4.234635369891269
+        6.457125057469984
+        9.742646776459974
+        77.95233103592048
+ 1.01e+10    
+         78.5367572374255
+         10.1018393723646
+        79.94979593039989
+        6.762142142986897
+        14.06906916462574
+        80.06266861342931
+         5.01288153779625
+        6.702002593205487
+        10.08449902887477
+        78.71962788984995
+ 1.06e+10    
+        71.81949044042904
+        5.505293058615679
+        72.65479941492411
+        3.507209198105161
+        10.91875361723849
+        72.78218172472999
+        3.512991682848697
+         3.41757387810189
+        5.492791905845868
+        72.08953591804642
+ 1.11e+10    
+        65.38391369498106
+       0.9617392035804087
+        65.61053493448925
+       0.1465266363375564
+        7.752965235456211
+        65.75383596216955
+        1.980119387781448
+      0.02680638723292628
+        0.954214455404033
+        65.74015922640436
+ 1.16e+10    
+        59.25737891439243
+       -3.509041623975814
+        58.84866085775177
+       -3.318984337710113
+        4.581619789486691
+        59.00915110883384
+       0.4163307616431164
+       -3.469197113772524
+       -3.511592150188038
+        59.69745533151519
+ 1.21e+10    
+        53.46291040672862
+       -7.888823432959039
+        52.39632872449253
+       -6.889398467024413
+        1.413800902902104
+        52.57512818223208
+       -1.176738476020045
+       -7.070285949378788
+       -7.886517723226063
+        53.98328912257312
+ 1.26e+10    
+        48.01947716179243
+       -12.16095073162888
+        46.27639963621113
+       -10.56587184545323
+       -1.742268695854571
+        46.47446956313158
+       -2.797915963998386
+       -10.77734077351139
+       -12.15399864007415
+        48.61569893068838
+ 1.31e+10    
+        42.94227590004397
+       -16.31034135757736
+        40.50769212954282
+        -14.3507344734171
+       -4.879253067940114
+        40.72583011385909
+       -4.446527020053935
+       -14.59235896096365
+       -16.29902104367387
+        43.60916622546332
+ 1.36e+10    
+        38.24301722075879
+       -20.32347870831839
+        35.10524971706981
+       -18.24759190036323
+       -7.990727924378829
+        35.34408742182177
+       -6.122430850862138
+        -18.5185477579784
+       -20.30811387271571
+        38.97488388037247
+ 1.41e+10    
+        33.93020871797519
+       -24.18839565481673
+        30.08061807990692
+       -22.26143805407679
+       -11.07120613657965
+        30.34062112233308
+       -7.826059245702012
+       -22.56042692997534
+       -24.16933376169507
+         34.7210189624861
+ 1.46e+10    
+        30.00943023795504
+       -27.89465222334274
+         25.4421236271043
+        -26.3987815693316
+       -14.11616546312354
+        25.72359301169021
+       -9.558458421810386
+       -26.72394280797108
+       -27.87224370239683
+        30.85296682957462
+ 1.51e+10    
+        26.48359755355848
+       -31.43330895171591
+        21.19514675107559
+       -30.66778819147441
+       -17.12207996665412
+        21.49822128085859
+       -11.32133477858518
+       -31.01659583391355
+       -31.40788721659884
+         27.3735940035353
+ 1.56e+10    
+        23.35321165103215
+       -34.79689766700012
+        17.34238455455478
+       -35.07844215002326
+       -20.08645653249753
+        17.66704365866432
+       -13.11710542263931
+       -35.44758393968327
+       -34.76875965969967
+        24.28346786400936
+ 1.61e+10    
+         20.6165915823477
+       -37.97939129813589
+         13.8840990821818
+       -39.64272977649115
+        -23.0078778756915
+        14.23016550790252
+       -14.94895444673573
+       -40.02796436550337
+       -37.94877816189206
+        21.58107168932681
+ 1.66e+10    
+        18.27008945043439
+       -40.97617422590491
+        10.81834815724948
+       -44.37484908118812
+       -25.88605343269214
+        11.18548998377568
+       -16.82089608124497
+       -44.77083682760171
+       -40.94325161504125
+        19.26300397644497
+ 1.71e+10    
+        16.30828658183936
+       -43.78401458706494
+        8.141196801806007
+       -49.29144950317026
+       -28.72187957820556
+        8.528928231079144
+       -18.73784598614716
+       -49.69155127523109
+       -43.74885203219624
+        17.32416130611014
+ 1.76e+10    
+        14.72417031762041
+       -46.40103988544394
+        5.846907922660563
+       -54.41190659862431
+       -31.51751068243735
+        6.254588291988163
+        -20.7057021112586
+       -54.80794382075852
+       -46.36358853884498
+        15.75790429197638
+ 1.81e+10    
+        13.50929113416481
+       -48.82671721884049
+        3.928111492302825
+       -59.75863701799094
+       -34.27644262080035
+        4.354941923996169
+        -22.7314367168035
+       -60.14060475972367
+        -48.7867852017672
+        14.55620636887001
+ 1.86e+10    
+        12.65390000647179
+       -51.06183940066629
+        2.375951869626427
+       -65.35745970674047
+       -37.00361045267564
+         2.82096892675851
+       -24.82320130298844
+       -65.71318288151178
+       -51.01906385332371
+        13.70978534543744
+ 1.91e+10    
+        12.14706606378187
+       -53.10851823150642
+        1.180213208665389
+       -71.23800979217634
+       -39.70550208038816
+        1.642278854973449
+       -26.99044632912469
+       -71.55273044398595
+       -53.06233302279882
+        13.20821777823085
+ 1.96e+10    
+        11.97677467959231
+       -54.97018614508582
+       0.3294231304594604
+       -77.43421198808169
+       -42.39028974638381
+       0.8072102002781829
+       -29.24405767812057
+       -77.69009314816789
+       -54.91978402560365
+        13.04003633255399
+ 2.01e+10    
+        12.13000620724028
+       -56.65160739561268
+          185.87993952924
+       -83.98482040341682
+       -45.06798117922371
+       0.3029072699044058
+       -31.59651179176196
+       -84.16034905048434
+       -56.59589517023863
+        13.19281039540314
+ 2.06e+10    
+        12.59279564734924
+       -58.15889983686294
+        196.9127933108171
+        -90.9340311229347
+       -47.75059197335608
+       0.1153751363756852
+       -34.06205119044962
+       -91.00329935857148
+       -58.09644488835549
+        13.65321032361838
+ 2.11e+10    
+        13.35027365393199
+       -59.49956811999868
+        208.2159229139332
+       -98.33217243605701
+       -50.45234026649615
+       0.2295132149699635
+       -36.65688157560007
+       -98.26401211931029
+       -59.42853433410501
+         14.4070558772221
+ 2.16e+10    
+        14.38668950862774
+       -60.68254873010074
+       0.1063527756321134
+       -106.2364745017162
+       -53.18986376886519
+       0.6291283336998372
+       -39.39939071318152
+       -105.9934163968788
+       -60.60061956322792
+        15.43934965396196
+ 2.21e+10    
+        15.68541710114248
+       -61.71826657704358
+       0.7688569366335898
+       -114.7119145855321
+       -55.98245742465422
+        1.296928684561782
+       -42.31038752850671
+       -114.2489388630658
+       -61.62255268987195
+        16.73429677534487
+ 2.26e+10    
+        17.22894567220824
+       -62.61870167772429
+        1.684288707853142
+       -123.8321243242683
+        -58.8523270112675
+        2.214500950523559
+       -45.41335688508578
+        -123.095165612563
+       -62.50563027529923
+        18.27531277874338
+ 2.31e+10    
+        18.99885829042925
+       -63.39746254905233
+        2.833593206634184
+        -133.680329528023
+       -61.82484917453571
+        3.362274407444884
+       -48.73472073560391
+       -132.6044977513195
+       -63.26264539909502
+        20.04502279509501
+ 2.36e+10    
+        20.97580302327205
+       -64.06985987659731
+        4.196613893973842
+       -144.3502674820158
+       -64.92882080073635
+        4.719478241094778
+       -52.30408878037522
+       -142.8577473860929
+       -63.90793706571735
+        22.02525685260689
+ 2.41e+10    
+        23.13946493717864
+       -64.65296924561035
+        5.752071607188915
+       -155.9469866033111
+       -68.19666885261876
+        6.264102191505442
+       -56.15447006444622
+       -153.9445874773111
+       -64.45742631878397
+        24.19704885722707
+ 2.46e+10    
+        25.46855202411049
+       -65.16566436171716
+        7.477563787582236
+       -168.5873714269808
+       -71.66457384112081
+        7.972876644811352
+       -60.32239910057044
+       -165.9637195555402
+       -64.92862197960699
+        26.54065090311035
+ 2.51e+10    
+        27.94081575923705
+       -65.62859103558517
+        9.349607283180028
+       -182.4001419808362
+       -75.37243315489327
+        9.821297454758334
+       -64.84790332460844
+       -179.0225506220032
+       -65.34056932552396
+        29.03558067288922
+ 2.56e+10    
+        30.53313843522079
+       -66.06403558793242
+         11.3437601465594
+       -197.5249365818548
+       -79.36355071565731
+        11.78373447452864
+       -69.77419918898956
+       -193.2360655733095
+       -65.71370098661643
+        31.66072861377392
+ 2.61e+10    
+        33.22173624124717
+       -66.49561709333427
+        13.43487519946153
+       -214.1098827581652
+       -83.68388202574494
+          13.833682809897
+       -75.14694716145763
+       -208.7244330966001
+       -66.06952923814157
+        34.39456433887923
+ 2.66e+10    
+        35.98255109600588
+       -66.94769850329179
+        15.59756243643701
+       -232.3067712415108
+        -88.3805831115414
+        15.94424427102128
+        -81.0128158414455
+        -225.608679308238
+       -66.43009088716977
+        37.21549943008087
+ 2.71e+10    
+        38.79193724281018
+       -67.44436486072171
+        17.80697000063984
+        -252.262553684319
+       -93.49950335795612
+        18.08896534291166
+       -87.41699757048015
+       -244.0034956503695
+       -66.81701857703598
+        40.10248744058362
+ 2.76e+10    
+        41.62779118882161
+       -68.00775692028502
+        20.04003465211813
+       -274.1053819213051
+       -99.08112522602821
+        20.24320779449999
+       -94.39918173829631
+       -264.0059188536443
+       -67.25006552616838
+        43.03597140353295
+ 2.81e+10    
+        44.47132287442338
+       -68.65547992726255
+        22.27739906388323
+         -297.92283522044
+       -105.1542996458405
+        22.38628528561083
+       -101.9873386770571
+         -285.67826434126
+       -67.74485846305774
+        45.99932204352336
+ 2.86e+10    
+        47.30971110538661
+       -69.39674594610408
+        24.50623401494132
+       -323.7294823595217
+       -111.7269921564521
+        24.50465111998523
+       -110.1885339872649
+        -309.023406722577
+       -68.30960854221917
+        48.98093826527509
+ 2.91e+10    
+        50.13990039681069
+       -70.22689236364822
+        26.72421305262328
+       -351.4208339951635
+       -118.7732300710319
+        26.59643729342522
+       -118.9759681957253
+       -333.9504950476411
+        -68.9405016846211
+        51.97718728617306
+ 2.96e+10    
+        52.97372530919011
+       -71.12002545064497
+        28.94481565942256
+       -380.7117240465035
+       -126.2156980603494
+        28.67756058362178
+       -128.2716916323732
+       -360.2298665999078
+       -69.61557481014657
+        54.99631024177638
+ 3.01e+10    
+        55.84430026262169
+       -72.01989458284467
+        31.20389968779707
+       -411.0603288198454
+       -133.9042554243689
+        30.78932207532312
+       -137.9252643427145
+       -387.4379262714848
+       -70.28715631912389
+         58.0632530885255
+ 3.06e+10    
+        58.81306372942813
+       -72.82988165283207
+         33.5669741961758
+       -441.5858564956307
+       -141.5924231086429
+        33.00679010660835
+        -147.690393554419
+       -414.8969292567256
+       -70.87353219086062
+        61.22502592770329
+ 3.11e+10    
+        61.97591467643704
+       -73.40432895474066
+        36.13572687524996
+       -470.9995317617035
+       -148.9169161851054
+        35.44615677857605
+       -157.2045890580376
+       -441.6216257044658
+       -71.25149661427969
+        64.55558113168537
+ 3.16e+10    
+        65.46559980956685
+       -73.54522070745188
+        39.05116511899939
+       -497.5837454424791
+       -155.3893517697427
+        38.26777466668908
+       -165.9809057139863
+       -466.2941980292601
+       -71.25280137983403
+        68.15835901896884
+ 3.21e+10    
+        69.44640504101575
+       -73.00977742394932
+         42.4896202217156
+       -519.2667360944904
+       -160.4128295903652
+         41.6702762315992
+       -173.4243892123099
+       -487.2977998703316
+       -70.66877707081464
+        72.16384023124213
+ 3.26e+10    
+        74.09739217371224
+       -71.53426646736645
+        46.64777814766654
+       -533.8361801757992
+       -163.3357825407194
+        45.87131794268421
+       -178.8855483324719
+       -502.8402201443049
+       -69.26750789962554
+        76.71928974739379
+ 3.31e+10    
+        79.58329468029396
+       -68.87534100339182
+         51.7151032689342
+       -539.2981340782165
+       -163.5470030222919
+        51.07367765173038
+       -181.7547463995672
+       -511.1829130114555
+       -66.82547225953677
+        81.96925828020672
+ 3.36e+10    
+        86.01808269495901
+       -64.86199481481626
+        57.83710343452189
+       -534.3152614513253
+        -160.597609712788
+        57.42214237607202
+       -181.5833840252964
+       -510.9512668390543
+       -63.16981886196795
+        88.02883432818507
+ 3.41e+10    
+        93.43268644753371
+       -59.44208357096726
+        65.07924468693105
+        -518.581783920844
+       -154.3145941307888
+        64.96423238991241
+       -178.1967520842151
+       -501.4497622729743
+       -58.22017932232271
+        94.95622236018606
+ 3.46e+10    
+        101.7604275522317
+       -52.70422760261748
+        73.40482987216058
+       -492.9732853843835
+       -144.8614469882316
+        73.63068279193152
+       -171.7543401084627
+        -482.871502958403
+       -52.01475567386238
+        102.7342365792634
+ 3.51e+10    
+        110.8477555455697
+       -44.86390913508254
+        82.67681846955681
+       -459.3880433137018
+       -132.7166752083277
+        83.24538425883514
+       -162.7285809638132
+       -456.3100669316855
+         -44.708977470522
+        111.2687197608402
+ 3.56e+10    
+        120.4864429983883
+       -36.21850705503802
+        92.68384364397713
+       -420.3374179755984
+       -118.5760140970217
+        93.56150801499149
+       -151.8077720591369
+       -423.5568775529107
+       -36.54600792191101
+         120.405394313818
+ 3.61e+10    
+        130.4541694690646
+       -27.08930282435965
+         103.180434541439
+       -378.4502061542368
+        -103.216579098659
+        104.3093349938901
+       -139.7611498541884
+       -386.7575632841152
+       -27.81028248204926
+        129.9588874450629
+ 3.66e+10    
+        140.5493159401227
+        -17.7706757517936
+        113.9271815001681
+       -336.0615250770351
+       -87.37048330120706
+        115.2390209253915
+        -127.313331924996
+       -348.0489163267643
+       -18.78053637085679
+        139.7435609850303
+ 3.71e+10    
+        150.6118038291974
+       -8.498689992461252
+        124.7198438779208
+       -294.9783446519555
+       -71.64028693789184
+        126.1477754072693
+       -115.0602933185628
+       -309.2807587082574
+       -9.695325555828425
+        149.5972612609946
+ 3.76e+10    
+        160.5294226595003
+       0.5594578690733361
+        135.4034561445048
+       -256.4209013098197
+       -56.46418329002626
+         136.889747454372
+       -103.4347460588193
+       -271.8688626794379
+      -0.7359624655790924
+        159.3940428859228
+ 3.81e+10    
+        170.2338486795326
+        9.300714885851008
+        145.8735402507723
+       -221.0844088796938
+       -42.12053475249935
+        147.3729312249228
+       -92.71061586457867
+       -236.7683031358195
+        7.975351395652076
+        169.0467217294921
+ 3.86e+10    
+        179.6916018631826
+        17.67360055136008
+        156.0692810560163
+       -189.2562534568121
+       -28.75477389369038
+        157.5491692913999
+       -83.02974786180512
+       -204.5266138299567
+        16.36778178233607
+        178.5026498135253
+ 3.91e+10    
+        188.8939753592287
+        25.66370926470869
+        165.9633968544713
+       -160.9407739400379
+       -16.41379404160846
+        167.4022358897396
+       -74.43606366235028
+       -175.3732072159298
+         24.4100663314555
+        187.7363632958379
+ 3.96e+10    
+        197.8481856269559
+        33.28071520949081
+         175.551956293874
+       -135.9661154284084
+       -5.078425616624946
+        176.9369677733108
+       -66.90782528207924
+          -149.3132753597
+        32.09854216491453
+        196.7417800617808
+ 4.01e+10    
+        206.5705694826955
+        40.54823454108766
+        184.8457962530522
+       -114.0647047783223
+        5.310281426545818
+        186.1706760240385
+       -60.38375127146068
+       -126.2089254834884
+        39.44699950162135
+        205.5254112232711
+ 4.06e+10    
+        215.0818238075878
+        47.49664203514389
+        193.8640453441339
+       -94.92846772520524
+        14.83185811743046
+        195.1269916903329
+       -54.78209921540664
+       -105.8414694777888
+        46.47899580309978
+        214.1011157979951
+ 4.11e+10    
+        223.4039255205682
+        54.15836786025451
+        202.6296239417126
+       -78.24377346525232
+        23.57347719745532
+        203.8317893093809
+       -50.01353013050938
+       -87.95528118426535
+        53.22250078273974
+        222.4863805404419
+ 4.16e+10    
+          231.55829059345
+        60.56505039319814
+        211.1663364468265
+       -63.71171361376924
+        31.62186730855424
+        212.3106844463219
+       -45.98915118254769
+       -72.28646172580571
+        59.70642878884224
+        230.6998654460283
+ 4.21e+10    
+        239.5647806681284
+        66.74597432034707
+        219.4971320616883
+       -51.05852424907368
+         39.0586847384247
+        220.5876325320607
+       -42.62512289095018
+       -58.58018394572455
+        65.95856103527943
+        238.7598981493528
+ 4.26e+10    
+        247.4412555957391
+        72.72734592119173
+        227.6431675453125
+       -40.03977671014614
+        45.95819585301353
+         228.684252263712
+        -39.8449699279258
+       -46.60017743905095
+        72.00442409410171
+        246.6836312706699
+ 4.31e+10    
+         255.203457966925
+        78.53208341904008
+        235.6233905733483
+       -30.44086364475461
+        52.38641918549965
+        236.6195997600273
+       -37.58044090461701
+       -36.13306268837218
+        77.86679036520837
+        254.4866374833242
+ 4.36e+10    
+        262.8650864355627
+        84.17990436286014
+        243.4544430953075
+       -22.07544448038099
+         58.4011363142724
+        244.4102063903833
+       -35.77150417544582
+       -26.98949023080851
+        83.56556151227359
+        262.1827787010623
+ 4.41e+10    
+        270.4379662911921
+        89.68756923639609
+        251.1507490227291
+       -14.78289668898685
+        64.05238121722765
+         252.070258382656
+       -34.36586749219578
+       -19.00342022631781
+        89.11787289789672
+        269.7842370203302
+ 4.46e+10    
+        277.9322612022393
+        95.06919416405212
+        258.7246983530916
+        -8.42540164418552
+        69.38316107375256
+        259.6118420598079
+       -33.31826700397234
+       -12.03041426887491
+        94.53831392047647
+         277.301633563474
+ 4.51e+10    
+        285.3566933650882
+        100.3365812183812
+        266.1868730358521
+       -2.885023372620313
+        74.43025876282502
+         267.045209179959
+       -32.58967445357111
+       -5.945485761108399
+        99.83919876707952
+        284.7441885661156
+ 4.56e+10    
+        292.7187540926049
+        105.4995376581192
+        273.5462820314597
+        1.939030641585361
+        79.22503086815193
+        274.3790366320143
+       -32.14650826630707
+      -0.6408363257178245
+        105.0308485690777
+        292.1198944416613
+ 4.61e+10    
+        300.0248959689421
+        110.5661695752097
+        280.8105873090179
+        6.132879653902549
+        83.79415518606196
+        281.6206670919258
+       -31.95989429747466
+        3.976336391472912
+        110.1218630441807
+        299.4356855691296
+ 4.66e+10    
+        307.2807030974399
+        115.5431439117948
+        287.9863114702306
+        9.770143324201371
+        88.16030633317318
+        288.7763247351283
+       -32.00499754711021
+        7.985863626454465
+        115.1193704309383
+        306.6975961720354
+ 4.71e+10    
+        314.4910390329316
+        120.4359176828433
+        295.0790231138312
+        12.91382407993013
+        92.34275256901228
+        295.8513044451718
+       -32.26043172842906
+         11.4564217138021
+        120.0292510161733
+        313.9109023367683
+ 4.76e+10    
+         321.660173619336
+        125.2489358747909
+        302.0934992043061
+        15.61792001296201
+        96.35787508776495
+         302.850135365008
+       -32.70774547825012
+        14.44713013782946
+         124.856333344981
+        321.0802469981805
+ 4.81e+10    
+         328.791890722249
+        129.9858007748436
+        309.0338654442031
+        17.92879723318886
+        100.2196152598605
+        309.7767208337378
+       -33.33097979422214
+        17.00893961637078
+        129.6045642806013
+        328.2097482843844
+ 4.86e+10    
+        335.8895791126185
+        134.6494159726682
+        315.9037165062475
+        19.88635229056055
+        103.9398571696489
+         316.634457260076
+       -34.11628942856946
+        19.18582732233951
+        134.2771551182249
+        335.3030924294728
+ 4.91e+10    
+        342.9563087489482
+         139.242108319937
+        322.7062183251961
+        21.52499408491943
+        107.5287533150284
+        323.4263345747871
+       -35.05162045047321
+        21.01582001222524
+        138.8767063677349
+        342.3636128219029
+ 4.96e+10    
+        349.9948945531249
+        143.7657309417017
+        329.4441946906968
+        22.87447208817376
+        110.9950010903675
+        330.1550207847834
+       -36.12643642211436
+        22.53186647775511
+        143.4053138749204
+        349.3943568545293
+ 5.01e+10    
+        357.0079495576849
+         148.221750089914
+        336.1202002671346
+        23.96057457454196
+        114.3460770753827
+        336.8229329298618
+       -37.33148623976029
+        23.76257974184323
+        147.8646588146322
+        356.3981421895592
+ 5.06e+10    
+        363.9979290693735
+        152.6113182965957
+        342.7365819736018
+        24.80571736995094
+        117.5884353777892
+        343.4322964762207
+       -38.65860744709943
+        24.73286762725817
+        152.2560838588709
+        363.3776039268925
+ 5.11e+10    
+        370.9671672653989
+        156.9353359475887
+        349.2955304369559
+        25.42944063329476
+        120.7276754893217
+        349.9851949142225
+       -40.10055961842247
+        25.46446822171741
+        156.5806575599474
+        370.3352340067063
+ 5.16e+10    
+        377.9179074289151
+        161.1945030889777
+         355.799123002775
+        25.84882848556534
+        123.7686843460804
+        356.4836110745075
+       -41.65088316960263
+        25.97640463038497
+        160.8392287210099
+        377.2734140120143
+ 5.21e+10    
+        384.8523268454809
+        165.3893630044335
+        362.2493595921707
+        26.07886395043617
+        126.7157565990155
+        362.9294614544463
+       -43.30377963343641
+         26.2853713957551
+        165.0324722813955
+         384.194442379518
+ 5.26e+10    
+        391.7725572192557
+         169.520338856058
+        368.6481924911795
+        26.13272963895323
+        129.5726964822995
+        369.3246246428367
+       -45.05401005346062
+        26.40606314326869
+        169.1609280155541
+        391.1005568820171
+ 5.31e+10    
+         398.680701331179
+        173.5877644798099
+        374.9975510031341
+        26.02206290155951
+        132.3429041394945
+        375.6709647606826
+       -46.89680866798313
+        26.35145440586242
+        173.2250331487649
+        397.9939531175099
+ 5.36e+10    
+        405.5788465423827
+        177.5919102451595
+        381.2993617472256
+        25.75717272079707
+        135.0294488134438
+        381.9703506913331
+       -48.82780951391911
+         26.1330381891347
+        177.2251498212452
+        404.8767996277065
+ 5.41e+10    
+        412.4690756504905
+        181.5330047459387
+        387.5555652654291
+        25.34722441310399
+          137.63513091876
+        388.2246717473258
+       -50.84298395640807
+        25.76102964866663
+        181.1615881856585
+        411.7512501718689
+ 5.46e+10    
+        419.3534755199538
+        185.4112529594154
+         393.768129495768
+        24.80039720067136
+        140.1625346926469
+        394.4358503164407
+       -52.93858747594125
+          25.244540239274
+        185.0346257987642
+         418.619453601048
+ 5.51e+10    
+        426.2341438425766
+        189.2268514116797
+        399.9390605797573
+        24.12401887668249
+        142.6140728500715
+        400.6058519478086
+       -55.11111431089682
+        24.59172684299342
+        188.8445238637566
+         425.483561705838
+ 5.56e+10    
+        433.1131943247856
+        192.9800007974125
+        406.0704114033084
+        23.32468109386938
+        144.9920244340182
+        406.7366932563436
+       -57.35725878214239
+        23.80991966428893
+        192.5915407898493
+        432.3457353540991
+ 5.61e+10    
+        439.9927605505268
+         196.670916430482
+        412.1642882024998
+        22.40833822773667
+        147.2985668703547
+         412.830447973192
+       -59.67388231270904
+         22.9057320789958
+        196.2759434640822
+        439.2081491841967
+ 5.66e+10    
+        446.8749987297051
+        200.2998368435425
+        418.2228555183363
+        21.38039228893351
+        149.5358030709199
+        418.8892514124086
+       -62.05798531171517
+        21.88515511979939
+        199.8980165667682
+        446.0729950790493
+ 5.71e+10    
+        453.7620895078632
+        203.8670308008972
+        424.2483397381104
+        20.24576596010649
+        151.7057842976459
+        424.9153035841824
+       -64.50668322722576
+        20.75363885783801
+        203.4580702098345
+        452.9424846094151
+ 5.76e+10    
+         460.656238986726
+        207.3728029518347
+        430.2430314258401
+          19.008965504213
+        153.8105293934994
+         430.910871149524
+       -67.01718617270825
+        19.51616258848645
+        206.9564461355951
+        459.8188506079053
+ 5.81e+10    
+        467.5596790793364
+         210.817498310825
+        436.2092866159697
+        17.67413501268757
+        155.8520408854386
+        436.8782883816643
+       -69.58678163616275
+        18.17729543172785
+        210.3935226746411
+        466.7043480093387
+ 5.86e+10    
+         474.474667308408
+        214.2015057293985
+        442.1495272131708
+        16.24510323834495
+        157.8323183955633
+        442.8199572748082
+       -72.21281984112485
+        16.74124871252742
+        213.7697186345505
+        473.6012540723984
+ 5.91e+10    
+        481.4034861356947
+        217.5252604918113
+        448.0662406261603
+          14.725424060179
+        159.7533697261519
+        448.7383469197913
+       -74.89270140639732
+        15.21192127703815
+        217.0854962610078
+        480.5118680812939
+ 5.96e+10    
+        488.3484419004589
+        220.7892461531844
+        453.9619787410682
+        13.11841147328226
+        161.6172199310643
+        454.6359922487337
+       -77.62386699480601
+        13.59293872726219
+        220.3413633956503
+        487.4385106098565
+ 6.01e+10    
+        495.3118634322971
+         223.993995717267
+        459.8393563268874
+        11.42716985858594
+        163.4259186431171
+        460.5154922396643
+       -80.40378868950467
+        11.88768741008583
+         223.537874935133
+        494.3835224205361
+ 6.06e+10    
+        502.2961003930472
+        227.1400922393457
+        465.7010489524005
+        9.654620177609194
+        165.1815458824134
+        466.3795076515794
+       -83.22996287439713
+         10.0993438742866
+        226.6756336802152
+        501.3492630583394
+ 6.11e+10    
+        509.3035213966597
+        230.2281689254666
+        471.5497904810263
+        7.803522641412599
+        166.8862165465026
+        472.2307583615245
+       -86.09990442416348
+        8.230900404041734
+         229.755290651744
+        508.3381091917977
+ 6.16e+10    
+        516.3365119466795
+        233.2589087900043
+         477.388370205099
+        5.876496325358969
+        168.5420837472961
+        478.0720203553976
+        -89.0111420359072
+         6.28518715126522
+        232.7775449396592
+        515.3524527463682
+ 6.21e+10    
+         523.397472228026
+        236.2330439262863
+        483.2196296702191
+        3.876036130428798
+        170.1513411404044
+        483.9061224251181
+       -91.96121455899002
+        4.264891312544524
+        235.7431431415426
+        522.3946988680624
+ 6.26e+10    
+         530.488814781286
+         239.151354434663
+        489.0464592332962
+        1.804527439111888
+        171.7162243778016
+        489.7359426123894
+       -94.94766819744221
+        2.172573737955464
+        238.6528784393814
+        529.4672637509456
+ 6.31e+10    
+        537.6129620879874
+        242.0146670492925
+        494.8717943958044
+       -0.335741235997169
+        173.2390117866095
+        495.5644044410391
+       -97.96805447044963
+      0.01068330103728954
+        241.5075893579229
+         536.572572356691
+ 6.36e+10    
+         544.772344086907
+        244.8238534971472
+        500.6986119443685
+        -2.54256735506906
+        174.7220243709597
+        501.3944729660564
+        -101.019928839264
+       -2.218430684059548
+        244.3081582399398
+        543.7130560510719
+ 6.41e+10    
+        551.9693956428787
+        247.5798286204356
+        506.5299259324574
+       -4.813824980973534
+        176.1676252230768
+        507.2291506719345
+       -104.1008499122172
+       -4.512507748487788
+        247.0555094720078
+        550.8911501792816
+ 6.46e+10    
+        559.2065539843296
+        250.2835482886449
+         512.368783524765
+       -7.147456745414493
+        177.5782184114382
+        513.0714732464604
+       -107.2083791518469
+       -6.869367046460525
+        249.7506074882405
+        558.1092915975449
+ 6.51e+10    
+         566.486256123471
+        252.9360071223896
+        518.2182607359376
+       -9.541466982250569
+        178.9562474102073
+        518.9245052497455
+       -110.3400810198334
+       -9.286899435596602
+         252.394454575561
+        565.3699161785584
+ 6.56e+10    
+        573.8109362732479
+        255.5382360504693
+        524.0814580754155
+       -11.99391588306393
+        180.3041931292648
+        524.7913357042734
+       -113.4935234966815
+       -11.76306069937587
+        254.9880885042827
+         572.675456303173
+ 6.61e+10    
+        581.1830232713339
+        258.0912997184915
+        529.9614961275904
+       -14.50291454740544
+        181.6245715867334
+        530.6750736189686
+       -116.6662789254278
+       -14.29586577027546
+        257.5325800012744
+        580.0283383520925
+ 6.66e+10    
+        588.6049380209963
+        260.5962937631075
+         535.861511075767
+       -17.06662081630187
+        182.9199312776552
+         536.578843468454
+       -119.8559251299485
+       -16.88338382806937
+        260.0290300823382
+        587.4309802072175
+ 6.71e+10    
+        596.0790909570773
+        263.0543419683572
+        541.7846501918103
+       -19.68323579273796
+        184.1928502654653
+        542.5057806396271
+       -123.0600467640001
+       -19.52373416736229
+        262.4785672613222
+        594.8857887719579
+ 6.76e+10    
+        603.6078795448656
+        265.4665933142431
+        547.7340673017685
+       -22.35100096250623
+        185.4459330414049
+         548.459026860992
+       -126.2762368561562
+       -22.21508273802249
+        264.8823446460608
+        602.3951575192798
+ 6.81e+10    
+        611.1936858179442
+        267.8342189321452
+         553.712918240121
+       -25.06819584006182
+        186.6818071745605
+        554.4417256250821
+       -129.5020985100189
+       -24.95563927531728
+        267.2415369353726
+        609.9614640734269
+ 6.86e+10    
+         618.838873960626
+        270.1584089739467
+        559.7243563101704
+       -27.83313607463055
+         187.903119782657
+        560.4570176195797
+       -132.7352467328548
+       -27.74365494514564
+        269.5573373279513
+        617.5870678331576
+ 6.91e+10    
+        626.5457879398547
+        272.4403694059688
+        565.7715277494054
+       -30.64417195626582
+        189.1125338509309
+        566.5080361705931
+       -135.9733103622021
+       -30.57742044197315
+        271.8309543506741
+        625.2743076389406
+ 6.96e+10    
+        634.3167491907789
+        274.6813187366781
+        571.8575672241539
+        -33.4996872712197
+         190.312724413965
+         572.597902714853
+       -139.2139340638672
+       -33.45526447876652
+        274.0636086185194
+          633.02549949272
+ 7.01e+10    
+        642.1540543597898
+        276.8824846837026
+        577.9855933499299
+       -36.39809846082984
+        191.5063746287027
+        578.7297223055119
+       -142.4547803813634
+       -36.37555262122341
+        276.2565295306876
+         640.842934330408
+ 7.06e+10    
+        650.0599731080554
+        279.0451007896805
+         584.158704253935
+       -39.33785404203245
+        192.6961717500903
+        584.9065791598582
+       -145.6935318116856
+       -39.33668641815637
+        278.4109519137636
+         648.728875853671
+ 7.11e+10    
+        658.0367459781068
+        281.1704029913799
+        590.3799731841492
+       -42.31743425515396
+        193.8848030283836
+        591.1315322593491
+       -148.9278928922816
+       -42.33710279080965
+        280.5281126154841
+        656.6855584216833
+ 7.16e+10    
+        666.0865823266294
+        283.2596261497816
+        596.6524441705099
+       -45.33535090506147
+        195.0749515438375
+        597.4076110043275
+       -152.1555922816827
+       -45.37527364343675
+        282.6092470584552
+        664.7151850077078
+ 7.21e+10    
+        674.2116583241982
+        285.3140005453764
+        602.9791277508541
+       -48.39014736858337
+        196.2692919893519
+         603.737810936016
+       -155.3743848170435
+       -48.44970566431832
+        284.6555857570961
+        672.8199252207438
+ 7.26e+10    
+        682.4141150256741
+        287.3347483459171
+        609.3629967615157
+       -51.48039874061078
+        197.4704864168183
+         610.125089524633
+       -158.5820535390586
+       -51.55894028910053
+        286.6683508047583
+         681.001913395362
+ 7.31e+10    
+        690.6960565098876
+        289.3230800484739
+        615.8069821997327
+       -54.60471209803452
+        198.6811799561813
+        616.5723620379736
+       -161.7764116703296
+       -54.70155379944028
+        288.6487523367766
+         689.263246751456
+ 7.36e+10    
+        699.0595480933689
+        291.2801909041879
+        622.3139691679264
+       -57.76172686020995
+        199.9039965188895
+        623.0824974878504
+       -164.9553045363118
+       -57.87615753707146
+        290.5979849727049
+        697.6059836251236
+ 7.41e+10    
+        707.5066146162483
+        293.2072573282708
+        628.8867929016629
+       -60.95011522627703
+        201.1415344957539
+        629.6583146644018
+       -168.1166114252095
+       -61.08139821063132
+        292.5172242430429
+         706.032141771322
+ 7.46e+10    
+        716.0392388028314
+        295.1054332986585
+        635.5282348819102
+       -64.16858267592906
+        202.3963624550833
+        636.3025782632212
+       -171.2582473744392
+       -64.31595827841363
+         294.407623006712
+        714.5436967402318
+ 7.51e+10    
+        724.6593596972837
+        296.9758467501582
+        642.2410190455425
+       -67.41586851573608
+        203.6710148561786
+        643.0179951050453
+       -174.3781648780367
+       -67.57855638946772
+        296.2703078599783
+        723.1425803280814
+ 7.56e+10    
+          733.36887117498
+        298.8195959667965
+        649.0278080932055
+       -70.69074645988182
+         204.967987777574
+        649.8072104593172
+       -177.4743555172123
+       -70.86794787065568
+        298.1063755451793
+        731.8306791025777
+ 7.61e+10    
+        742.1696205299885
+        300.6377459748774
+        655.8911998940239
+       -73.99202523215361
+        206.2897346747013
+        656.6728044699827
+        -180.544851499057
+       -74.18292524433357
+         299.916889360169
+        740.6098330043035
+ 7.66e+10    
+        751.0634071395981
+        302.4313249443336
+        662.8337240059302
+       -77.31854917992807
+        207.6386621694503
+        663.6172886907096
+        -183.587727112222
+       -77.52231876507815
+        301.7028755731574
+        749.4818340240098
+ 7.71e+10    
+        760.0519812057545
+        304.2013205985975
+        669.8578382955415
+       -80.66919888790267
+        209.0171258809025
+        670.6431027337148
+       -186.6011000881402
+       -80.88499696662187
+        303.4653198501144
+        758.4484249571547
+ 7.76e+10    
+        769.1370425738794
+        305.9486766384798
+        676.9659256784486
+       -84.04289178764171
+        210.4274262981493
+          677.75261102993
+       -189.5831328749334
+       -84.26986720730379
+        305.2051636923711
+        767.5112982344218
+ 7.81e+10    
+        778.3202396295532
+        307.6742891853176
+        684.1602909763501
+       -87.43858274891652
+        211.8718047118569
+        684.9480997146629
+       -192.5320338168777
+       -87.67587620691241
+        306.9233008944594
+        776.6720948307714
+ 7.86e+10    
+        787.6031682734481
+        309.3790032435317
+        691.4431578897213
+       -90.85526465117968
+         213.352439196348
+        692.2317736307208
+       -195.4460582461955
+       -91.10201056555627
+        308.6205740227379
+        785.9324032514101
+ 7.91e+10    
+        796.9873709735479
+        311.0636091905023
+        698.8166661007732
+       -94.29196892594607
+        214.8714406585282
+        699.6057534608652
+       -198.3235094834523
+       -94.54729726003566
+        310.2977709195667
+        795.2937585957108
+ 7.96e+10    
+        806.4743358971232
+        312.7288392949761
+        706.2828684983378
+       -97.74776606592997
+        216.4308489533919
+        707.0720729863526
+       -201.1627397509734
+       -98.01080410811241
+        311.9556212371699
+        804.7576416998892
+ 8.01e+10    
+        816.0654961200963
+        314.3753642684039
+        713.8437285356561
+       -101.2217660939457
+        218.0326290738148
+        714.6326764812318
+       -203.9621510009839
+       -101.4916401983438
+        313.5947930044898
+        814.3254783570857
+ 8.06e+10    
+        825.7622289157987
+        316.0037898555204
+        721.5011177215584
+       -104.7131189888231
+        219.6786674159846
+         722.289416237989
+       -206.7201956609156
+       -104.9889562772054
+        315.2158892324384
+         823.998638616612
+ 8.11e+10    
+        835.5658551223127
+        317.6146534632126
+        729.2568132439553
+       -108.2210150632978
+        221.3707681297454
+        730.0440502310382
+       -209.4353772988241
+        -108.501945091901
+        316.8194445592626
+        833.7784361621347
+ 8.16e+10    
+        845.4776385894568
+         319.208420838523
+        737.1124957375063
+       -111.7446852899868
+        223.1106495530051
+        737.8982399236231
+       -212.1062512138249
+       -112.0298416816933
+         318.405921943547
+        843.6661277681941
+ 8.21e+10    
+        855.4987857044655
+        320.7854827934967
+        745.0697471871889
+       -115.2834015722198
+        224.8999407402946
+        745.8535482158176
+       -214.7314249511886
+       -115.5719236155878
+        319.9757094050183
+        853.6629128359973
+ 8.26e+10    
+        865.6304449976143
+        322.3461519854947
+        753.1300489826757
+       -118.8364769564009
+        226.7401780866654
+        753.9114375375264
+        -217.309558751269
+       -119.1275111733878
+         321.529116822179
+         863.769933009392
+ 8.31e+10    
+        875.8737068275028
+        323.8906597562276
+        761.2947801112848
+       -122.4032657833474
+        228.6328020489619
+        762.0732680904874
+       -219.8393659313178
+       -122.6959674646331
+        323.0663727858372
+         873.988271868737
+ 8.36e+10    
+        886.2296031460721
+        325.4191530329414
+        769.5652155097205
+       -125.9831637762625
+        230.5791539763938
+        770.3402962424127
+       -222.3196132079278
+       -126.2766984855317
+        324.5876215185166
+        884.3189547068446
+ 8.41e+10    
+        896.6991073443485
+        326.9316912981097
+        777.9425245583436
+       -129.5756080618043
+        232.5804730441489
+        778.7136730714591
+       -224.7491209622853
+       -129.8691531092527
+        326.0929198600949
+        894.7629483824377
+ 8.46e+10    
+        907.2831341780276
+        328.4282436313107
+        786.4277697401402
+       -133.1800771238196
+        234.6378933038599
+        787.1944430686857
+       -227.1267634516531
+       -133.4728230066407
+        327.5822343268238
+        905.3211612562772
+ 8.51e+10    
+        917.9825397745666
+        329.9086858280409
+        795.0219054474589
+       -136.7960906866669
+        236.7524408485023
+        795.7835429974756
+       -229.4514689739459
+        -137.087242498432
+        329.0554382475879
+        915.9944432061521
+ 8.56e+10    
+        928.7981217205188
+        331.3727976015855
+        803.7257769536543
+       -140.4232095263745
+        238.9250310987649
+        804.4818009132655
+       -231.7222199865613
+       -140.7119883331267
+        330.5123089826654
+         926.783585723834
+ 8.61e+10    
+        939.7306192312695
+        332.8202598719535
+        812.5401195458817
+       -144.0610352084333
+        241.1564662154526
+        813.2899353455084
+       -233.9380531861042
+       -144.3466793906152
+        331.9525252305257
+        937.6893220925422
+ 8.66e+10    
+        950.7807134012701
+        334.2506521473807
+        821.4655578210791
+       -147.7092097511431
+        243.4474326381242
+        822.2085546471261
+       -236.0980595490346
+       -147.9909763103174
+        333.3756644273254
+        948.7123276459681
+ 8.71e+10    
+        961.9490275379243
+         335.663450004701
+        830.5026051494996
+       -151.3674152108373
+        245.7984987597597
+         831.238156505479
+       -238.2013843421036
+       -151.6445810413394
+        334.7812002448154
+        959.8532201101161
+ 8.76e+10    
+        973.2361275760582
+        337.0580226725752
+        839.6516633065257
+       -155.0353731915529
+        248.2101127375749
+        840.3791276299182
+       -240.2472271011233
+       -155.3072363132561
+          336.16850019144
+        971.1125600258048
+ 8.81e+10    
+        984.6425225770155
+         338.433630725332
+          848.91302227754
+       -158.7128442752908
+        250.6826004436449
+        849.6317436036381
+       -242.2348415872988
+       -158.9787250273464
+        337.5368233242445
+        982.4908512544897
+ 8.86e+10    
+         996.168665309714
+        339.7894238907086
+        858.2868602356983
+       -162.3996273699092
+        253.2161635628365
+        858.9961689160745
+       -244.1635357145319
+       -162.6588695645116
+         338.885318074553
+        993.9885415672708
+ 8.91e+10    
+        1007.814952915736
+        341.1244389797708
+        867.7732436943082
+       -166.0955589800286
+        255.8108778395287
+        868.4724571652001
+       -246.0326714642408
+       -166.3475310142788
+        340.2130201966877
+        1005.606023316608
+ 8.96e+10    
+        1019.581727658189
+        342.4375979439125
+        877.3721278403713
+       -169.8005123936813
+        258.4666914769317
+        878.0605514416693
+       -247.8416647790998
+        -170.044608315103
+        341.5188508423377
+        1017.343634192012
+ 9.01e+10    
+        1031.469277755543
+        343.7277060656136
+        887.0833570455964
+        -173.514396786346
+        261.1834236963273
+        887.7602848933935
+       -249.5899854421709
+       -173.7500373146192
+        342.8016147698984
+        1029.201658058819
+ 9.06e+10    
+        1043.477838299126
+        344.9934502896315
+        896.9066655644127
+       -177.2371562421393
+        263.9607634547615
+        897.5713814681221
+       -251.2771569476787
+       -177.4637897434403
+        344.0599986927859
+        1041.180325883011
+ 9.11e+10    
+        1055.607592256756
+        346.2333976997324
+        906.8416784126069
+       -180.9687686911991
+        266.7982683336559
+        907.4934568462668
+       -252.9027563573613
+       -181.1858721004613
+        345.2925697748582
+        1053.279816738592
+ 9.16e+10    
+         1067.85867156105
+        347.4459941500154
+         916.887912437614
+       -184.7092447606041
+        269.6953635933319
+        917.5260195540716
+       -254.4664141522391
+       -184.9163244557151
+        346.4977742788616
+        1065.500258901631
+ 9.21e+10    
+        1080.231158284322
+        348.6295630553018
+        927.0447775717973
+       -188.4586265419744
+         272.651341403188
+        927.6684722721143
+        -255.967814077428
+       -188.6552191628171
+        347.6739363748709
+        1077.841731028961
+ 9.26e+10    
+        1092.725085898583
+        349.7823043495168
+        937.3115782886161
+       -192.2169862722219
+        275.6653602530185
+        937.9201133257552
+       -257.4066929818276
+       -192.4026594838874
+        348.8192571154528
+        1090.304263422382
+ 9.31e+10    
+        1105.340440623521
+        350.9022936181117
+         947.687515238709
+       -195.9844249267244
+        278.7364445447819
+         948.280138376025
+       -258.7828406537914
+       -196.1587781293675
+        349.9318135840845
+        1102.887839378826
+ 9.36e+10    
+        1118.077162859542
+        351.9874814111342
+        958.1716870935311
+       -199.7610707288143
+        281.8634843728106
+         958.747642299714
+       -260.0960996566744
+       -199.9237357043187
+         351.009558226486
+        1115.592396627021
+ 9.41e+10    
+        1130.935148709267
+        353.0356927464325
+        968.7630925793873
+       -203.5470775684334
+        285.0452354948653
+        969.3216212671325
+        -261.346365159228
+       -203.6977190711775
+        352.0503183678537
+        1128.417828849639
+ 9.46e+10    
+        1143.914251585135
+        354.0446268077845
+        979.4606327166543
+       -207.3426233361866
+        288.2803195017435
+        980.0009750185695
+       -262.5335847684446
+       -207.4809396190549
+         353.051795928166
+        1141.363987293833
+ 9.51e+10    
+        1157.014283905488
+        355.0118568475203
+        990.2631132558282
+       -211.1479081689974
+        291.5672241838699
+        990.7845093380076
+       -263.6577583585971
+       -211.2736314465267
+        354.0115673391628
+        1154.430682466064
+ 9.56e+10    
+        1170.235018876971
+        355.9348303008927
+        1001.169247322311
+       -214.9631526075131
+        294.9043041041974
+         1001.67093873001
+        -264.718937903189
+       -215.0760494551725
+        354.9270836726309
+        1167.617685915544
+ 9.61e+10    
+        1183.576192366473
+        356.8108691189168
+        1012.177658261269
+       -218.7885956657196
+        298.2897813812817
+        1012.658889303786
+       -265.7172273013637
+       -218.8884673520925
+        355.7956709874877
+        1180.924732104301
+ 9.66e+10    
+        1197.037504858438
+        357.6371703286787
+        1023.286882695881
+       -222.6244928146085
+         301.721746682339
+        1023.746901848328
+       -266.6527822101125
+       -222.7111755651041
+        356.6145309031045
+        1194.351520363228
+ 9.71e+10    
+        1210.618623501572
+        358.4108068289372
+        1034.495373787648
+       -226.4711138753568
+        305.1981604388543
+        1034.933435131588
+       -267.5258098709298
+       -226.5444790685335
+        357.3807414068636
+        1207.897716936457
+ 9.76e+10    
+        1224.319184243113
+        359.1287284283157
+         1045.80150471443
+       -230.3287408264014
+         308.716854278008
+          1046.2168693928
+       -268.3365689337803
+        -230.388695119986
+        358.0912579039095
+        1221.562957111308
+ 9.81e+10    
+        1238.138794049761
+        359.7877631346493
+        1057.203572352939
+         -234.19766552453
+        312.2755326862501
+        1057.595510050359
+         -269.08536928512
+       -234.2441509097758
+        358.7429145165862
+        1235.346847435871
+ 9.86e+10    
+        1252.077033216671
+        360.3846187034838
+        1068.699801179065
+       -238.0781873352707
+        315.8717748985265
+        1069.067591615859
+       -269.7725718650129
+       -238.1111811218533
+        359.3324256418574
+        1249.248968021661
+ 9.91e+10    
+         1266.13345776342
+         360.915884454546
+        1080.288347382746
+       -241.9706106817553
+         319.503037026033
+        1080.631281822728
+       -270.3985884878276
+       -241.9901254072404
+        359.8563877776462
+         1263.26887493424
+ 9.96e+10    
+        1280.307601915954
+          361.37803336114
+        1091.967303192742
+       -245.8752425033744
+        323.1666544179608
+        1092.284685960965
+       -270.9638816509079
+       -245.8813257726803
+        360.3112816178383
+        1277.406102667696
+ 1.001e+11   
+        1294.598980676076
+        361.7674244269398
+        1103.734701425835
+       -249.7923896308679
+        326.8598442708673
+        1104.025851430169
+       -271.4689643420709
+       -249.7851238806845
+        360.6934744357495
+        1291.660166705786
+ 1.006e+11   
+        1309.007092475381
+        362.0803053504943
+        1115.588520244485
+       -253.7223560767347
+         330.579708481577
+         1115.85277249877
+       -271.9143998367701
+       -253.7018582675686
+        360.9992227531229
+        1306.030566167201
+ 1.011e+11   
+        1323.531421915457
+        362.3128154917842
+        1127.526688136896
+        -257.665440241985
+        334.3232367500311
+        1127.763395280701
+       -272.3008014862091
+       -257.6318614762945
+        361.2246753102593
+        1320.516786534895
+ 1.016e+11   
+        1338.171442590474
+        362.4609891451004
+        1139.547089113091
+       -261.6219320394273
+        338.0873099389961
+        1139.755622922349
+       -272.6288324985025
+       -261.5754571067506
+        361.3658763409123
+        1335.118302468652
+ 1.021e+11   
+        1352.926619996672
+        362.5207591290867
+        1151.647568118445
+       -265.5921099359563
+        341.8687036910554
+        1151.827321006688
+        -272.899205699725
+       -265.5329567832823
+        361.4187691622367
+        1349.834580700187
+ 1.026e+11   
+        1367.796414520154
+        362.4879606973967
+        1163.825936662259
+       -269.5762379136859
+        345.6640923049241
+        1163.976323160816
+        -273.112683290447
+        -269.504657045169
+        361.3792000846448
+        1364.665083010172
+ 1.031e+11   
+        1382.780284509668
+        362.3583357832017
+        1176.079978669324
+       -273.5745623528185
+        349.4700528772645
+        1176.200436883654
+       -273.2700765785812
+       -273.4908361556603
+        361.2429226538612
+        1379.609269284701
+ 1.036e+11   
+        1397.877689427582
+        362.1275375792347
+        1188.407456536812
+       -277.5873088363709
+        353.2830697151441
+        1188.497449581878
+       -273.3722457006995
+       -277.4917508357815
+        361.0056022268347
+        1394.666600650947
+ 1.041e+11   
+        1413.088093080278
+        361.7911354676556
+        1200.806117419601
+       -281.6146788780783
+         357.099539014805
+        1200.865134813644
+        -273.420099317303
+       -281.5076329218017
+        360.6628208941887
+         1409.83654269226
+ 1.046e+11   
+        1428.410966924871
+        361.3446202969805
+        1213.273699715588
+       -285.6568465798879
+        360.9157738176508
+        1213.301258737907
+        -273.414594294107
+       -285.5386859517579
+        360.2100827514196
+        1425.118568736498
+ 1.051e+11   
+        1443.845793454172
+        360.7834100244781
+         1225.80793977092
+        -289.713955211332
+        364.7280092396956
+        1225.803586775864
+       -273.3567353517591
+       -289.5850816784949
+        359.6428195291301
+        1440.512163220664
+ 1.056e+11   
+        1459.392069651377
+        360.1028557200302
+        1238.406578790193
+       -293.7861137253153
+        368.5324079819804
+        1238.369890469574
+       -273.2475746971349
+        -293.646956516271
+        358.9563965869762
+        1456.016825128741
+ 1.061e+11   
+        1475.049310519903
+        359.2982479462465
+        1251.067369956308
+        -297.873393202145
+        372.3250661180993
+        1250.997954542361
+       -273.0882116216613
+       -297.7244079210328
+        358.1461192783052
+         1471.63207149818
+ 1.066e+11   
+        1490.817052680533
+        358.3648235125936
+        1263.788085748635
+       -301.9758232306809
+        376.1020191648349
+        1263.685584158772
+       -272.8797920708613
+       -301.8174907058796
+        357.2072396911899
+        1487.357440996101
+ 1.071e+11   
+        1506.694858036311
+        357.2977726157086
+        1276.566525467789
+       -306.0933882269014
+        379.8592484397535
+        1276.430612374106
+       -272.6235081851322
+       -305.9262132984254
+        356.1349637689951
+        1503.192497561281
+ 1.076e+11   
+        1522.682317500968
+        356.0922463671384
+        1289.400522948395
+       -310.2260236930696
+        383.5926876929371
+        1289.230907775067
+       -272.3205977995425
+       -310.0505339405544
+        354.9244588186809
+        1519.136834108505
+ 1.081e+11   
+         1538.77905479022
+        354.7433647136525
+        1302.287954467599
+       -314.3736124218597
+        387.2982300347851
+        1302.084382303754
+       -271.9723439141219
+       -314.1903568325179
+        353.5708614094424
+        1535.190076293867
+ 1.086e+11   
+        1554.984730269385
+        353.2462247545431
+        1315.226746840153
+       -318.5359806483211
+        390.9717351391488
+        1314.988999259245
+       -271.5800741218128
+       -318.3455282304195
+        352.0692856647397
+        1551.351886338292
+ 1.091e+11   
+        1571.299044857575
+        351.5959094561439
+        1328.214885684823
+       -322.7128941515733
+        394.6090367360221
+        1327.942781476651
+       -271.1451599942104
+       -322.5158324940893
+        350.4148319520382
+         1567.62196690288
+ 1.096e+11   
+        1587.721743981462
+        349.7874967719622
+        1341.250423875465
+       -326.9040543149011
+        398.2059503824088
+        1340.943819662456
+       -270.6690164283025
+        -326.700988095846
+        348.6025959729886
+        1584.000065016465
+ 1.101e+11   
+        1604.252621578148
+        347.8160691619312
+        1354.331490146982
+       -331.1090941434627
+        401.7582815178467
+        1353.990280901837
+        -270.153100945996
+       -330.9006435895967
+        346.6276782531619
+        1600.485976048714
+ 1.106e+11   
+        1620.891524139105
+         345.676723521472
+        1367.456297869039
+       -335.3275742473596
+        405.2618337973937
+        1367.080417301407
+       -269.5989129434784
+       -335.1143735494088
+        344.4851940339912
+        1617.079547725025
+ 1.111e+11   
+        1637.638354794846
+        343.3645815083452
+        1380.623153959499
+       -339.5589787954164
+        408.7124176999318
+        1380.212574789351
+       -269.0079928987672
+       -339.3416744776427
+        342.1702835698622
+        1633.780684180633
+ 1.116e+11   
+        1654.493077430803
+        340.8748002777797
+        1393.830467943096
+       -343.8027114401517
+        412.1058594103335
+        1393.385202033907
+       -268.3819215189064
+       -343.5819606934787
+        339.6781228208125
+        1650.589350046526
+ 1.121e+11   
+        1671.455720834436
+        338.2025836168679
+        1407.076761138359
+       -348.0580912287858
+         415.438009965345
+        1406.596859491028
+        -267.722318844155
+       -347.8345602041927
+        337.0039345479632
+        1667.505574562955
+ 1.126e+11   
+        1688.526382862897
+        335.3431934750104
+        1420.360675960628
+       -352.3243484947911
+        418.7047546673609
+        1419.846228562388
+       -267.0308432851813
+       -352.0987105634734
+        334.1429998025708
+        1684.529455717299
+ 1.131e+11   
+        1705.705234629781
+        332.2919618903588
+        1433.680985333019
+       -356.6006207468192
+         421.902022751291
+         1433.13212085068
+       -266.3091906175567
+       -356.3735547306943
+        331.0906698067973
+        1701.661164396514
+ 1.136e+11   
+        1722.992524701231
+        329.0443033001386
+         1447.03660218603
+       -360.8859485548842
+        425.0257972950412
+        1446.453487495525
+       -265.5590929056846
+        -360.658136928419
+        327.8423782164913
+        1718.900948549656
+ 1.141e+11   
+        1740.388583297655
+        325.5957272334693
+        1460.426589040752
+        -365.179271442753
+        428.0721253834988
+        1459.809428588119
+       -264.7823173748599
+       -364.9513985124896
+        324.3936537650386
+        1736.249137356725
+ 1.146e+11   
+        1757.893826491374
+        321.9418513727855
+         1473.85016764986
+       -369.4794237979905
+        431.0371284872541
+        1473.199202636307
+       -263.9806652198536
+       -369.2521738591475
+        320.7401332752871
+        1753.706145393303
+ 1.151e+11   
+        1775.508760394896
+        318.0784149763548
+        1487.306728689141
+       -373.7851307991078
+         433.917013073526
+        1486.622236069546
+       -263.1559703538231
+       -373.5591862793049
+        316.8775750246634
+        1771.272476781966
+ 1.156e+11   
+        1793.233985330762
+        314.0012926484973
+         1500.79584147653
+       -378.0950043796714
+        436.7080814222037
+        1500.078132769475
+        -262.310098091895
+       -377.8710439641193
+        312.8018724623372
+        1788.948729330689
+ 1.161e+11   
+        1811.070199974235
+        309.7065084410691
+        1514.317263700983
+       -382.4075392258283
+        439.4067426322108
+        1513.566683600875
+        -261.444943770584
+       -382.1862359776121
+        308.5090682537315
+        1806.735598639018
+ 1.166e+11   
+        1829.018205462858
+        305.1902502768664
+        1527.870951145024
+       -386.7211088273764
+        442.0095238151629
+        1527.087875927634
+       -260.5624313086752
+       -386.5031283009026
+        303.9953686400594
+        1824.633882173918
+ 1.171e+11   
+        1847.078909457884
+        300.4488846635061
+        1541.457067376007
+        -391.033961587061
+        444.5130814468691
+        1540.641903091898
+       -259.6645117015624
+       -390.8199599375283
+        299.2571580957558
+        1842.644483297278
+ 1.176e+11   
+        1865.253330154933
+        295.4789716917304
+        1555.075993383312
+       -395.3442169978267
+        446.9142128663064
+        1554.229173838582
+       -258.7531614499358
+       -395.1348390946921
+        294.2910142599692
+        1860.768415242138
+ 1.181e+11   
+        1883.542600228532
+        290.2772802843902
+        1568.728337143193
+       -399.6498618996158
+        449.2098679019744
+         1567.85032164991
+       -257.8303809293553
+        -399.445739446349
+        289.0937231213117
+        1879.006805023761
+ 1.186e+11   
+        1901.947970701566
+        284.8408036725634
+        1582.414943079424
+       -403.9487468304436
+          451.39716059854
+        1581.506213982271
+       -256.8981926956978
+       -403.7504964939755
+        283.6622944285837
+        1897.360897275218
+ 1.191e+11   
+        1920.470814728559
+        279.1667750727208
+          1596.1369014003
+       -408.2385824786297
+        453.4733810282614
+        1595.197961364859
+       -255.9586397327996
+       -408.0468040326821
+        277.9939772972182
+         1915.83205799919
+ 1.196e+11   
+        1939.112631282359
+        273.2526835294984
+        1609.895557279115
+       -412.5169362506476
+        455.4360071518355
+         1608.92692634237
+       -255.0137836392643
+       -412.3322107386631
+        272.0862759857754
+        1934.421778220012
+ 1.201e+11   
+        1957.875048727227
+         267.096289890568
+        1623.692519852234
+       -416.7812289685014
+        457.2827167075786
+        1622.694732225766
+       -254.0657027606655
+       -416.6041168888211
+        265.9369657986042
+        1953.131677529266
+ 1.206e+11   
+        1976.759828274238
+        260.6956428774457
+        1637.529671004089
+       -421.0287317060972
+         459.011399095813
+        1636.503271631492
+       -253.1164902670003
+       -420.8597712252785
+        259.5441090846358
+        1971.963507507244
+ 1.211e+11   
+        1995.768867296148
+        254.0490952039852
+        1651.409173904225
+       -425.2565627846799
+        460.6201672279079
+        1650.354714766549
+       -252.1682521862759
+        -425.096267982733
+        252.9060712852594
+        1990.919155010247
+ 1.216e+11   
+        2014.904202495863
+        247.1553197062316
+        1665.333481272145
+       -429.4616849336479
+          462.10736929435
+        1664.251517433433
+       -251.2231053852338
+       -429.3105440852094
+        246.0215369903312
+        2010.000645311152
+ 1.221e+11   
+        2034.168012910402
+        240.0133254246689
+        1679.305343321244
+       -433.6409026386261
+        463.4716004295627
+        1678.196428722472
+       -250.2831755169601
+        -433.499376536779
+         238.889525947121
+        2029.210145074857
+ 1.226e+11   
+        2053.562622737261
+        232.6224735923397
+        1693.327815363431
+       -437.7908596872696
+        464.7117142163631
+         1692.19249835074
+       -249.3505949318246
+       -437.6593800112942
+         231.509408975172
+        2048.549965161605
+ 1.231e+11   
+        2073.090503968552
+        224.9824934675297
+        1707.404265020482
+       -441.9080369268743
+        465.8268339934754
+        1706.243083618468
+       -248.4275005629601
+       -441.7870046644948
+         223.880923725909
+        2068.022563234628
+ 1.236e+11   
+        2092.754278816327
+        217.0934979481237
+        1721.538379016317
+       -445.9887502553524
+        466.8163639160404
+        1720.351855935998
+        -247.516031785532
+        -445.878534178766
+        216.0041902226273
+        2087.630546165364
+ 1.241e+11   
+        2112.556721915349
+        208.9559989011086
+        1735.734169506381
+       -450.0291488554722
+        467.6799997161706
+        1734.522806894312
+       -246.6183282785943
+       -449.9300840592362
+         207.879726119801
+         2107.37667221488
+ 1.246e+11   
+        2132.500762286853
+         200.570922135836
+        1749.995979900345
+       -454.0252136900592
+        468.4177391103592
+        1748.760253831822
+       -245.7365278737786
+        -453.937600196934
+        199.5084616031228
+        2127.263852979831
+ 1.251e+11   
+        2152.589485045668
+        191.9396219406083
+        1764.328490143266
+       -457.9727562745964
+        469.0298917907547
+        1763.068844851935
+       -244.8727644198743
+       -457.8968577134737
+        190.8917538550981
+        2147.295155083199
+ 1.256e+11   
+        2172.826132837485
+        183.0638951012744
+        1778.736721402283
+       -461.8674177444256
+        469.5170889384202
+        1777.453563266487
+        -244.029165667608
+       -461.8034601046916
+        182.0314010072875
+        2167.473801597704
+ 1.261e+11   
+        2193.214106987428
+        173.9459943125372
+        1793.226040132549
+       -465.7046682282857
+        469.8802921949756
+        1791.919731403844
+       -243.2078511942312
+       -465.6528386994386
+        172.9296554821712
+        2187.803173183359
+ 1.266e+11   
+        2213.756968343704
+        164.5886408851666
+        1807.802161454579
+       -469.4798065483703
+        470.1208020075509
+        1806.473013750523
+       -242.4109303796066
+       -469.4402524497561
+        163.5892366366376
+        2208.286808922131
+ 1.271e+11   
+        2234.458437802375
+        154.9950366499925
+        1822.471151822727
+       -473.1879602586002
+        470.2402652885866
+        1821.119419380283
+        -241.640500444121
+       -473.1607880629106
+          154.01334260442
+        2228.928406836855
+ 1.276e+11   
+        2255.322396493795
+        145.1688749495016
+        1837.239430916862
+       -476.8240860385147
+         470.240682285013
+        1835.865303624271
+       -240.8986445849713
+       -476.8093604996578
+        144.2056612273826
+        2249.731824074423
+ 1.281e+11   
+        2276.352885617121
+        135.1143506016291
+        1852.113772735564
+       -480.3829704539611
+        470.1244125969311
+        1850.717368939226
+       -240.1874302100659
+       -480.3807138395163
+        134.1703799652666
+        2270.701076740894
+ 1.286e+11   
+        2297.554105906866
+        124.8361687147158
+         1867.10130582175
+       -483.8592310983568
+        469.8941802215207
+        1865.682664933598
+       -239.5089073070391
+       -483.8694225415499
+        123.9121946584288
+        2291.840339370562
+ 1.291e+11   
+        2318.930416715909
+        114.3395522246229
+        1882.209512593143
+       -487.2473181311192
+          469.55307754629
+        1880.768587501796
+       -238.8651069714175
+       -487.2698930992137
+        113.4363170183302
+        2313.153944016406
+ 1.296e+11   
+        2340.486334702336
+         103.630248017255
+         1897.44622772822
+       -490.5415162130555
+        469.1045681835985
+        1895.982877032175
+       -238.2580401058294
+       -490.5763661075875
+        102.7484807066775
+        2334.646378946168
+ 1.301e+11   
+        2362.226532103927
+        92.71453148967736
+        1912.819635556064
+       -493.7359468611585
+        468.5524885224488
+        1911.333615637516
+       -237.6896963410215
+       -493.7829187487615
+        91.85494586203896
+        2356.322286931779
+ 1.306e+11   
+          2384.1558345918
+         81.5992094020324
+        1928.338266425929
+       -496.8245712174439
+        467.9010478931162
+        1926.829223377274
+       -237.1620431961086
+       -496.8834677058889
+        80.76250192079557
+        2378.186463119676
+ 1.311e+11   
+        2406.279218689348
+        70.29162085504662
+        1944.010991997885
+       -499.8011932449765
+        467.1548272152028
+        1942.478453422861
+       -236.6770255152529
+       -499.8717725049734
+        69.47846857024349
+        2400.243852471819
+ 1.316e+11   
+         2428.60180874675
+        58.79963622526366
+        1959.847019422951
+       -502.6594633513146
+        466.3187759942443
+        1958.290386141302
+       -236.2365652273353
+       -502.7414392933838
+        58.01069466835281
+        2422.499546766031
+ 1.321e+11   
+        2451.128873467482
+        47.13165388263693
+        1975.855884386704
+       -505.3928824351734
+        465.3982075367163
+        1974.274422056596
+       -235.8425614516797
+        -505.485925049805
+        46.36755495399449
+        2444.958781151889
+ 1.326e+11   
+        2473.865821975614
+        35.29659449993479
+        1992.047442964619
+       -507.9948063576709
+        464.3987922237903
+        1990.440273654441
+       -235.4968910188804
+       -508.0985422219767
+        34.55794435527595
+         2467.62693025221
+ 1.331e+11   
+        2496.818199424757
+        23.30389276127755
+        2008.431862277581
+       -510.4584508260689
+        463.3265487055891
+        2006.797956015119
+       -235.2014094286088
+       -510.5724637857592
+        22.59126970989816
+        2490.509503810314
+ 1.336e+11   
+        2519.991682146116
+        11.16348626546479
+        2025.019609917992
+       -512.7768966808705
+        462.1878328358832
+        2023.357776245259
+       -234.9579523197891
+        -512.900728715008
+        10.47743868952121
+         2513.61214188243
+ 1.341e+11   
+        2543.392072339325
+       -1.114198591504441
+        2041.821442120297
+       -514.9430955682956
+        460.9893241939096
+        2040.130321693249
+       -234.7683374850701
+       -515.0762478377887
+       -1.773154287646392
+        2536.940609573665
+ 1.346e+11   
+        2567.025292312544
+       -13.51826397405483
+        2058.848390675164
+       -516.9498759746936
+        459.7380099974612
+         2057.12644693461
+       -234.6343675179667
+       -517.0918100668638
+       -14.14964536871078
+        2560.500791331554
+ 1.351e+11   
+        2590.897378277462
+        -26.0373614402284
+        2076.111748567593
+       -518.7899495972127
+        458.4411662331147
+        2074.357259530495
+       -234.5578331239445
+       -518.9400889679102
+       -26.64072204405068
+        2584.298684797454
+ 1.356e+11   
+        2615.014473721231
+       -38.65971648640148
+        2093.623054358085
+       -520.4559180166121
+        457.1063357961179
+        2091.834104558769
+       -234.5405172018783
+       -520.6136496319339
+       -39.23464761975251
+        2608.340394239756
+ 1.361e+11   
+        2639.382822366435
+       -51.37315705795559
+        2111.394075291547
+       -521.9402796247366
+        455.7413034390719
+        2109.568547927161
+       -234.5841997333552
+       -522.1049558144194
+       -51.91928964255854
+        2632.632123578804
+ 1.366e+11   
+        2664.008760749138
+       -64.16514627850631
+        2129.436789181545
+        -523.235436766197
+        454.3540673108762
+        2127.572358495943
+       -234.6906635855522
+       -523.4063772820282
+       -64.68215252898224
+         2657.18016903519
+ 1.371e+11   
+        2688.898710441385
+       -77.02281966917306
+        2147.763365075602
+       -524.3337030252742
+        452.9528068625609
+        2145.857489045328
+       -234.8617013053804
+       -524.5101973176809
+       -77.51041466337132
+        2681.990911427816
+ 1.376e+11   
+        2714.059169959998
+       -89.93302712799513
+        2166.386142764065
+       -525.2273106007286
+        451.5458468856544
+        2164.436056122547
+       -235.0991229927827
+       -525.4086203037562
+       -90.39097024204628
+        2707.070808159529
+ 1.381e+11   
+        2739.496706399158
+       -102.8823799540081
+        2185.317611175446
+       -525.9084176800729
+        450.1416174340657
+        2183.320318841453
+       -235.4047653467861
+       -526.0937793158245
+       -103.3104761399275
+        2732.426384933498
+ 1.386e+11   
+        2765.217946845813
+       -115.8573032034544
+        2204.570385734466
+       -526.3691157315046
+        448.7486093796309
+        2202.522656695128
+       -235.7805020036754
+       -526.5577436260592
+       -116.2554040897879
+        2758.064227254715
+ 1.391e+11   
+        2791.229569632472
+       -128.8440936729078
+         2224.15718477149
+       -526.6014366085514
+         447.375325338716
+        2222.055546482854
+         -236.22825526477
+       -526.7925260197477
+       -129.2120984673628
+        2783.990971773256
+ 1.396e+11   
+        2817.538295503348
+       -141.8289838113908
+        2244.090805085688
+       -526.5973593489603
+        446.0302256900438
+        2241.931538454032
+       -236.7500093243028
+       -526.7900898057096
+       -142.1668399800803
+        2810.213297540995
+ 1.401e+11   
+        2844.150878767746
+       -154.7982118652549
+        2264.384096794122
+       -526.3488165509373
+        444.7216694063719
+        2262.163231795351
+       -237.3478251489211
+       -526.5423553896562
+       -155.1059155664606
+        2836.737917263778
+ 1.406e+11   
+        2871.074098537128
+       -167.7380985656867
+        2285.049937597786
+       -525.8477001639724
+        443.4578494080894
+        2282.763249619912
+       -238.0238571098978
+       -526.0412062682074
+       -168.0156948091185
+        2863.571568633587
+ 1.411e+11   
+        2898.314750149402
+       -180.6351306643437
+        2306.101206665135
+       -525.0858665515668
+        442.2467221354421
+        2303.744213621158
+       -238.7803715271851
+       -525.2784942737211
+       -180.8827131742893
+         2890.72100585193
+ 1.416e+11   
+        2925.879636889636
+       -193.4760516407813
+        2327.550758295947
+       -524.0551406380749
+         441.095931027527
+        2325.118718598348
+       -239.6197672757266
+       -524.2460439024546
+       -193.6937623859677
+        2918.192991453308
+ 1.421e+11   
+        2953.775562150678
+       -206.2479598754144
+        2349.411395616982
+       -522.7473189461989
+        440.0127236004379
+        2346.899307077977
+       -240.5445985962003
+       -522.9356555141266
+       -206.4359882454095
+        2945.994288561761
+ 1.426e+11   
+        2982.009322164646
+       -218.9384146131158
+         2371.69584455074
+       -521.1541713085539
+        439.0038617880272
+        2369.098444288972
+       -241.5576002839944
+       -521.3391071925287
+       -219.0969961997879
+        2974.131653724376
+ 1.431e+11   
+        3010.587699477792
+       -231.5355500085712
+        2394.416728350486
+       -519.2674410193561
+        438.0755252229396
+        2391.728493779647
+       -242.6617154424376
+       -519.4481550317432
+       -231.6649649678932
+        3002.611830481451
+ 1.436e+11   
+        3039.517457342894
+       -244.0281975559672
+        2417.586543028535
+       -517.0788431648405
+        437.2332071177275
+        2414.801694010723
+       -243.8601259608226
+        -517.254531578149
+       -244.1287685083624
+        3031.441543854537
+ 1.441e+11   
+        3068.805335227111
+       -256.4060171867729
+        2441.217634033893
+       -514.5800608523612
+        436.4816024001381
+        2438.330136271029
+       -245.1562859288614
+       -514.7499421509224
+       -256.4781066278485
+        3060.627495942251
+ 1.446e+11   
+        3098.458045651768
+       -268.6596373155536
+        2465.322174587702
+       -511.7627390327754
+        435.8244877685541
+        2462.325744340942
+       -246.5539581831767
+       -511.9260587329362
+       -268.7036444915527
+        3090.176362844756
+ 1.451e+11   
+        3128.482272603505
+       -280.7808040871777
+         2489.91214612049
+       -508.6184755851656
+         435.264593308661
+        2486.800256331095
+       -248.0572541973023
+       -508.7745110973326
+       -280.7971613024915
+        3120.094793151025
+ 1.456e+11   
+        3158.884671774785
+       -292.7625400694806
+        2514.999321312838
+       -505.1388093073488
+        434.8034653309017
+         2511.76520920754
+       -249.6706775430349
+       -505.2868748080702
+       -292.7517083842654
+        3150.389408246879
+ 1.461e+11   
+        3189.671872917702
+       -304.5993126117579
+        2540.595250272845
+       -501.3152044250458
+        434.4413200750042
+        2537.231926535972
+       -251.3991711428055
+       -501.4546557174211
+       -304.5617768868226
+        3181.066804723832
+ 1.466e+11   
+        3220.850484617977
+       -316.2872120591296
+        2566.711250462385
+       -497.1390312114247
+        434.1768879500231
+        2563.211510047459
+       -253.2481685662917
+       -497.2692705307637
+        -316.223475307177
+        3212.133559196402
+ 1.471e+11   
+         3252.42710182244
+       -327.8241399847807
+        2593.358401015837
+       -492.6015422692555
+        434.0072479612555
+        2589.714835675647
+       -255.2236496141633
+       -492.7220230084008
+       -327.7347169855103
+        3243.596235857312
+ 1.476e+11   
+         3284.40831648086
+       -339.2100075694117
+        2620.547542183014
+         -487.69384400533
+        433.9276519965279
+         2616.75255478959
+       -257.3322004447764
+       -487.8040753213929
+       -339.0954176994748
+        3275.461397127257
+ 1.481e+11   
+        3316.800731688527
+       -350.4469442139558
+        2648.289280651271
+       -482.4068627953641
+        433.9313386556895
+        2644.335101372357
+       -259.5810785209935
+       -482.5064140623782
+       -350.3077034531003
+        3307.735617786094
+ 1.486e+11   
+        3349.610979747722
+       -361.5395164272796
+        2676.594001621412
+       -476.7313053005819
+        434.0093363151922
+        2672.472706021055
+       -261.9782826436151
+       -476.8198103672013
+       -361.3761284873963
+        3340.425502999137
+ 1.491e+11   
+        3382.845744595207
+       -372.4949569801499
+        2705.471888533965
+        -470.657612369266
+        434.1502551440222
+        2701.175417647882
+       -264.5326283567304
+       -470.7347735899777
+       -372.3079035178049
+        3373.537710680314
+ 1.496e+11   
+        3416.511789070775
+       -383.3234042621721
+        2734.932951447438
+       -464.1759059218613
+        434.3400677935481
+        2730.453133884859
+        -267.253829010807
+       -464.2414979194291
+       -383.1131341228343
+         3407.07897867066
+ 1.501e+11   
+         3450.61598754182
+       -394.0381517104246
+        2764.987065130446
+       -457.2759281886246
+         434.561878528246
+        2760.315641247279
+       -270.1525827853363
+       -457.3298013141642
+       -393.8050691610545
+        3441.056157232619
+ 1.506e+11   
+        3485.165364417577
+       -404.6559071165815
+        2795.644018022821
+       -449.9469726271757
+         434.795680577487
+        2790.772666190805
+       -273.2406659614149
+       -449.9890560802137
+       -404.4003590183132
+        3475.476247402757
+ 1.511e+11   
+        3520.167139134008
+        -415.197061536868
+        2826.913573286369
+       -442.1778058268935
+        435.0181015291266
+        2821.833938280182
+       -276.5310327484914
+       -442.2081104001157
+       -414.9193234131292
+         3510.34644576948
+ 1.516e+11   
+        3555.628778211212
+       -425.6859674495892
+        2858.805543274306
+       -433.9565796589893
+        435.2021366192549
+        2853.509266783403
+       -280.0379219718324
+        -433.975200079985
+       -425.3862284059427
+         3545.67419627718
+ 1.521e+11   
+        3591.558055022442
+       -436.1512257181313
+         2891.32987881257
+       -425.2707329123973
+        435.3168698213361
+        2885.808632061655
+       -283.7769709104855
+       -425.2778497505131
+       -435.8295721684589
+        3581.467249696387
+ 1.526e+11   
+        3627.963117947048
+       -446.6259808155506
+        2924.496774786514
+       -416.1068816169125
+        435.3271826826169
+        2918.742293254909
+       -287.7653366020346
+        -416.102762727954
+       -446.2823789733932
+        3617.733731417144
+ 1.531e+11   
+        3664.852567606342
+       -457.1482236648047
+        2958.316793629059
+        -406.450697223571
+        435.1934509005071
+        2952.320913802293
+       -292.0218248921974
+       -406.4356987158457
+       -456.7825007608158
+         3654.48221827131
+ 1.536e+11   
+        3702.235543915018
+       -467.7611013436241
+        2992.801008367435
+       -396.2867717886297
+        434.8712287176356
+        2986.555706473244
+       -296.5670275307484
+       -396.2613384877989
+       -467.3729255316977
+        3691.721825104982
+ 1.541e+11   
+        3740.121823706967
+       -478.5132327766337
+        3027.961167012271
+       -385.5984692744341
+         434.310921241357
+        3021.458599640438
+       -301.4234675747061
+        -385.563134680886
+        -478.102091693847
+        3729.462301855518
+ 1.546e+11   
+        3778.521929718589
+       -489.4590294230311
+        3063.809880125514
+       -374.3677620589901
+        433.4574449012925
+        3057.042426624968
+       -306.6157533696719
+       -374.3231477878847
+       -489.0242073724895
+        3767.714141915858
+ 1.551e+11   
+        3817.447251740488
+       -500.6590198302542
+        3100.360833530281
+       -362.5750517248488
+         432.249876306531
+        3093.321140038996
+       -312.1707413515156
+         -362.52186643153
+       -500.1995735608693
+        3806.488702588429
+ 1.556e+11   
+        3856.910180762294
+       -512.1801768005062
+        3137.629028173038
+       -350.1989731749156
+        430.6210898633541
+        3130.310053105049
+       -318.1177078971276
+        -350.138010970555
+       -511.6949098583144
+        3845.798338449937
+ 1.561e+11   
+          3896.9242569535
+        -524.096245765075
+         3175.63104925834
+       -337.2161811121846
+         428.497384592678
+        3168.026110046571
+       -324.4885304045193
+       -337.1483194855757
+       -523.5836814015466
+        3885.656548467543
+ 1.566e+11   
+        3937.504332334755
+       -536.4880728306198
+        3214.385366828079
+         -323.60111790825
+        425.7981006821674
+         3206.48818767955
+       -331.3178777901988
+       -323.5273151742888
+       -535.9464254543346
+        3926.078137713883
+ 1.571e+11   
+        3978.666748997444
+       -549.4439308112992
+        3253.912670030536
+       -309.3257618814691
+        422.4352264040408
+         3245.71743042022
+       -338.6434105179297
+        -309.247054183458
+       -548.8710759742718
+        3967.079394538634
+ 1.576e+11   
+        4020.429533726515
+       -563.0598414176623
+        3294.236237388469
+       -294.3593550057219
+        418.3129961330765
+          3285.7376209648
+       -346.5059902577259
+        -294.276852908393
+       -562.4532843415726
+        4008.678284044073
+ 1.581e+11   
+        4062.812609875388
+       -577.4398916299032
+        3335.382345392481
+       -278.6681090835578
+         413.327480287123
+        3326.575588940592
+       -354.9498992112782
+        -278.582993799089
+       -576.7967342730519
+        4050.894658716976
+ 1.586e+11   
+        4105.838027322482
+       -592.6965421406344
+        3377.380717806221
+       -262.2148894323402
+        407.3661681470393
+         3368.26165985164
+       -364.0230691007075
+       -262.1284087293362
+        -592.013448826712
+        4093.750487036123
+ 1.591e+11   
+        4149.530211311139
+       -608.9509256204353
+        3420.265018045017
+       -244.9588751568187
+        400.3075445860228
+          3410.8301466496
+       -373.7773197372075
+       -244.8723390083412
+       -608.2240872475555
+        4137.270100864347
+ 1.596e+11   
+         4193.91623093878
+       -626.3331324310778
+         3464.07338700277
+       -226.8551951267904
+        392.0206618654628
+        3454.319886240374
+       -384.2686070345149
+       -226.7699711596152
+       -625.5582292944639
+        4181.480462382332
+ 1.601e+11   
+        4239.026088009538
+       -644.9824812895661
+        3508.849028658306
+        -207.854538821208
+          382.36470775788
+        3498.774823215136
+       -395.5572802561545
+       -207.7720476365735
+       -644.1546445602382
+        4226.411451284009
+ 1.606e+11   
+        4284.893026904206
+       -665.0477722970337
+        3554.640845715676
+       -187.9027412745741
+        371.1885713414503
+        3544.244642995191
+       -407.7083481813906
+       -187.8244517072899
+       -664.1615442036933
+        4272.096172885023
+ 1.611e+11   
+        4331.553866041315
+       -686.6875196430634
+        3601.504127448243
+       -166.9403414283542
+         358.330407922415
+        3590.785456518728
+       -420.7917538084214
+        -166.867765827668
+       -685.7368124211616
+        4318.571287722001
+ 1.616e+11   
+        4379.049351414715
+       -710.0701612511399
+        3649.501291773635
+       -144.9021133095838
+        343.6172046208467
+        3638.460538428966
+       -434.8826570868592
+       -144.8368029120714
+       -709.0482149258196
+         4365.87736312551
+ 1.621e+11   
+        4427.424532578405
+       -735.3742425679601
+        3698.702683420526
+       -121.7165695535785
+        326.8643482380775
+        3687.341120569106
+       -450.0617250728289
+       -121.6601100364368
+       -734.2735816601656
+        4414.059247147239
+ 1.626e+11   
+        4476.729161322631
+       -762.7885717152791
+        3749.187429795093
+       -97.30543695200308
+        307.8751970841369
+        3737.507242336852
+       -466.4154287632484
+       -97.25944423990741
+       -761.6009609548281
+        4463.166465084624
+ 1.631e+11   
+        4527.018113139649
+       -792.5123432165908
+        3801.044355913159
+        -71.5831038642814
+        286.4406585050442
+        3789.048659213917
+       -484.0363457577229
+       -71.54922026854996
+       -791.2287423723764
+        4513.253638706357
+ 1.636e+11   
+        4578.351831398848
+       -824.7552275870921
+        3854.372959398311
+       -44.45603951665635
+        262.3387738890257
+        3842.065810398952
+       -503.0234677063572
+       -44.43593028578236
+       -823.3657455268146
+        4564.380928107381
+ 1.641e+11   
+        4630.796793966619
+       -859.7374241627173
+        3909.284446158248
+        -15.8221854605113
+        235.3343129452951
+        3896.670846122195
+       -523.4825113970364
+       -15.81753580288968
+       -858.2312722692037
+        4616.614495928538
+ 1.646e+11   
+        4684.426001776871
+       -897.6896746898755
+        3965.902826873295
+        14.42968029527461
+        205.1783790588927
+        3952.988714717585
+       -545.5262321305054
+        14.41716765042025
+       -896.0551197700253
+        4670.026993460159
+ 1.651e+11   
+         4739.31948861752
+       -938.8532353825902
+        4024.366073881748
+        46.42060566574921
+        171.6080275174828
+        4011.158308993776
+       -569.2747378679982
+        46.38921231929001
+       -937.0775522148094
+        4724.698067896963
+ 1.656e+11   
+        4795.564851120191
+        -983.479805390763
+        4084.827337408649
+         80.2821522222504
+        134.3458983563845
+        4071.333670809651
+       -594.8558024502978
+         80.2301453331288
+       -981.5492290719407
+        4780.714889741235
+ 1.661e+11   
+        4853.257797631062
+        -1031.83140992185
+        4147.456219360322
+        116.1571067386754
+        93.09986553145113
+        4133.685252056273
+       -622.4051759830246
+        116.0827396076518
+       -1029.731088171733
+        4838.172699039903
+ 1.666e+11   
+         4912.50271430557
+       -1084.180236583785
+         4212.44010208386
+        154.2002145829815
+        47.56270404686929
+        4198.401229405045
+       -652.0668902837231
+        154.1017265925437
+        -1081.89418218502
+        4897.175368804893
+ 1.671e+11   
+        4973.413246386644
+       -1140.808423931577
+        4279.985528562962
+        194.5789324963518
+       -2.588223410657649
+        4265.688869300063
+       -683.9935570715608
+        194.4545484297303
+       -1138.319467481511
+        4957.835983589159
+ 1.676e+11   
+        5036.112892225016
+        -1202.00780163226
+        4350.319629498182
+         237.474197763909
+       -57.69125888454531
+        4335.775938627761
+       -718.3466563577887
+        237.3221265606976
+       -1199.297544788424
+        5020.277430780972
+ 1.681e+11   
+        5100.735607138322
+       -1268.079582173285
+         4423.69159155438
+        283.0812101789737
+       -118.1007192705896
+        4408.912155372334
+       -755.2968122884914
+         282.899643217332
+       -1265.128351576657
+        5084.633001728573
+ 1.686e+11   
+        5167.426413725749
+       -1339.334004567439
+        4500.374159836394
+          331.61022253768
+       -184.1871429034935
+        4485.370672337909
+       -795.0240534646166
+        331.3973315772855
+       -1336.120806626469
+        5151.046999320807
+ 1.691e+11   
+         5236.34201471892
+       -1416.089931100449
+        4580.665166240051
+        383.2873346659877
+       -256.3375114838018
+        4565.449585638374
+       -837.7180545472538
+        383.0412696411702
+       -1412.592407813785
+        5219.675348117604
+ 1.696e+11   
+        5307.651403880221
+       -1498.674398770238
+        4664.889073872016
+        438.3552851791166
+       -334.9554462891548
+        4649.473458215622
+       -883.5783557554864
+        438.0741720936442
+       -1494.868784761119
+        5290.686202558794
+ 1.701e+11   
+        5381.536469847489
+       -1587.422127702456
+        4753.398526115644
+        497.0742342899792
+        -420.461377692272
+        4737.794847044565
+       -932.8145566602417
+        496.7561735444818
+       -1583.283208621021
+        5364.260548167398
+ 1.706e+11   
+        5458.192587171291
+       -1682.674989462491
+        4846.575887221695
+        559.7225300339462
+       -513.2926870125683
+        4830.795821020603
+       -985.6464805094801
+        559.3655956116518
+       -1678.176061902246
+        5440.592790017762
+ 1.711e+11   
+        5537.829188105207
+       -1784.781438816785
+        4944.834759514028
+        626.5974492331495
+       -613.9038197114304
+        4928.889454748388
+       -1042.304305141641
+        626.1996892933383
+        -1779.89427186344
+         5519.89132205511
+ 1.716e+11   
+        5620.670307981582
+       -1894.095913103474
+        5048.621460402705
+        698.0159034179396
+       -722.7663688448017
+        5032.521281585767
+       -1103.028656416752
+         697.575342983387
+       -1888.790711611936
+        5602.379070135947
+ 1.721e+11   
+        5706.955096259136
+       -2010.978203934119
+         5158.41644047172
+        774.3150987122929
+        -840.369127506058
+        5142.170687388014
+        -1168.07066000701
+        773.8297453353897
+       -2005.223573595315
+        5688.294000917408
+ 1.726e+11   
+        5796.938284555399
+       -2135.792806447967
+        5274.735621907796
+        855.8531374122342
+       -967.2181087273106
+        5258.352224434511
+       -1237.691947275573
+         855.320990926253
+       -2129.555720661604
+        5777.889587964013
+ 1.731e+11   
+        5890.890602188173
+        -2268.90825175646
+        5398.131634551804
+        943.0095476037811
+       -1103.836530920545
+        5381.616823037234
+       -1312.164610983134
+        942.4286153690564
+        -2262.15402028302
+        5871.435225659737
+ 1.736e+11   
+        5989.099128967829
+       -2410.696428515913
+        5529.194924853579
+         1036.18572569896
+       -1250.764766442456
+        5512.552876376523
+       -1391.771106549699
+        1035.554045134366
+       -2403.388667819558
+        5969.216580754251
+ 1.741e+11   
+        6091.867574199152
+       -2561.531899745746
+         5668.55471111018
+        1135.805275175871
+       -1408.560250221444
+        5651.787172197015
+       -1476.804094666538
+        1135.120945864111
+        -2553.63250486884
+        6071.535870603131
+ 1.746e+11   
+        6199.516470100573
+        -2721.79122102551
+        5816.879756521274
+        1242.314223110592
+       -1577.797344621562
+        5799.985643186659
+       -1567.566221167624
+        1241.575451412916
+        -2713.26033875642
+        6178.712056440098
+ 1.751e+11   
+        6312.383267126764
+       -2891.852266055801
+        5974.878929934306
+        1356.181094190488
+       -1759.067155795583
+        5957.853906178132
+        -1664.36983024535
+        1355.386254176703
+       -2882.648269050185
+         6291.08093933194
+ 1.756e+11   
+        6430.822318017552
+       -3072.093565213728
+        6143.301522676943
+        1477.896819827767
+       -1952.977295725926
+        6126.137558845935
+       -1767.536607326301
+        1477.044535472818
+       -3062.173026608033
+        6408.995145844298
+ 1.761e+11   
+        6555.204736780517
+        -3262.89366219082
+         6322.93728864374
+        1607.974457561884
+       -2160.151583007254
+         6305.62220129115
+       -1877.397148223889
+        1607.063712730545
+       -3252.211330098911
+        6532.823989895856
+ 1.766e+11   
+         6685.91811827837
+       -3464.630493008644
+        6514.616173903327
+        1746.948693110091
+       -2381.229674125634
+         6497.13314896779
+       -1994.290451572595
+        1745.978977981524
+       -3453.139264105374
+         6662.95319681914
+ 1.771e+11   
+        6823.366103598393
+       -3677.680790715787
+         6719.20770152874
+        1895.375093894443
+       -2616.866615698651
+        6701.534802726679
+       -2118.563331981617
+        1894.346599429466
+        -3665.33168186553
+        6799.784475270394
+ 1.776e+11   
+        6967.967775931572
+       -3902.419517804717
+        6937.619977185939
+        2053.829078367239
+       -2867.732306780482
+        6919.729641452326
+       -2250.569751907823
+        2052.742954548282
+       -3889.161634379541
+        6943.734922343735
+ 1.781e+11   
+        7120.156871207971
+       -4139.219326903844
+        7170.798281269911
+        2222.904559428892
+       -3134.510859056597
+        7152.656802789589
+       -2390.670070867987
+        2221.763258821643
+        -4124.99982600352
+        7095.236247006662
+ 1.786e+11   
+        7280.380787138965
+       -4388.450048536091
+        7419.723214012989
+        2403.212211895517
+       -3417.899841591521
+        7401.290217730887
+       -2539.230211360065
+          2402.0199484194
+         -4373.2140947313
+        7254.733796731603
+ 1.791e+11   
+         7449.09937341395
+       -4650.478202692984
+        7685.408360968165
+        2595.377302114288
+       -3718.609395835004
+        7666.636265309329
+       -2696.620741707692
+        2594.140666954018
+       -4634.168913082636
+        7422.685371831917
+ 1.796e+11   
+        7626.783484313954
+       -4925.666528588969
+        7968.897447431317
+         2800.03700054976
+       -4037.361205978454
+        7949.730913969879
+       -2863.215877031057
+        2798.765794789881
+       -4908.224902784346
+        7599.559811347342
+ 1.801e+11   
+        7813.913272442986
+       -5214.373524134241
+        8271.260951438251
+        3017.837072543188
+       -4374.887309543417
+        8251.636316027098
+       -3039.392400639153
+        3016.545442262865
+       -5195.738353060639
+        7785.835333027158
+ 1.806e+11   
+        8010.976197869097
+       -5516.952983190962
+        8593.592145500932
+        3249.427803907125
+       -4731.928733439217
+        8573.436820194582
+       -3225.528509343299
+        3248.135802736446
+        -5497.06072808287
+        7981.997607550724
+ 1.811e+11   
+        8218.464719449741
+       -5833.753514197148
+        8937.002536443162
+        3495.458959376786
+       -5109.233941696845
+        8916.234363264502
+       -3422.002587440662
+        3494.194723160098
+       -5812.538143429423
+        8188.537542764878
+ 1.816e+11   
+        8436.873622420979
+       -6165.118017586692
+        9302.616669320774
+        3756.573481951368
+       -5507.557082692809
+         9281.14319368912
+        -3629.19191519857
+        3755.376291840329
+       -6142.510783380812
+        8405.948746130831
+ 1.821e+11   
+        8666.696915142884
+       -6511.383090395193
+        9691.566253432036
+        4033.399502211547
+       -5927.656025720153
+        9669.283863766779
+       -3847.471318190796
+        4032.324154839151
+       -6487.312219033426
+        8634.724620656889
+ 1.826e+11   
+        8908.424192785269
+       -6872.878312352792
+        10104.98355263834
+         4326.54001180038
+       -6370.290178564756
+        10081.77639813011
+       -4077.211762784033
+         4325.66313778762
+        -6847.26856885941
+        8875.355028038968
+ 1.831e+11   
+        9162.536308142217
+       -7249.925344649579
+        10543.99395360545
+        4636.559224795292
+       -6836.218077492295
+        10519.73249589174
+       -4318.778898213887
+        4635.988545534407
+       -7222.697414068754
+        9128.322417304047
+ 1.836e+11   
+        9429.500096623446
+       -7642.836733175449
+         11009.7075765467
+        4963.964152976119
+       -7326.194734260841
+        10984.24653935854
+       -4572.531531977652
+        4963.852206798046
+       -7613.906333425414
+        9394.097259958668
+ 1.841e+11   
+        9709.761756396072
+       -8051.914238981712
+        11503.20971322441
+        5309.179211320138
+       -7840.968700650064
+        11476.38504664504
+       -4838.819991235175
+        5309.743892967985
+       -8021.190844271571
+        9673.132542218795
+ 1.846e+11   
+         10003.7382713247
+       -8477.446395590425
+        12025.54975552278
+        5672.510798957995
+       -8381.278743480629
+        11997.17400453723
+       -5117.984242069455
+        5674.066171536801
+       -8444.831412157489
+          9965.8569287917
+ 1.851e+11   
+        10311.80601015536
+       -8919.704772680192
+        12577.72811721988
+        6054.098239543464
+       -8947.849849428625
+        12547.58327625812
+       -5410.351449680215
+        6057.100217876234
+       -8885.089008114219
+        10272.66602967241
+ 1.856e+11   
+        10634.28555368225
+       -9378.938042563921
+        13160.68051940425
+        6453.849206900717
+       -9541.387848019662
+        13128.50720123894
+       -5716.232224410953
+         6458.96034267174
+       -9342.198484492468
+        10593.91103245736
+ 1.861e+11   
+        10971.42281037361
+       -9855.362344192445
+        13775.25922029328
+        6871.368859686899
+       -10162.57089902863
+        13740.74147631252
+       -6035.913795800059
+        6879.538610580781
+       -9816.359063929422
+        10929.88411085429
+ 1.866e+11   
+        11323.37188616111
+       -10349.14582302918
+        14422.21246592701
+         7305.93501225457
+       -10812.03368285696
+        14384.96162940437
+       -6369.646169289388
+        7318.456285792635
+       -10307.72259358745
+         11280.8016238329
+ 1.871e+11   
+        11690.20533066124
+       -10860.38627804123
+        15102.17030385562
+        7756.710832114448
+       -11490.33523611039
+        15061.72792052564
+       -6717.613233977977
+        7775.090441438644
+       -10816.38674481634
+        11646.79294568027
+ 1.876e+11   
+         12072.0368260386
+       -11389.09151103133
+         15815.6671604365
+        8223.750564856327
+       -12197.89521913936
+        15771.59928206528
+       -7079.877013373014
+          8248.8930373367
+       -11342.42225949612
+        12027.92560837261
+ 1.881e+11   
+         12469.4502967331
+       -11935.21828374393
+        16563.28840186668
+        8710.880695278898
+       -12934.89549766014
+        16515.54557175002
+       -7456.299993565697
+        8740.554306380838
+       -11886.01078639271
+        12424.35783318661
+ 1.886e+11   
+        12884.32465974596
+       -12498.93550080009
+        17346.10282686703
+        9230.322791530565
+       -13701.24950941798
+        17295.74884212434
+       -7846.554551652156
+        9254.840753159206
+       -12447.76485508634
+        12836.79485332476
+ 1.891e+11   
+        13319.92715058571
+       -13081.21777658137
+        18166.33703028491
+        9801.040907940671
+       -14496.95757409583
+        18115.70150282549
+       -8250.502167360546
+        9804.092106824832
+       -13028.91561572589
+        13267.21856651964
+ 1.896e+11   
+        13778.19257974728
+       -13683.93519485407
+        19027.11886324233
+        10430.10162808083
+       -15322.83443638186
+        18977.55145794883
+       -8668.833305673901
+        10404.40697901522
+       -13630.60059452891
+         13718.6450938943
+ 1.901e+11   
+        14257.29477537703
+       -14308.28179354772
+        19929.91942850836
+        11101.09662316367
+       -16180.43753022707
+        19879.69516355358
+       -9102.849216720804
+        11058.86278488674
+       -14252.91647489992
+        14192.43122590356
+ 1.906e+11   
+        14754.18875415351
+       -14953.64335333929
+         20872.9502192511
+        11793.92060515724
+       -17070.92867012264
+        20819.25416112491
+       -9553.358622731956
+        11751.49820731539
+       -14895.23032230542
+        14686.58855205893
+ 1.911e+11   
+        15267.33943456907
+       -15618.80312955145
+        21853.57746564921
+        12500.48041281785
+       -17994.56047100516
+        21794.77736295417
+        -10020.3282192056
+        12465.30673890247
+       -15556.93538781044
+        15198.31833252928
+ 1.916e+11   
+        15796.53180933298
+        -16303.0991220887
+        22870.45013508012
+        13221.17835105852
+       -18951.11452902969
+        22806.05539006407
+       -10503.38094977206
+        13193.72180634326
+       -16237.73892996644
+        15726.22798168437
+ 1.921e+11   
+        16341.98643741965
+       -17006.40507059805
+        23923.26977349597
+        13958.70022752034
+       -19940.32044404283
+        23853.23820353897
+       -11002.17905022352
+        13937.16174590203
+       -16937.59595301795
+        16270.08739236627
+ 1.926e+11   
+        16903.92257269026
+       -17728.80642543841
+        25012.04342328904
+        14715.43240656358
+        -20961.9608106244
+        24936.40221987375
+       -11516.49319096755
+        14697.93593667424
+       -17656.56710102637
+        16830.05348526484
+ 1.931e+11   
+        17482.44265383054
+       -18470.41825483318
+        26136.70832524761
+        15492.97133914381
+       -22015.84265793281
+        26055.43910230056
+       -12046.16054474943
+        15478.10000707856
+       -18394.72817090219
+        17406.28172767158
+ 1.936e+11   
+        18077.52845709921
+        -19231.3239289427
+        27297.02937819872
+        16292.24017831969
+       -23101.75622417685
+        27210.05503522287
+          -12591.04170582
+        16279.02202890327
+       -19152.13237800154
+        17998.81926955156
+ 1.941e+11   
+        18689.06173953944
+       -20011.56266579113
+        28492.59611075148
+        17113.68286007825
+        -24219.4484637569
+        28399.79387105877
+       -13150.99544275792
+        17101.47019264787
+       -19928.79924188961
+        18607.59997395148
+ 1.946e+11   
+        19316.84474852876
+       -20811.13144983097
+         29722.8435339288
+        17957.41529432156
+       -25368.60947456651
+        29624.06024204264
+        -13725.8663963491
+        17945.77768092649
+       -20724.71353318339
+        19232.46325882821
+ 1.951e+11   
+        19960.61615462383
+       -21629.98971498122
+        30987.07432280056
+        18823.32679186326
+       -26548.86676558903
+        30882.13855356279
+       -14315.47987835972
+         18811.9758881624
+       -21539.82723908877
+        19873.17357123489
+ 1.956e+11   
+        20620.06296785941
+       -22468.06369048994
+        32284.47779488311
+        19711.14579170181
+       -27759.78395048866
+        32173.20853140414
+       -14919.64028632039
+        19699.88611196944
+       -22374.06208837977
+        20529.43589727869
+ 1.961e+11   
+        21294.82970730913
+       -23325.24990070737
+        33614.14588739235
+        20620.48289313928
+       -29000.86199912182
+        33496.35858860076
+       -15538.13135081907
+        20609.18023921667
+       -23227.31193451165
+        21200.90758577493
+ 1.966e+11   
+        21984.52583915119
+       -24201.41795971002
+        34975.08711607255
+        21550.86000677215
+       -30271.54207068733
+        34850.59797402186
+       -16170.71733729749
+        21539.42121694059
+       -24099.44488272783
+        21887.20756989404
+ 1.971e+11   
+        22688.73215060472
+       -25096.41289042405
+        36366.23932654713
+        22501.73108055431
+       -31571.20940652757
+        36234.86829608398
+       -16817.14476618289
+        22490.09091399567
+       -24990.30520992929
+        22587.92389990044
+ 1.976e+11   
+        23407.00646317162
+       -26010.05715203624
+        37786.48175279553
+        23472.49767347459
+       -32899.19798207789
+        37648.05474139862
+       -17477.14442544855
+        23460.61019486168
+       -25899.71514982608
+        23302.62020118901
+ 1.981e+11   
+        24138.88891463059
+        -26942.1524984221
+        39234.64666149791
+        24462.52131913301
+       -34254.79572355242
+         39088.9971293227
+       -18150.43354965557
+        24450.35414587149
+       -26827.47660079322
+        24030.84143419096
+ 1.986e+11   
+        24883.90693041291
+       -27892.48174157089
+        40709.53070222413
+        25471.13382744574
+       -35637.25014536306
+        40556.50083232583
+        -18836.7180875557
+        25458.66422085204
+       -27773.37279258927
+        24772.11917272766
+ 1.991e+11   
+        25641.57993868995
+       -28860.81046002312
+         42209.9059838493
+        26497.64619996299
+       -37045.77428832824
+        42049.34752550418
+       -19535.69500394726
+        26484.85836132934
+        -28737.1699300245
+        25525.97651628208
+ 1.996e+11   
+        26411.42384404436
+       -29846.88866998843
+        43734.53083822104
+         27541.3565517332
+       -38479.55285075923
+        43566.30569060644
+       -20247.05457364567
+        27528.23971772839
+       -29718.61881846202
+        26291.93268986679
+ 2.001e+11   
+        27192.95525201551
+       -30850.45246273276
+        45282.16019919796
+        28601.55726306795
+       -39937.74841153841
+         45106.1407805378
+       -20970.48263232816
+        28588.10433975817
+       -30717.45646721908
+         27069.5073485483
+ 2.006e+11   
+        27985.69542493169
+        -31871.2256033738
+        46851.55550962402
+        29677.54148284736
+       -41419.50764978878
+        46667.62494323638
+       -21705.66275359791
+         29663.7480485001
+       -31733.40766157039
+        27858.22458301804
+ 2.011e+11   
+        28789.17394444087
+       -32908.92108162136
+        48441.49406476984
+        30768.60904465385
+       -42923.96747131017
+        48249.54620508449
+       -22452.27832529429
+        30754.47260924746
+       -32766.18649126525
+        28657.61661206133
+ 2.016e+11   
+        29602.93205560936
+       -33963.24260302167
+        50050.77770445369
+        31874.07182227338
+       -44450.26095837334
+        49850.71702103297
+       -23210.01450151312
+         31859.5912688276
+       -33815.49782257459
+        29467.22714371352
+ 2.021e+11   
+        30426.52566982353
+       -35033.88600906687
+        51678.24077494922
+        32993.25853242607
+       -45997.52306695798
+         51469.9821095839
+       -23978.56001027107
+        32978.43368952473
+       -34881.03870134939
+        30286.61438698607
+ 2.026e+11   
+        31259.52800794318
+       -36120.54061557367
+        53322.75729410683
+        34125.51898407502
+       -47564.89600407706
+        53106.22550439335
+       -24757.60880033998
+        34110.35029496235
+       -35962.49967599524
+        31115.35369877209
+ 2.031e+11   
+        32101.53187048855
+       -37222.89046053355
+        54983.24726758469
+        35270.22777158046
+       -49151.53422727042
+        54758.37676949943
+       -25546.86151447265
+        35254.71603589421
+       -37059.56603132462
+        31953.03985488601
+ 2.036e+11   
+        32952.15152757602
+       -38340.61545496115
+        56658.68211972443
+        36426.78741089912
+       -50756.60901845909
+        56425.41634127642
+        -26346.0267799948
+        36410.93358229809
+       -38171.91892669271
+        32799.28893944855
+ 2.041e+11   
+        33811.02422743983
+       -39473.39243279776
+        58348.08921862924
+        37594.63092234206
+       -52379.31259482303
+        58106.37997647229
+       -27154.82231145537
+        37578.43595017077
+       -39299.23643444484
+        33653.73985248793
+ 2.046e+11   
+        34677.81132840519
+       -40620.89609853445
+        60050.55549079818
+        38773.22386900961
+       -54018.86172993697
+        59800.36230158036
+        -27972.9758236353
+         38756.6885754797
+       -40441.19447734986
+        34516.05544132533
+ 2.051e+11   
+        35552.19906487413
+       -41782.79987372483
+         61765.2301357368
+        39962.06586614458
+       -55674.50086879016
+        61506.51947386921
+       -28800.22575662496
+         39945.1908528006
+       -41597.46766620415
+        35385.92326677235
+ 2.056e+11   
+         36433.8989630847
+       -42958.77664586606
+        63491.32646491018
+        41160.69158274965
+       -57345.50473027835
+        63224.07097828915
+       -29636.32181782532
+        41143.47716156152
+       -42767.73004111044
+        36263.05602019125
+ 2.061e+11   
+         37322.6479269773
+       -44148.49942514854
+        65228.12290192928
+        42368.67126252794
+       -59031.18040007774
+        64952.30059691398
+       -30481.02534854185
+         42351.1174080337
+       -43951.65572193419
+         37147.1916119145
+ 2.066e+11   
+        38218.20801837162
+       -45351.64191625118
+        66974.96319174573
+        43585.61079626566
+       -60730.86892530489
+        66690.55659835995
+       -31334.10952528661
+        43567.71711593343
+        -45148.9194751106
+        38038.09295529078
+ 2.071e+11   
+        39120.36595877075
+       -46567.87901366706
+          68731.255875745
+        44811.15138202377
+       -62443.94642990494
+        68438.25120363022
+       -32195.35940793962
+        44792.91710251034
+       -46359.19720525187
+        38935.54747366374
+ 2.076e+11   
+        40028.93238245496
+       -47796.88722996486
+        70496.47309689707
+        46044.96881284508
+       -64169.82477619737
+        70194.85939200092
+        -33064.5718485445
+        46026.39278017876
+       -47582.16638091562
+        39839.36635988141
+ 2.081e+11   
+        40943.74087210398
+       -49038.34506692219
+        72270.14880454259
+        47286.77243406435
+       -65907.95180337162
+        71959.91711588419
+       -33941.55527570471
+        47267.85312601899
+        -48817.5064043985
+        40749.38361946784
+ 2.086e+11   
+         41864.6468090386
+       -50291.93333964475
+        74051.87643201502
+        48536.30381375417
+       -67657.81117797254
+        73733.01899714417
+       -34826.12937033353
+        48517.03936284747
+       -50064.89893558084
+        41665.45492941198
+ 2.091e+11   
+         42791.5260703357
+       -51557.33546362188
+         75841.3061222105
+        49793.33517037334
+        -69418.9218945442
+        75513.81557918803
+       -35718.12464889985
+        49773.72339603978
+       -51324.02817967765
+        42587.45634467246
+ 2.096e+11   
+        43724.27360461462
+       -52834.23771422049
+        77638.14157655036
+        51057.66760137353
+       -71190.83746665499
+        77302.01020943004
+        -36617.3819703364
+        51037.70604994992
+       -52594.58114827806
+        43515.28288402758
+ 2.101e+11   
+         44662.8019172883
+       -54122.32946741734
+        79442.13660169466
+        52329.12915545687
+       -72973.14484959049
+          79097.355625608
+       -37523.75198247872
+         52308.8151466882
+       -53876.24790235615
+        44448.84702589046
+ 2.106e+11   
+        45607.03949459703
+       -55421.30342967626
+        81253.09142602785
+        53607.57278944978
+       -74765.46313614634
+        80899.65031707649
+       -38437.09452331275
+        53586.90346828304
+       -55168.72178503269
+        45388.07714323376
+ 2.111e+11   
+        46556.92919387759
+       -56730.85586382709
+        83070.84885454284
+         54892.8742484735
+       -76567.44206628708
+        82708.73472880182
+       -39357.27799147954
+        54871.84664096357
+       -56471.69965081721
+        46332.91590490717
+ 2.116e+11   
+        47512.42662534946
+       -58050.68681666465
+        84895.29032648406
+        56184.92990535931
+       -78378.76039007257
+        84524.48737153057
+       -40284.17869945704
+           56163.54097757
+       -57784.88209692238
+        47283.31866846982
+ 2.121e+11   
+        48473.49854830222
+       -59380.50035278425
+        86726.33193516279
+        57483.65459218013
+       -80199.12412129894
+        86346.82089668213
+       -41217.68022165935
+        57461.90131102152
+        -59107.9737010447
+        48239.25188727016
+ 2.126e+11   
+        49440.12130201786
+       -60720.00479796714
+        88563.92046391354
+        58788.97945345278
+       -82028.26471687856
+        88175.67818910613
+       -42157.67274840568
+        58766.85884846165
+       -60440.68326881108
+        49200.69155197181
+ 2.131e+11   
+        50412.27928912859
+       -62068.91299424514
+        90408.02948637966
+        60100.84984710005
+       -83865.93721418928
+        90011.02852511308
+       -43104.05245535445
+        60078.35907223659
+       -61782.72409291275
+        50167.62168410445
+ 2.136e+11   
+        51389.96352646219
+       -63426.94256765523
+        92258.65557336877
+        61419.22331573961
+       -85711.91835558471
+        91852.86383729124
+       -44056.72089661142
+        61396.35971034675
+       -63133.81422483973
+        51140.03289658528
+ 2.141e+11   
+        52373.17027581157
+       -64793.81620865731
+        94115.81464253324
+        62744.06764736191
+        -87566.0047260502
+        93701.19512169807
+       -45015.58442834146
+        62720.82879550925
+       -64493.67675910785
+        52117.92103356039
+ 2.146e+11   
+        53361.89976453424
+       -66169.26196425926
+        95979.53848122843
+        64075.35904103689
+        -89428.0109267135
+        95556.04901717624
+        -45980.5536683586
+        64051.74282854774
+       -65862.04012894299
+         53101.2858993971
+ 2.151e+11   
+         54356.1550034785
+       -67553.01354007608
+        97849.87146719146
+        65413.08039000721
+       -91297.76780364514
+        97417.46458090151
+       -46951.54299587932
+        65389.08505854964
+       -67238.63841159557
+        54090.13008427033
+ 2.156e+11   
+        55355.94070748244
+        -68944.8106098784
+        99726.86750624946
+        66757.21969143418
+       -93175.12074818982
+        99285.49027890284
+       -47928.47009440864
+        66732.84388913486
+       -68623.21164078792
+        55084.45789154683
+ 2.161e+11   
+         56361.2623216077
+       -70344.39912962353
+          101610.58720116
+        68107.76858917701
+       -95059.92808198303
+        101160.1812052572
+       -48911.25553959933
+        68083.01141729963
+       -70015.50612325383
+        56084.27437010521
+ 2.166e+11   
+        57372.12515439393
+       -71751.53165255736
+        103501.0952609851
+        69464.72105336434
+       -96952.05953691198
+        103041.5965390277
+       -49899.82243291102
+         69439.5821086714
+        -71415.2747559354
+        57089.58445286545
+ 2.171e+11   
+        58388.53361773332
+       -73165.96764168124
+        105398.4581561093
+        70828.07219813787
+       -98851.39483756659
+         104929.797243785
+       -50894.09608097955
+        70802.55161063316
+       -72822.27734011736
+        58100.39220112867
+ 2.176e+11   
+        59410.49057149703
+       -74587.47377571954
+        107302.7420201746
+        72197.81723685411
+       -100757.8223912571
+        106824.8440107782
+       -51894.00371981594
+         72171.9157026769
+       -74236.28088863382
+        59116.70015287198
+ 2.181e+11   
+         60437.9967697763
+       -76015.82424466813
+        109214.0107968118
+        73573.95057219485
+       -102671.2380884311
+        108726.7954434835
+       -52899.47428227004
+        73547.66938150805
+       -75657.05992223442
+        60138.50877188356
+ 2.186e+11   
+        61471.05040454215
+        -77450.8010310628
+        111132.3246261157
+        74956.46501708124
+       -104591.5442143459
+        110635.7064783786
+       -53910.43820662943
+         74929.8060768617
+       -77084.39675126283
+        61165.81599357323
+ 2.191e+11   
+        62509.64674165742
+       -78892.19417324521
+        113057.7384633053
+        76345.35114097975
+        -106518.648471114
+        112551.6270343396
+        -54926.8272837652
+        76318.31699268313
+       -78518.08173895036
+        62198.61686243167
+ 2.196e+11   
+        63553.77784349023
+        -80339.8020071278
+        114990.3009199376
+        77740.59673513321
+       -108452.4631077545
+        114474.6008810211
+       -55948.57453988009
+        77713.19056726046
+        -79957.9135428516
+        63236.90325543121
+ 2.201e+11   
+        64603.43237186453
+       -81793.43138324446
+        116930.0533163646
+        79142.18638942218
+       -110392.9041546357
+        116404.6647149448
+       -56975.61415165818
+        79114.41204507007
+       -81403.69933124464
+        64280.66368515472
+ 2.206e+11   
+        65658.59546472772
+       -83252.89785621538
+        118877.0289328126
+        80550.10117295128
+        -112339.890757676
+        118341.8474307467
+       -58007.88139044472
+        80521.96315247421
+       -82855.25497165836
+        65329.88317608373
+ 2.211e+11   
+        66719.24867969569
+       -84718.02584412761
+        120831.2524454998
+        81964.31841003078
+       -114293.3446068575
+         120286.169574095
+       -59045.31259199312
+        81935.82186898567
+       -84312.40518907127
+        66384.54320726352
+ 2.216e+11   
+        67785.36999754746
+       -86188.64875574344
+        122792.7395335433
+        83384.81154297991
+       -116253.1894529953
+        122237.6429621576
+       -60087.84514829698
+        83355.96228555984
+        -85774.9836917315
+        67444.62171447316
+ 2.221e+11   
+         68856.9338787642
+       -87664.60908387188
+        124761.4966420355
+        84811.55007308669
+       -118219.3507062737
+        124196.2704571425
+       -61135.41751806834
+        84782.35454128294
+       -87242.83326297838
+        68510.09314505193
+ 2.226e+11   
+        69933.91136631582
+       -89145.75846366544
+        126737.5208865149
+        86244.49957109445
+       -120191.7551097712
+        126162.0458782992
+       -62187.96925251424
+        86214.96482985275
+       -88715.80581786679
+         69580.9285586437
+ 2.231e+11   
+        71016.27022810173
+       -90631.95769503836
+        128720.8000841476
+        87683.62174874822
+        -122170.330481075
+        128134.9540378726
+       -63245.44103320599
+         87653.7554674061
+       -90193.76242383392
+        70657.09576732053
+ 2.236e+11   
+         72103.9751327089
+       -92123.07672881837
+        130711.3128971706
+        89128.87458317973
+       -124155.0055150572
+        130114.9708867483
+       -64307.77471900685
+        89098.68501349031
+       -91676.57328505836
+        71738.55950880228
+ 2.241e+11   
+        73196.98785246864
+       -93618.99461665156
+        132709.0290745702
+        90580.21248624474
+       -126145.7096409826
+          132102.06375595
+       -65374.91339922792
+        90549.70843730462
+       -93164.11769056894
+        72825.28164680679
+ 2.246e+11   
+        74295.26748815051
+       -95119.59942505925
+        134713.9097784852
+        92037.58651131816
+        -128142.372927292
+        134096.1916806792
+       -66446.80145040521
+        92006.77732172662
+       -94656.28392653883
+        73917.22139291688
+ 2.251e+11   
+        75398.77071001918
+       -96624.78811440716
+        136725.9079824622
+        93500.94459049593
+       -130144.9260276537
+        136097.3057942187
+       -67523.38459432808
+        93469.84009807724
+       -96152.96915355492
+        75014.33554473624
+ 2.256e+11   
+        76507.45201039159
+       -98134.46638387362
+        138744.9689293955
+        94970.23179563286
+       -132153.3001621877
+        138105.3497797291
+       -68604.60995519931
+        94938.84230505639
+       -97654.07924998121
+        76116.57873551489
+ 2.261e+11   
+        77621.26396325097
+       -99648.54848380125
+        140771.0306377455
+        96445.39061714357
+       -134167.4271281097
+        140120.2603687257
+       -69690.42611405505
+        96413.72686577454
+       -99159.52862282518
+         77223.9036908389
+ 2.266e+11   
+        78740.15748690159
+       -101166.9569970818
+         142804.024445433
+        97926.36125501379
+       -136187.2393344383
+         142141.967875823
+       -70780.78315882508
+        97894.43437732289
+       -100669.2399877796
+        78336.26148840567
+ 2.271e+11   
+        79864.08210607617
+       -102689.6225914539
+        144843.8755816313
+        99413.08191698618
+       -138212.6698558037
+        144170.3967601493
+       -71875.63272866167
+        99380.90340784086
+       -102183.1441203398
+        79453.60181732608
+ 2.276e+11   
+        80992.98621032135
+       -104216.4837447922
+        146890.5037575114
+        100905.4891194034
+       -140243.6525008268
+        146205.4662046653
+       -72974.92805140234
+        100873.0707965542
+       -103701.1795800887
+        80575.87323380957
+ 2.281e+11   
+        82126.81730589508
+       -105747.4864456233
+        148943.8237678203
+        102403.5179866961
+       -142280.1218909512
+        148247.0907054335
+       -74078.62397326111
+          102370.87195276
+       -105223.2924104006
+        81703.02341048964
+ 2.286e+11   
+        83265.52225880283
+       -107282.5838712451
+        151003.7460960011
+        103907.1025460009
+       -144322.0135460476
+        150295.1806637074
+       -75186.67698006288
+        103874.2411502325
+       -106749.4358159452
+         82834.9993770374
+ 2.291e+11   
+        84409.04752696639
+       -108821.7360459096
+        153070.1775163414
+        105416.1760138566
+       -146369.2639735089
+        152349.6429744772
+       -76299.04520953349
+        105383.1118139832
+       -108279.5698204628
+        83971.74775007486
+ 2.296e+11   
+        85557.33937987598
+       -110364.9094816129
+        155143.0216874209
+        106930.6710723889
+       -148421.8107579757
+        154410.3816058852
+       -77415.68845435233
+          106897.41679677
+       -109813.6609073527
+        85113.21495075364
+ 2.301e+11   
+        86710.34410440132
+       -111912.0768040617
+        157222.1797318496
+         108450.520132806
+       -150479.5926492037
+         156477.298164632
+         -78536.568155842
+        108417.0886431626
+       -111351.6816456474
+        86259.34740868419
+ 2.306e+11   
+        87868.00819574665
+       -113463.2163664097
+        159307.5507979931
+        109975.6555844367
+        -152542.549645965
+         158550.292443195
+       -79661.64738833134
+        109942.0598393787
+       -112893.6103039627
+        87410.09175121016
+ 2.311e+11   
+        89030.27853281026
+       -115018.3118533373
+        161399.0326000295
+        111506.0100278984
+       -154610.6230742134
+        160629.2629453122
+       -80790.89083436198
+        111472.2630474604
+       -114439.4304549909
+        88565.39497729318
+ 2.316e+11   
+        90197.10253747094
+        -116577.351878019
+        163496.5219333018
+        113041.5164913335
+       -156683.7556580741
+        162714.1073867998
+       -81924.26475103803
+        113007.6313227121
+       -115989.1305730765
+         89725.2046155329
+ 2.321e+11   
+        91368.42831755476
+       -118140.3295744679
+        165599.9151624962
+        114582.1086289577
+       -158761.8915825198
+        164804.7231693292
+       -83061.73692792511
+        114548.0983136248
+       -117542.7036273534
+        90889.46886607636
+ 2.326e+11   
+        92544.20479343945
+       -119707.2421876719
+         167709.108680702
+        116127.7209014403
+       -160844.9765468617
+        166901.0078252986
+       -84203.27663699409
+        116093.5984437897
+       -119100.1466728489
+        92058.13672637183
+ 2.331e+11   
+        93724.38180844352
+       -121278.0906638517
+        169823.9993378913
+        117678.2887378982
+       -162932.9578084475
+        169002.8594324163
+       -85348.85457518582
+        117644.0670755632
+       -120661.4604418697
+         93231.1581009107
+ 2.336e+11   
+        94908.91022330805
+       -122852.8792430664
+        171944.4848377983
+        119233.7486795039
+        -165025.784216179
+        171110.1769970399
+       -86498.44280023637
+        119199.4406554676
+       -122226.6489378862
+        94408.48389525947
+ 2.341e+11   
+        96097.74199521649
+       -124431.6150562809
+        174070.4641025668
+        120794.0385049052
+       -167123.4062336641
+        173222.8608057011
+       -87652.01466044816
+        120759.6568415054
+       -123795.7190340113
+        95590.06609481956
+ 2.346e+11   
+        97290.83024192022
+       -126014.3077288809
+        176201.8376048967
+        122359.0973378295
+       -169225.7759520001
+        175340.8127445956
+       -88809.54471913238
+        122324.6546127447
+       -125368.6800780482
+        96775.85782887533
+ 2.351e+11   
+         98488.1292916399
+       -127600.9689925014
+        178338.5076677401
+        123928.8657373934
+        -171332.847092346
+        177463.9365871311
+        -89971.0086744741
+         123894.374361679
+       -126945.5435059522
+        97965.81342058908
+ 2.356e+11   
+        99689.59471948938
+        -129191.612306882
+        180480.3787318652
+        125503.2857717621
+       -173444.5749985691
+        179592.1382498933
+       -91136.38327558216
+        125468.7579699884
+       -128526.3224654098
+        99159.88842368078
+ 2.361e+11   
+        100895.1833712425
+       -130786.2524933339
+        182627.3575918649
+         127082.301075909
+       -175560.9166203777
+        181725.3260176305
+       -92305.64623549454
+        127047.7488684386
+       -130111.0314510995
+        100358.0396465991
+ 2.366e+11   
+        102104.8533753029
+       -132384.9053812496
+        184779.3536013862
+        128665.8568943071
+       -177681.8304874387
+        183863.4107380611
+        -93478.7761419013
+        128631.2920817348
+       -131699.6859530493
+        101560.2251650348
+ 2.371e+11   
+        103318.5641437862
+       -133987.5874689452
+        186936.2788485503
+        130253.9001094602
+       -179807.2766750736
+        186006.3059874932
+       -94655.75236634034
+        130219.3342592202
+       -133292.3021193683
+        102766.4043236693
+ 2.376e+11   
+        104536.2763636327
+       -135594.3155999758
+        189098.0483026716
+        131846.3792572155
+       -181937.2167621703
+        188153.9282083728
+       -95836.55497259604
+        131811.8236923532
+       -134888.8964344726
+        103976.5377280685
+ 2.381e+11   
+        105757.9519786914
+       -137205.1066559174
+        191264.5799335181
+        133443.2445298508
+       -184071.6137820166
+        190306.1968200189
+        -97021.1646250081
+        133408.7103199369
+        -136489.485413786
+        105190.5872276437
+ 2.386e+11   
+        106983.5541637092
+        -138819.977266468
+        193435.7948044566
+        135044.4477679382
+       -186210.4321667826
+        192463.0343038857
+       -98209.56249736722
+        135009.9457220974
+       -138094.0853157534
+        106408.5158906063
+ 2.391e+11   
+        108213.0472911573
+       -140438.9435375754
+        195611.6171408998
+        136649.9424420032
+       -188353.6376864109
+        194624.3662647765
+       -99401.73018303759
+        136615.4831040134
+       -139702.7118718605
+        107630.2879718301
+ 2.396e+11   
+        109446.3968918019
+       -142062.0207981636
+        197791.9743755335
+        138259.6836249903
+       -190501.1973826776
+        196790.1214694777
+       -100597.6496069056
+        138225.2772704002
+       -141315.3800352157
+         108855.868874519
+ 2.401e+11   
+        110683.5696099124
+       -143689.2233658967
+        199976.7971718477
+        139873.6279565408
+       -192653.0794991999
+        198960.2318643349
+       -101797.3029397154
+        139839.2845917438
+       -142932.1037481246
+        110085.2251065578
+ 2.406e+11   
+        111924.5331539601
+       -145320.5643322867
+         202166.019427505
+         141491.733600061
+       -194809.2534081447
+        201134.6325732937
+       -103000.6725153027
+        141457.4629632542
+       -144552.8957289495
+        111318.3242323899
+ 2.411e+11   
+         113169.256243633
+       -146956.0553673334
+        204359.5782591038
+        143113.9601935392
+       -196969.6895343921
+        203313.2618779487
+       -104207.7407511931
+        143079.7717574897
+       -146177.7672784306
+        112555.1348212317
+ 2.416e+11   
+        114417.7085539507
+       -148595.7065437666
+        206557.4139698829
+        144740.2687950341
+       -199134.3592778797
+        205496.0611811354
+       -105418.4900729865
+        144706.1717715646
+       -147806.7281055315
+        113795.6263923997
+ 2.421e+11   
+        115669.8606572159
+       -150239.5261808434
+        208759.4700018909
+        146370.6218237156
+       -201303.2349348253
+        207682.9749555718
+       -106632.9028428945
+        146336.6251698193
+       -149439.7861727529
+        115039.7693584744
+ 2.426e+11   
+        116925.6839635013
+       -151887.5207075618
+        210965.6928741358
+        148004.9829973034
+       -203476.2896185013
+        209873.9506790458
+       -107850.9612927541
+        147971.0954227881
+       -151076.9475607652
+        116287.5349669894
+ 2.431e+11   
+        118185.1506603155
+       -153539.6945450393
+        213176.0321081724
+        149643.3172666939
+       -205653.4971801861
+        212068.9387575869
+       -109072.6474617895
+        149609.5472432549
+       -152718.2163521056
+        117538.8952412806
+ 2.436e+11   
+        119448.2336520474
+       -155196.0500077275
+        215390.4401425676
+        151285.5907485292
+       -207834.8321308989
+        214267.8924380439
+       -110297.9431393484
+        151251.9465201427
+        -154363.594533604
+        118793.8229210849
+ 2.441e+11   
+        120714.9064997362
+       -156856.5872230429
+         217608.872237614
+        152931.7706563997
+       -210020.2695644585
+        216470.7677114111
+       -111526.8298127906
+         152898.260250928
+       -156013.0819171118
+        120052.2914034291
+ 2.446e+11   
+        121985.1433616626
+       -158521.3040689174
+        219831.2863716201
+        154581.8252313268
+       -212209.7850823842
+        218677.5232082166
+       -112759.2886206598
+        154548.4564732225
+       -157666.6760780348
+        121314.2746842943
+ 2.451e+11   
+        123258.9189352122
+       -160190.1961287093
+        222057.6431300481
+        156235.7236721236
+       -214403.3547211046
+        220888.1200872141
+       -113995.3003112319
+        156202.5041961189
+       -159324.3723111104
+        122579.7473015031
+ 2.456e+11   
+        124536.2084004036
+       -161863.2566628439
+        224287.9055887021
+        157893.4360661681
+       -216600.9548818905
+         223102.521918559
+       -115234.8452064809
+        157860.3733318336
+       -160986.1636027913
+        123848.6842792147
+ 2.461e+11   
+        125816.9873654344
+       -163540.4765965032
+        226522.0391921106
+        159554.9333210836
+       -218802.5622638924
+        225320.6945625913
+       -116477.9031714735
+        159522.0346281414
+       -162652.0406195617
+        125121.0610743748
+ 2.466e+11   
+        127101.2318145441
+       -165221.8445226368
+        228760.0116281857
+        161220.1870977629
+       -221008.1538006116
+        227542.6060452767
+       -117724.4535891602
+        161187.4596020374
+       -164321.9917114496
+         126396.853525417
+ 2.471e+11   
+        128388.9180584513
+       -166907.3467195171
+        231001.7927001627
+        162889.1697451259
+       -223217.7066000906
+        229768.2264312949
+       -118974.4753404942
+        162856.6204750182
+       -165996.0029299695
+        127676.0378034678
+ 2.476e+11   
+        129680.0226875748
+       -168596.9671820319
+        233247.3541967732
+        164561.8542369473
+       -225431.1978890656
+        231997.5276956905
+       -120227.9467897807
+        164529.4901103186
+       -167674.0580596803
+        128958.5903662616
+ 2.481e+11   
+        130974.5225282112
+       -170290.6876658773
+        235496.6697615203
+        166238.2141110543
+       -227648.6049612818
+        234230.4835949482
+       -121484.8457751251
+        166206.0419524059
+        -169356.138662532
+         130244.487914937
+ 2.486e+11   
+        132272.3946017956
+       -171988.4877437876
+        237749.7147618781
+        167918.2234111356
+       -229869.9051301276
+        236467.0695382694
+       -122745.1496038206
+        167886.2499689763
+       -171042.2241341349
+        131533.7073538386
+ 2.491e+11   
+        133573.6160873399
+       -173690.3448729217
+        240006.4661591481
+        169601.8566313719
+       -232095.0756857111
+        238707.2624597813
+       -124008.8350524939
+        169570.0885956655
+       -172732.2917710808
+         132826.225753418
+ 2.496e+11   
+        134878.1642871049
+       -175396.2344725156
+        242266.9023796679
+        171289.0886640513
+       -234324.0938564558
+        240951.0406923298
+       -125275.8783717972
+        171257.5326836392
+       -174426.3168484235
+        134122.0203162882
+ 2.501e+11   
+        136186.0165955304
+        -177106.130010901
+        244531.0031879809
+        172979.8947502987
+       -236556.9367752641
+        243198.3838434586
+       -126546.2552954255
+        172948.5574501963
+       -176124.2727064287
+        135421.0683464593
+ 2.506e+11   
+        137497.1504714164
+        -178820.003100984
+        246798.7495625289
+        174674.2504340046
+       -238793.5814502577
+        245449.2726741026
+       -127819.9410532077
+        174643.1384324768
+       -177826.1308456907
+        136723.3472217448
+ 2.511e+11   
+        138811.5434133232
+       -180537.8236032881
+        249070.1235743687
+        176372.1315190191
+       -241034.0047400758
+         247703.688980481
+        -129096.910388016
+        176341.2514443393
+       -179531.8610297257
+        138028.8343693111
+ 2.516e+11   
+        140129.1729381288
+       -182259.5597356648
+        251345.1082693539
+        178073.5140296312
+       -243278.1833336821
+        249961.6154796071
+       -130377.1375762173
+        178042.8725364372
+       -181241.4313941521
+        139337.5072443089
+ 2.521e+11   
+        141450.0165626648
+       -183985.1781887877
+        253623.6875541706
+        179778.3741743363
+       -245526.0937346006
+         252223.035698784
+       -131660.5964513848
+        179747.9779594971
+       -182954.8085615779
+        140649.3433115085
+ 2.526e+11   
+        142774.0517883248
+       -185714.6442465586
+        255905.8460865636
+        181486.6883128603
+       -247777.7122494752
+        254487.9338694023
+       -132947.2604309759
+        181456.5441307785
+       -184671.9577613339
+        141964.3200298389
+ 2.531e+11   
+        144101.2560885291
+       -187447.9219105759
+        258191.5691700469
+         183198.432926397
+       -250033.0149808372
+        256756.2948253136
+       -134237.1025456806
+        183168.5476036682
+        -186392.842953206
+        143282.4148397129
+ 2.536e+11   
+        145431.6068989067
+       -189184.9740278267
+        260480.8426533305
+        184913.5845909779
+       -252291.9778239178
+         259028.103905994
+       -135530.0954711371
+         184883.965040343
+       -188117.4269543377
+         144603.605153007
+ 2.541e+11   
+         146765.081610048
+        -190925.762420798
+        262773.6528346729
+        186632.1199538931
+       -254554.5764673542
+        261303.3468646873
+       -136826.2115617113
+        186602.7731874169
+       -189845.6715685026
+        145927.8683455499
+ 2.546e+11   
+        148101.6575626663
+       -192670.2480192149
+        265069.9863713054
+          188354.01571305
+       -256820.7863975959
+        263582.0097816602
+       -138125.4228860362
+        188324.9488544705
+       -191577.5377169664
+        147255.1817519623
+ 2.551e+11   
+        149441.3120450015
+       -194418.3909926564
+        267369.8301940564
+         190079.248599155
+       -259090.5829068212
+        265864.0789826754
+       -139427.7012640099
+        190050.4688953501
+       -193312.9855701885
+        148585.5226626861
+ 2.556e+11   
+         150784.022292288
+       -196170.1508833136
+        269673.1714272523
+        191807.7953605808
+       -261363.9411041462
+        268149.5409627471
+       -140733.0183049535
+        191779.3101921069
+       -195051.9746796426
+        149918.8683230288
+ 2.561e+11   
+        152129.7654881062
+       -197925.4867381948
+        271979.9973139461
+        193539.6327507801
+       -263640.8359299126
+        270438.3823152155
+       -142041.3454466326
+        193511.4496414413
+       -196794.4641090641
+        151255.1959340461
+ 2.566e+11   
+        153478.5187674353
+       -199684.3572401168
+        274290.2951464944
+        195274.7375180942
+       -265921.2421728153
+        272730.5896661415
+       -143352.6539948607
+        195246.8641435077
+       -198540.4125644682
+        152594.4826550852
+ 2.571e+11   
+        154830.2592212172
+       -201446.7208368446
+        276604.0522024718
+        197013.0863978003
+       -268205.1344896412
+        275026.1496140032
+       -144666.9151633986
+        196985.5305929272
+       -200289.7785223126
+        153936.7056078064
+ 2.576e+11   
+        156184.9639022516
+       -203212.5358677879
+        278921.2556858883
+        198754.6561062333
+       -270492.4874273659
+         277325.048674638
+       -145984.1001138831
+        198727.4258718545
+        -202042.520355214
+        155281.8418815005
+ 2.581e+11   
+        157542.6098322322
+       -204981.7606876899
+        281241.8926736517
+        200499.4233368241
+       -272783.2754473691
+        279627.2732313703
+       -147304.1799955227
+        200472.5268449401
+       -203798.5964546656
+        156629.8685395241
+ 2.586e+11   
+        158903.1740097451
+       -206754.3537867843
+        283565.9500671942
+        202247.3647578811
+       -275077.4729515105
+         281932.809490222
+        -148627.125984309
+         202220.810356025
+       -205557.9653502316
+        157980.7626266747
+ 2.591e+11   
+        160266.6334190509
+       -208530.2739069283
+        285893.4145491658
+        203998.4570119547
+       -277375.0543098199
+        284241.6434401029
+       -149952.9093215077
+        203972.2532264125
+       -207320.5858247372
+        159334.5011773318
+ 2.596e+11   
+        161632.9650394786
+       -210309.4801532621
+        288224.2725450792
+        205752.6767166192
+       -279675.9938895468
+        286553.7608178532
+       -151281.5013512017
+        205726.8322545539
+       -209086.4170250057
+         160691.061224198
+ 2.601e+11   
+        163002.1458552624
+       -212091.9321009718
+         290558.510189773
+        207510.0004665061
+       -281980.2660853168
+        288869.1470779949
+       -152612.8735566721
+        207484.5242169927
+       -210855.4185677286
+        162050.4198074752
+ 2.606e+11   
+        164374.1528656642
+       -213877.5898967785
+        292896.1132985537
+        209270.4048364357
+       -284287.8453501493
+        291187.7873670418
+       -153946.9975954203
+        209245.3058704129
+       -212627.5506400922
+        163412.5539843225
+ 2.611e+11   
+        165748.9630952284
+       -215666.4143548054
+        295237.0673428556
+        211033.8663854858
+       -286598.7062270863
+        293509.6665022002
+       -155283.8453326428
+        211009.1539546435
+       -214402.7740948198
+        164777.4408384476
+ 2.616e+11   
+        167126.5536040243
+       -217458.3670465117
+        297581.3574302579
+        212800.3616618554
+       -288912.8233811947
+        295834.7689542914
+       -156623.3888729897
+        212776.0451964717
+       -216181.0505393214
+        166145.0574896921
+ 2.621e+11   
+        168506.9014977455
+       -219253.4103844184
+        299928.9682886854
+        214569.8672083722
+       -291230.1716317018
+        298163.0788347107
+       -157965.6005904482
+        214545.9563141293
+       -217962.3424186788
+        167515.3811034809
+ 2.626e+11   
+        169889.9839375356
+         -221051.50769938
+        302279.8842546083
+        216342.3595685114
+       -293550.7259840315
+        300494.5798862354
+       -159310.4531562097
+        216318.8640223161
+       -219746.6130922252
+        168888.3889000133
+ 2.631e+11   
+        171275.7781494299
+       -222852.6233111969
+        304634.0892650613
+        218117.8152927947
+        -295874.461661519
+        302829.2554774928
+       -160657.9195643935
+        218094.7450376383
+       -221533.8269035144
+        170264.0581630855
+ 2.636e+11   
+        172664.2614333063
+       -224656.7225923871
+        306991.5668532896
+        219896.2109454476
+       -298201.3541365843
+        305167.0886008898
+       -162007.9731555147
+        219873.5760843424
+       -223323.9492435044
+        171642.3662484444
+ 2.641e+11   
+        174055.4111712495
+       -226463.7720249718
+         309352.300147827
+        221677.5231111967
+        -300531.379161148
+        307508.0618738023
+       -163360.5876375961
+        221655.3339002312
+       -225116.9466068088
+        173023.2905915772
+ 2.646e+11   
+         175449.204835249
+       -228273.7392501591
+        311716.2718748145
+         223461.728402108
+       -302864.5127960944
+        309852.1575428313
+       -164715.7371048446
+        223439.9952426662
+       -226912.7866409055
+        174406.8087148633
+ 2.651e+11   
+        176845.6199941519
+       -230086.5931108395
+         314083.464363363
+        225248.8034643601
+       -305200.7314395772
+        312199.3574909176
+       -166073.3960538196
+        225227.5368945549
+       -228711.4381882123
+        175792.8982340112
+ 2.656e+11   
+        178244.6343198149
+       -231902.3036868293
+        316453.8595537627
+        227038.7249848694
+       -307540.0118539858
+        314549.6432471191
+       -167433.5393970402
+        227017.9356702431
+        -230512.871320976
+        177181.5368637267
+ 2.661e+11   
+        179646.2255923986
+       -233720.8423228366
+        318827.4390083456
+        228831.4696976843
+       -309882.3311913896
+        316902.9959988494
+        -168796.142473992
+        228811.1684212333
+       -232317.0573689401
+        178572.7024225611
+ 2.666e+11   
+        181050.3717047673
+       -235542.1816491351
+        321204.1839248076
+        230627.0143900772
+       -312227.6670172934
+        319259.3966063811
+       -170161.1810595021
+        230607.2120416604
+       -234123.9689397854
+        179966.3728369019
+ 2.671e+11   
+        182457.0506659633
+       -237366.2955949689
+        323584.0751517978
+        232425.3359082732
+       -314575.9973325384
+         321618.825619419
+       -171528.6313694718
+        232406.0434734658
+        -235933.579932362
+        181362.5261440772
+ 2.676e+11   
+        183866.2406037331
+       -239193.1593947238
+         325967.093206585
+        234226.4111627588
+       -316927.3005931973
+        323981.2632955486
+       -172898.4700639652
+        234207.6397112199
+       -237745.8655427498
+        182761.1404945579
+ 2.681e+11   
+         185277.919766102
+       -241022.7495869317
+        328353.2182946199
+        236030.2171331299
+       -319281.5557283224
+        326346.6896203762
+       -174270.6742476623
+        236011.9778065501
+       -239560.8022632156
+        184162.1941532498
+ 2.686e+11   
+         186692.066521993
+       -242855.0440061884
+        330742.4303308096
+        237836.7308724397
+       -321638.7421554076
+        328715.0843291731
+       -175645.2214677031
+        237819.0348721395
+       -241378.3678741402
+        185565.6654998758
+ 2.691e+11   
+        188108.6593609001
+       -244690.0217680835
+        333134.7089623204
+        239645.9295110177
+       -323998.8397934386
+        331086.4269298421
+       -177022.0897089539
+        239628.7880852712
+       -243198.5414290244
+        186971.5330284621
+ 2.696e+11   
+        189527.6768916417
+       -246527.6632472702
+        335530.0335927477
+        241457.7902597451
+       -326361.8290734182
+        333460.6967270378
+        -178401.257386744
+        241441.2146909034
+       -245021.3032326883
+        188379.7753459496
+ 2.701e+11   
+        190949.0978402139
+        -248367.950048805
+        337928.3834074746
+        243272.2904127701
+       -328727.6909462535
+        335837.8728472636
+        -179782.703337127
+        243256.2920042619
+       -246846.6348128015
+        189790.3711699579
+ 2.706e+11   
+         192372.901046789
+       -250210.8649729109
+        340329.7374000587
+        245089.4073496614
+       -331096.4068879052
+        338217.9342647855
+       -181166.4068047315
+        245073.9974129483
+       -248674.5188848928
+        191203.2993257423
+ 2.711e+11   
+           193799.0654619
+       -252056.3919733346
+        342734.0743994911
+        246909.1185370032
+       -333467.9589017085
+        340600.8598281982
+       -182552.3474282793
+        246894.3083785723
+       -250504.9393110067
+        192618.5387423886
+ 2.716e+11   
+        195227.5701418679
+       -253904.5161094728
+        345141.3730981724
+        248731.4015294443
+       -335842.3295177835
+        342986.6282874975
+       -183940.5052238526
+        248717.2024379188
+       -252337.8810521849
+         194036.068448302
+ 2.721e+11   
+        196658.3942435316
+       -255755.2234924625
+        347551.6120804563
+        250556.2339702164
+       -338219.5017894536
+        345375.2183215027
+        -185330.860566003
+        250542.6572036659
+       -254173.3301149594
+        195455.8675660488
+ 2.726e+11   
+        198091.5170183484
+       -257608.5012254387
+        349964.7698516257
+        252383.5935911481
+       -340599.4592866095
+        347766.6085654923
+       -186723.3941668035
+        252370.6503646864
+       -256011.2734920629
+        196877.9153066228
+ 2.731e+11   
+        199526.9178059419
+         -259464.33733817
+        352380.8248671567
+         254213.458212205
+       -342982.1860859558
+        350160.7776389151
+        -188118.087052949
+        254201.1596859558
+       -257851.6990975621
+        198302.1909632071
+ 2.736e+11   
+        200964.5760271777
+       -261322.7207162975
+        354799.7555621492
+        256045.8057405934
+       -345367.6667580869
+        352557.7041730462
+       -189514.9205410218
+        256034.1630081138
+        -259694.595696638
+        199728.6739045182
+ 2.741e+11   
+        202404.4711768542
+       -263183.6410254003
+        357221.5403807863
+        257880.6141694658
+       -347755.8863513435
+        354957.3668384604
+       -190913.8762110394
+        257869.6382467121
+       -261539.9528302354
+        201157.3435678135
+ 2.746e+11   
+        203846.5828161027
+       -265047.0886301335
+         359646.157805721
+        259717.8615762851
+       -350146.8303724176
+        357359.7443722144
+       -192314.9358784136
+        259707.5633912061
+       -263387.7607348174
+        202588.1794516588
+ 2.751e+11   
+        205290.8905645916
+        -266913.054508671
+        362073.5863872588
+        261557.5261208869
+       -352540.4847636602
+        359764.8156046087
+       -193718.0815644494
+        261547.9165037361
+       -265238.0102574662
+        204021.1611085516
+ 2.756e+11   
+        206737.3740926434
+        -268781.530162708
+        364503.8047722421
+        263399.5860433101
+        -354936.835877078
+        362172.5594854376
+       -195123.2954655222
+        263390.6757177609
+       -267090.6927665701
+        205456.2681375014
+ 2.761e+11   
+        208186.0131133631
+        -270652.507523271
+        366936.7917325258
+         265244.019661449
+       -357335.8704449892
+        364582.9551096185
+       -196530.5599210711
+        265235.8192366009
+       -268945.8000583508
+        206893.4801766752
+ 2.766e+11   
+        209636.7873748972
+       -272525.9788525893
+        369372.5261929477
+        267090.8053685939
+       -359737.5755473239
+        366995.9817421016
+       -197939.8573805526
+        267083.3253319577
+       -270803.3242594743
+        208332.7768962132
+ 2.771e+11   
+        211089.6766529312
+       -274401.9366422885
+        371810.9872587071
+        268939.9216309306
+        -362141.938575562
+        369411.6188419775
+       -199351.1703695037
+        268933.1723424807
+       -272663.2577260119
+        209774.1379913356
+ 2.776e+11   
+        212544.6607435466
+       -276280.3735081655
+        374252.1542420622
+        270791.3469850708
+       -364548.9471933026
+        371829.8460856911
+       -200764.4814548623
+        270785.3386724496
+       -274525.5929389942
+        211217.5431758483
+ 2.781e+11   
+        214001.7194565572
+       -278161.2820818002
+        376696.0066882598
+        272645.0600356875
+       -366958.5892934622
+        374250.6433892866
+       -202179.7732096983
+        272639.8027906495
+       -276390.3223968256
+        212662.9721761721
+ 2.786e+11   
+        215460.8326094447
+       -280044.6548992699
+        379142.5244006299
+        274501.0394533332
+       -369370.8529521084
+        376673.9909296027
+       -203597.0281775104
+         274496.543229516
+       -278257.4385048109
+        214110.4047260145
+ 2.791e+11   
+        216921.9800220229
+       -281930.4842872267
+        381591.6874647664
+        276359.2639725219
+       -371785.7263789363
+        379099.8691643547
+       -205016.2288362439
+        276355.5385846281
+       -280126.9334620541
+        215559.8205618072
+ 2.796e+11   
+        218385.1415119519
+       -283818.7622465977
+        384043.4762717334
+        278219.7123901592
+       -374203.1978644052
+        381528.2588510372
+       -206437.3575621891
+        278216.7675146335
+       -281998.7991459875
+        217011.1994190345
+ 2.801e+11   
+        219850.2968912352
+       -285709.4803341639
+        386497.8715402262
+        280082.3635643991
+       -376623.2557235433
+        383959.1410645818
+       -207860.3965939168
+        280080.2087416883
+       -283873.0269947829
+        218464.5210295789
+ 2.806e+11   
+        221317.4259638235
+       -287602.6295422808
+        388954.8543376386
+        281947.1964140201
+       -379045.8882364492
+        386392.4972137216
+       -209285.3279964123
+        281945.8410524948
+       -285749.6078879048
+         219919.765120212
+ 2.811e+11   
+        222786.5085244614
+       -289498.2001769936
+        391414.4060999766
+         283814.189918403
+       -381471.0835855117
+        388828.3090560065
+       -210712.1336255669
+        283813.6433000272
+       -287628.5320250535
+        221376.9114123578
+ 2.816e+11   
+        224257.5243589024
+       -291396.1817347996
+        393876.5086505751
+        285683.3231182019
+       -383898.8297893735
+        391266.5587114261
+       -212140.7950931872
+        285683.5944060287
+       -289509.7888037484
+        222835.9396232566
+ 2.821e+11   
+        225730.4532456247
+       -293296.5627783068
+        396341.1442175625
+        287554.5751167956
+       -386329.1146336708
+         393707.228674593
+       -213571.2937326828
+         287555.673364372
+       -291393.3666958033
+        224296.8294686627
+ 2.826e+11   
+        227205.2749591821
+       -295199.3308110409
+        398808.2954500476
+        289427.9250826108
+       -388761.9255985811
+        396150.3018254532
+       -215003.6105655919
+        289429.8592453698
+       -293279.2531229305
+        225759.5606672003
+ 2.831e+11   
+        228681.9692753177
+       -297104.4721516388
+        401277.9454329782
+        291303.3522524094
+       -391197.2497832199
+        398595.7614384866
+       -216437.7262691033
+        291306.1312011266
+       -295167.4343317201
+        227224.1129465105
+ 2.836e+11   
+        230160.5159779729
+       -299011.9718076728
+        403750.0777006446
+        293180.8359356267
+       -393635.0738269158
+        401043.5911903667
+       -217873.6211447364
+        293184.4684720206
+       -297057.8952682306
+        228690.4660513169
+ 2.841e+11   
+        231640.8948683218
+       -300921.8133493389
+        406224.6762488008
+        295060.3555198587
+       -396075.3838274182
+        403493.7751660561
+       -219311.2750883338
+        295064.8503944095
+       -298950.6194524224
+        230158.5997535412
+ 2.846e+11   
+        233123.0857759664
+       -302833.9787832453
+        408701.7255453721
+        296941.8904775862
+       -398518.1652560713
+        405946.2978633127
+        -220750.667561525
+        296947.2564096435
+       -300845.5888526646
+        231628.4938645917
+ 2.851e+11   
+        234607.0685724127
+        -304748.448426526
+        411181.2105397333
+        298825.4203742283
+       -400963.4028700066
+        408401.1441955882
+       -222191.7775648203
+        298831.6660744885
+       -302742.7837605439
+        233100.1282499617
+ 2.856e+11   
+        236092.8231869659
+       -306665.2007815035
+        413663.1166705351
+        300710.9248776205
+       -403411.0806214023
+        410858.2994933047
+       -223634.5836124838
+        300718.0590730373
+       -304642.1826661914
+        234573.4828462545
+ 2.861e+11   
+        237580.3296251711
+       -308584.2124111278
+        416147.4298720698
+        302598.3837690061
+       -405861.1815638588
+        413317.7495034986
+       -225079.0637093472
+        302606.4152302121
+       -306543.7621343508
+        236048.5376807713
+ 2.866e+11   
+        239069.5679899218
+       -310505.4578153955
+        418634.1365791595
+        304487.7769556384
+        -408313.687755949
+        415779.4803878216
+       -226525.1953297102
+        304496.7145269378
+       -308447.4966813941
+        237525.2728937787
+ 2.871e+11   
+        240560.5185053732
+       -312428.9093089728
+        421123.2237305661
+        306379.0844850833
+       -410768.5801619965
+         418243.478718902
+       -227972.9553984867
+        306388.9371170905
+       -310353.3586535047
+        239003.6687635909
+ 2.876e+11   
+        242053.1615437751
+       -314354.5369002208
+        423614.6787709151
+        308272.2865613135
+       -413225.8385501383
+        420709.7314750553
+        -229422.320274741
+        308283.0633462999
+         -312261.31810622
+        240483.7057345793
+ 2.881e+11   
+        243547.4776553593
+       -316282.3081718312
+         426108.489651138
+        310167.3635626941
+       -415685.4413877411
+        423178.2260333596
+         -230873.26573777
+        310179.0737727071
+       -314171.3426855454
+        241965.3644482437
+ 2.886e+11   
+        245043.4476014013
+       -318212.1881632737
+        428604.6448274383
+        312064.2960619481
+       -418147.3657342305
+        425648.9501610998
+       -232325.7669758767
+        312076.9491897644
+        -316083.397510832
+        243448.6257774597
+ 2.891e+11   
+        246541.0523905791
+       -320144.1392552428
+        431103.1332587842
+        313963.0648481932
+       -420611.5871313955
+        428121.8920055854
+       -233779.7985779855
+        313976.6706511705
+       -317997.4450596113
+        244933.4708640288
+ 2.896e+11   
+         248040.273318756
+       -322078.1210563053
+        433603.9444029477
+        315863.6509511531
+       -423078.0794912488
+         430597.040082371
+       -235235.3345282465
+        315878.2194980358
+       -319913.4450545799
+        246419.8811596508
+ 2.901e+11   
+        249541.0920123086
+       -324014.0902919326
+        436107.0682111059
+        317766.0356676291
+       -425546.8149815072
+        433074.3832618909
+       -236692.3482037761
+        317781.5773883679
+       -321831.3543529168
+        247907.8384704389
+ 2.906e+11   
+        251043.4904751189
+       -325952.0006961009
+        438612.4951210205
+        319670.2005903318
+       -428017.7639087698
+        435553.9107545334
+       -238150.8123756798
+        319686.7263289728
+       -323751.1268381203
+        249397.3250050983
+ 2.911e+11   
+        252547.4511393566
+       -327891.8029056464
+        441120.2160488285
+        321576.1276391686
+       -430490.8945994747
+        438035.6120941878
+       -239610.6992135066
+        321593.6487098671
+       -325672.7133145423
+        250888.3234268876
+ 2.916e+11   
+        254052.9569201679
+       -329833.4443575496
+        443630.2223794677
+        323483.7990950827
+       -432966.1732787124
+        440519.4771202912
+       -241071.9802932755
+        323502.3273412932
+        -327596.061404797
+        252380.8169094809
+ 2.921e+11   
+        255559.9912743942
+       -331776.8691893262
+        446142.5059557763
+        325393.1976365409
+       -435443.5639469844
+        443005.4959584184
+       -242534.6266092247
+         325412.745493436
+       -329521.1154502184
+        253874.7891968494
+ 2.926e+11   
+         257068.538263438
+       -333722.0181426975
+        448657.0590662998
+        327304.3063787692
+       -437923.0282549937
+        445493.6589994525
+       -243998.6085894248
+        327324.8869389363
+       -331447.8164145386
+        255370.2246672809
+ 2.931e+11   
+         258578.582620394
+        -335668.828470709
+         451173.874431852
+        329217.1089158333
+       -440404.5253765567
+        447983.9568773849
+       -245463.8961154023
+        329238.7359982971
+       -333376.1017909534
+        256867.1084016527
+ 2.936e+11   
+        260090.1098215605
+       -337617.2338484602
+        453692.9451908723
+        331131.5893656603
+       -442888.0118797324
+        450476.3804457897
+       -246930.4585459115
+        331154.2775882778
+        -335305.905512738
+          258365.42625607
+ 2.941e+11   
+        261603.1061624523
+       -339567.1642876146
+        456214.2648836328
+        333047.7324181027
+        -445373.441596261
+        452970.9207530289
+       -248398.2647450004
+        333071.4972733745
+       -337237.1578675759
+        259865.1649389884
+ 2.946e+11   
+        263117.5588384138
+       -341518.5460548328
+        458737.8274353343
+        334965.5233861335
+       -447860.7654894106
+        455467.5690162392
+       -249867.2831145019
+        334990.3813204771
+       -339169.7854157548
+        261366.3120929241
+ 2.951e+11   
+         264633.456029953
+        -343471.301594296
+        461263.6271381621
+        336884.9482602727
+       -450349.9315203272
+        457966.3165941577
+       -251337.4816310848
+        336910.9167567936
+       -341103.7109123758
+        262868.8563808599
+ 2.956e+11   
+        266150.7869928853
+       -345425.3494544464
+        463791.6586323304
+        338805.9937663228
+       -452840.8845129798
+        460467.1549588373
+       -252808.8278879894
+        338833.0914311301
+       -343038.8532337231
+        264372.7875774481
+ 2.961e+11   
+          267669.54215339
+       -347380.6042190862
+        466321.9168861791
+         340728.647426502
+        -455333.566017797
+        462970.0756663058
+       -254281.2891415609
+        340756.8940786014
+       -344975.1273079196
+        265878.0966650961
+ 2.966e+11   
+        269189.7132080533
+       -349336.9764429521
+        468854.3971753537
+         342652.897624039
+       -457827.9141740682
+        465475.0703262117
+       -255754.8323626841
+        342682.3143888412
+       -346912.4440499894
+         267384.775935022
+ 2.971e+11   
+        270711.2932289679
+       -351294.3725918633
+        471389.0950611045
+        344578.7336712853
+       -460323.8635711879
+        467982.1305704867
+       -257229.4242932023
+        344609.3430777656
+       -348850.7103014282
+        268892.8190933392
+ 2.976e+11   
+        272234.2767739394
+       -353252.6949875344
+        473926.0063677226
+        346506.1458813862
+       -462821.3451088039
+        470491.2480210579
+        -258705.031507383
+        346537.9719629263
+       -350789.8287743633
+        270402.2213722224
+ 2.981e+11   
+        273758.6600018177
+       -355211.8417570885
+        476465.1271590972
+        348435.1256435104
+       -465320.2858558887
+        473002.4142565886
+       -260181.6204784571
+        348468.1940424559
+       -352729.6980003502
+        271912.9796461712
+ 2.986e+11   
+        275284.4407929453
+       -357171.7067873068
+        479006.4537143772
+        350365.6655016272
+       -467820.6089087575
+        475515.6207782369
+       -261659.1576502247
+        350400.0035775874
+       -354670.2122838278
+        273425.0925533638
+ 2.991e+11   
+        276811.6188746771
+        -359132.179683572
+        481549.9825026496
+         352297.759236757
+       -470322.2332479862
+        478030.8589743526
+       -263137.6095136722
+        352333.3961786801
+       -356611.2616602057
+        274938.5606220526
+ 2.996e+11   
+        278340.1959518623
+       -361093.1457334332
+        484095.7101565285
+          354231.40195258
+       -472825.0735941557
+        480548.1200840023
+       -264616.9426884708
+        354268.3688946216
+       -358552.7318584906
+        276453.3864018922
* NOTE: Solution at 1e+08 Hz used as DC point.
* NOTE: Repaired negative diagonal entries at these frequencies:
*  2e+10 Hz, 2.1e+10 Hz, 2.1e+10 Hz

.model l_m4lines_veryHighFreq_W_1 sp N=4 SPACING=nonuniform VALTYPE=real
+ INTERPOLATION=spline
+ INFINITY =
+     1.24059880231526e-05
+   -1.528022937622716e-05
+     2.24060214148671e-05
+      1.5191092713225e-05
+   -2.097553049136751e-05
+    2.232836754302833e-05
+   -1.088364074586691e-05
+    1.518777564363861e-05
+    -1.52218532717874e-05
+    1.236102136755522e-05
+ DATA = 600
+ 0           
+     4.20266069931064e-07
+     1.49892505860857e-07
+    4.170768222841771e-07
+    4.555134050645788e-08
+     9.33939986199654e-08
+    4.170888506778619e-07
+    2.471028786369816e-08
+    4.556334226522421e-08
+      1.4993074974344e-07
+    4.202232793369385e-07
+ 6e+08       
+    4.137728548351578e-07
+    1.492708365372005e-07
+    4.104530110976688e-07
+     4.52905365811054e-08
+     9.25207309980272e-08
+     4.10472762753663e-07
+    2.461315040040524e-08
+    4.530446051117568e-08
+    1.493103845007641e-07
+    4.137069439857984e-07
+ 1.1e+09     
+    4.126244509636713e-07
+    1.492173472978974e-07
+    4.092758395422161e-07
+    4.524248514961317e-08
+    9.238747072701994e-08
+    4.092976176969652e-07
+    2.459662301950652e-08
+    4.525665291771942e-08
+    1.492564261725866e-07
+    4.125521743247561e-07
+ 1.6e+09     
+    4.121750728235947e-07
+    1.492709864442246e-07
+     4.08800328950587e-07
+    4.519612391949503e-08
+    9.235320059979149e-08
+    4.088232304346868e-07
+    2.456910508441308e-08
+    4.521044478206623e-08
+    1.493098591877597e-07
+    4.120988884779976e-07
+ 2.1e+09     
+    4.117776864397868e-07
+    1.492446039238189e-07
+    4.083876531910376e-07
+    4.518032054575695e-08
+    9.230697865427897e-08
+    4.084110328715542e-07
+    2.455797025243276e-08
+    4.519486841510102e-08
+    1.492832639661574e-07
+    4.116991604201628e-07
+ 2.6e+09     
+    4.114730702905467e-07
+    1.492122763326093e-07
+    4.080769108938253e-07
+    4.519174658367004e-08
+    9.227809755200503e-08
+    4.081003184866233e-07
+    2.456926817988529e-08
+    4.520648936955566e-08
+    1.492507536817829e-07
+    4.113933687193145e-07
+ 3.1e+09     
+     4.11259854088199e-07
+    1.492002449354272e-07
+    4.078623258588693e-07
+    4.522736172053641e-08
+    9.227351546494369e-08
+    4.078855220655792e-07
+    2.460396312584708e-08
+     4.52422694626706e-08
+    1.492385657162871e-07
+    4.111796244189016e-07
+ 3.6e+09     
+    4.111248971147498e-07
+    1.492166256017472e-07
+    4.077279506952679e-07
+    4.528510629361827e-08
+    9.229539577144972e-08
+    4.077508318609027e-07
+    2.466101083036246e-08
+    4.530015927770827e-08
+    1.492548093126842e-07
+    4.110444438160116e-07
+ 4.1e+09     
+    4.110547112432908e-07
+    1.492634686531503e-07
+    4.076592347367265e-07
+     4.53639540736727e-08
+     9.23461924290262e-08
+    4.076817683576236e-07
+    2.473893597314369e-08
+    4.537914078847674e-08
+    1.493015329828699e-07
+    4.109741586994824e-07
+ 4.6e+09     
+    4.110383566212247e-07
+    1.493408556734908e-07
+    4.076451817146062e-07
+    4.546358571847223e-08
+    9.242893832980684e-08
+    4.076673681602417e-07
+    2.483640212235767e-08
+    4.547890054393931e-08
+    1.493788201734081e-07
+    4.109577479229974e-07
+ 5.1e+09     
+    4.110675278814131e-07
+    1.494480676961413e-07
+    4.076774911265828e-07
+    4.558370933650535e-08
+    9.254438922828138e-08
+    4.076993437325702e-07
+    2.495229175713058e-08
+    4.559915058902342e-08
+    1.494859547590938e-07
+    4.109868757557435e-07
+ 5.6e+09     
+    4.111359702603132e-07
+    1.495837978424644e-07
+    4.077492659026733e-07
+    4.572345620906127e-08
+     9.26881657256158e-08
+    4.077708008677062e-07
+    2.508563524448641e-08
+    4.573902444661221e-08
+    1.496216304991523e-07
+    4.110552802845713e-07
+ 6.1e+09     
+    4.112389082592219e-07
+    1.497462580623919e-07
+    4.078546868192754e-07
+    4.588162033293626e-08
+    9.285297756863277e-08
+    4.078759174305414e-07
+    2.523562625083437e-08
+    4.589731701148803e-08
+    1.497840541598155e-07
+    4.111581873309013e-07
+ 6.6e+09     
+    4.113726198218682e-07
+    1.499333297512874e-07
+    4.079894036172784e-07
+    4.605741308108181e-08
+     9.30339905123391e-08
+    4.080103361318821e-07
+    2.540171434973479e-08
+    4.607323974713961e-08
+    1.499710931707929e-07
+    4.112918772319126e-07
+ 7.1e+09     
+    4.115341210643493e-07
+    1.501426134952328e-07
+    4.081504760569297e-07
+    4.625065729538214e-08
+    9.323055741259585e-08
+    4.081711070585963e-07
+    2.558362044399649e-08
+    4.626661552465196e-08
+    1.501803264599115e-07
+    4.114533670146062e-07
+ 7.6e+09     
+    4.117209805059166e-07
+    1.503715454529629e-07
+    4.083358621144828e-07
+    4.646142913087039e-08
+    9.344427627502937e-08
+    4.083561793699695e-07
+    2.578128729750871e-08
+    4.647752148862196e-08
+    1.504091707749235e-07
+     4.11640226500467e-07
+ 8.1e+09     
+    4.119313107402051e-07
+    1.506178729278335e-07
+    4.085440846433313e-07
+    4.668975017673128e-08
+    9.367703737060978e-08
+    4.085640738052813e-07
+    2.599486875115079e-08
+      4.6705981694101e-08
+    1.506553747796244e-07
+     4.11850575237082e-07
+ 8.6e+09     
+    4.121639016742112e-07
+    1.508804503011236e-07
+    4.087742342345746e-07
+    4.693554647524229e-08
+    9.393028317402522e-08
+    4.087938898227176e-07
+    2.622478970475343e-08
+    4.695192315610689e-08
+    1.509178280971092e-07
+    4.120832195639344e-07
+ 9.1e+09     
+    4.124183431962331e-07
+    1.511598921000274e-07
+    4.090260793771636e-07
+    4.719882139975483e-08
+    9.420499917507315e-08
+     4.09045412396398e-07
+    2.647185187309692e-08
+    4.721533698758624e-08
+    1.511972008794427e-07
+    4.123377708003081e-07
+ 9.6e+09     
+     4.12694966780804e-07
+    1.514585417711409e-07
+    4.093000350167233e-07
+    4.748001503522429e-08
+    9.450193445547068e-08
+    4.093190699961506e-07
+    2.673736321921395e-08
+    4.749661214563698e-08
+    1.514958728352864e-07
+    4.126145738455468e-07
+ 1.01e+10    
+    4.129796793319785e-07
+    1.517557829651655e-07
+    4.095849853130342e-07
+     4.77472106636134e-08
+    9.479328297952915e-08
+    4.096037851608875e-07
+    2.699310527978731e-08
+    4.776384162367628e-08
+    1.517931397096729e-07
+    4.128989981582042e-07
+ 1.06e+10    
+    4.132194239673054e-07
+    1.519718564017253e-07
+    4.098350610067127e-07
+     4.78922514101228e-08
+    9.498365903173492e-08
+    4.098537624640855e-07
+    2.713968926344471e-08
+    4.790937733487321e-08
+    1.520089864090429e-07
+    4.131365315724783e-07
+ 1.11e+10    
+    4.134676443349587e-07
+    1.521955757680202e-07
+    4.100907212704122e-07
+    4.804225703475203e-08
+     9.51804717456942e-08
+    4.101092989848254e-07
+    2.729079797685548e-08
+    4.805992587708687e-08
+    1.522325074113614e-07
+    4.133828304428554e-07
+ 1.16e+10    
+     4.13724007883129e-07
+    1.524266673096013e-07
+    4.103515694318296e-07
+    4.819698847643358e-08
+    9.538344621185501e-08
+    4.103699986769501e-07
+    2.744611956320201e-08
+    4.821524955678689e-08
+    1.524634269619907e-07
+    4.136375431402382e-07
+ 1.21e+10    
+    4.139881997283174e-07
+    1.526648641915497e-07
+    4.106172489955454e-07
+     4.83562048787339e-08
+    9.559231162714905e-08
+    4.106355058732364e-07
+    2.760533866458407e-08
+    4.837510906878737e-08
+     1.52701476235551e-07
+    4.139003352632263e-07
+ 1.26e+10    
+    4.142599240139137e-07
+    1.529099070769148e-07
+    4.108874416355019e-07
+    4.851966425973665e-08
+    9.580680179798677e-08
+    4.109055032313605e-07
+    2.776813745055491e-08
+    4.853926420183159e-08
+    1.529463939686722e-07
+    4.141708915298451e-07
+ 1.31e+10    
+    4.145389046642303e-07
+    1.531615445477268e-07
+    4.111618648793102e-07
+    4.868712415960734e-08
+    9.602665556677851e-08
+    4.111797093748673e-07
+     2.79341966062811e-08
+    4.870747451782353e-08
+    1.531979269192175e-07
+    4.144489169177014e-07
+ 1.36e+10    
+    4.148248856294526e-07
+    1.534195333919273e-07
+    4.114402695966584e-07
+    4.885834227451025e-08
+    9.625161717556637e-08
+    4.114578763424607e-07
+    2.810319628154639e-08
+    4.887950001462722e-08
+    1.534558301790836e-07
+    4.147341371783138e-07
+ 1.41e+10    
+    4.151176307152923e-07
+    1.536836387779657e-07
+    4.117224373874946e-07
+    4.903307708715224e-08
+    9.648143657955484e-08
+    4.117397869413048e-07
+    2.827481700199439e-08
+     4.90551017827941e-08
+     1.53719867364903e-07
+    4.150262988452892e-07
+ 1.46e+10    
+    4.154169230858753e-07
+    1.539536343379867e-07
+     4.12008177947928e-07
+    4.921108850484614e-08
+    9.671586972243304e-08
+    4.120252520830226e-07
+    2.844874054515911e-08
+    4.923404266792206e-08
+    1.539898107102574e-07
+    4.153251688463357e-07
+ 1.51e+10    
+    4.157225645198781e-07
+    1.542293021779598e-07
+    4.122973264768756e-07
+    4.939213851827846e-08
+    9.695467878395744e-08
+    4.123141081643832e-07
+    2.862465078441895e-08
+    4.941608795122206e-08
+    1.542654410795141e-07
+    4.156305338165706e-07
+ 1.56e+10    
+    4.160343744906794e-07
+    1.545104328322629e-07
+    4.125897411717913e-07
+    4.957599189573867e-08
+    9.719763241062198e-08
+    4.126062145420858e-07
+    2.880223450509514e-08
+    4.960100606319004e-08
+    1.545465479220423e-07
+    4.159421991974217e-07
+ 1.61e+10    
+    4.163521891312149e-07
+     1.54796825177589e-07
+    4.128853008504264e-07
+    4.976241693133493e-08
+    9.744450593943338e-08
+    4.129014511371393e-07
+    2.898118219792492e-08
+    4.978856934737403e-08
+    1.548329291832365e-07
+    4.162599881927955e-07
+ 1.66e+10    
+    4.166758601348033e-07
+     1.55088286320399e-07
+    4.131839027244589e-07
+    4.995118626837062e-08
+    9.769508162535434e-08
+    4.131997161950483e-07
+    2.916118883654017e-08
+    4.997855489454066e-08
+    1.551243911868426e-07
+    4.165837406416315e-07
+ 1.71e+10    
+     4.17005253634193e-07
+    1.553846314702391e-07
+    4.134854603431672e-07
+    5.014207782547063e-08
+     9.79491488840389e-08
+    4.135009242194428e-07
+     2.93419546472041e-08
+    5.017074547206224e-08
+    1.554207485017135e-07
+    4.169133118553564e-07
+ 1.76e+10    
+    4.173402490935231e-07
+    1.556856838111533e-07
+    4.137899017181977e-07
+    5.033487585881771e-08
+    9.820650456260725e-08
+    4.138050040899237e-07
+    2.952318588151522e-08
+    5.036493057857422e-08
+    1.557218238053724e-07
+    4.172485714593998e-07
+ 1.81e+10    
+    4.176807382411174e-07
+    1.559912743825573e-07
+    4.140971676358291e-07
+    5.052937220250792e-08
+    9.846695325327196e-08
+       4.141118973706e-07
+    2.970459560518556e-08
+    5.056090766134304e-08
+    1.560274477556069e-07
+    4.175894022696052e-07
+ 1.86e+10    
+    4.180266240655242e-07
+    1.563012419812093e-07
+    4.144072101599715e-07
+    5.072536774072187e-08
+    9.873030766804057e-08
+    4.144215568119243e-07
+    2.988590451951843e-08
+    5.075848354304327e-08
+     1.56337458881725e-07
+    4.179356992283704e-07
+ 1.91e+10    
+    4.183778198934137e-07
+    1.566154330966346e-07
+    4.147199913265833e-07
+    5.092267417884189e-08
+    9.899638909613239e-08
+    4.147339450473249e-07
+    3.006684183691327e-08
+    5.095747611610573e-08
+    1.566517035072486e-07
+    4.182873684199543e-07
+ 1.96e+10    
+    4.187342485649662e-07
+    1.569337018938688e-07
+    4.150354820300797e-07
+    5.112111619999071e-08
+    9.926502797126568e-08
+      4.1504903348482e-07
+    3.024714623672492e-08
+    5.115771637776238e-08
+    1.569700357168956e-07
+    4.186443261811777e-07
+ 2.01e+10    
+    4.190958417207158e-07
+     1.57255910259099e-07
+    4.153536611028324e-07
+    5.132053411635391e-08
+     9.95360645827425e-08
+    4.153668013957689e-07
+    3.042656693532243e-08
+    5.135905089787513e-08
+    1.572923173824346e-07
+    4.190064983209898e-07
+ 2.06e+10    
+    4.194625392138004e-07
+    1.575819279272544e-07
+     4.15674514590152e-07
+    5.152078715531734e-08
+    9.980934997290188e-08
+    4.156872352037771e-07
+    3.060486491264086e-08
+    5.156134483487133e-08
+    1.576184182646321e-07
+    4.193738194617639e-07
+ 2.11e+10    
+    4.198342886624895e-07
+    1.579116327145394e-07
+    4.159980352269673e-07
+    5.172175755905826e-08
+    1.000847470743669e-07
+    4.160103279812795e-07
+    3.078181434923299e-08
+    5.176448564521934e-08
+    1.579482162118274e-07
+     4.19746232515159e-07
+ 2.16e+10    
+     4.20211045160431e-07
+    1.582449108844495e-07
+    4.163242221258927e-07
+    5.192335572493467e-08
+    1.003621321550965e-07
+    4.163360791659629e-07
+    3.095720434122414e-08
+    5.196838766807403e-08
+    1.582815974802657e-07
+    4.201236883068651e-07
+ 2.21e+10    
+    4.205927711661375e-07
+    1.585816576829267e-07
+    4.166530806923273e-07
+     5.21255266761102e-08
+    1.006413966558182e-07
+    4.166644945149012e-07
+    3.113084097888418e-08
+    5.217299781238466e-08
+    1.586184572074408e-07
+    4.205061453673138e-07
+ 2.26e+10    
+    4.209794365986892e-07
+    1.589217780873601e-07
+    4.169846227895384e-07
+    5.232825822820238e-08
+    1.009224495270723e-07
+    4.169955863236226e-07
+    3.130254989537944e-08
+    5.237830262800271e-08
+    1.589587000766114e-07
+    4.208935699093472e-07
+ 2.31e+10    
+     4.21371019174579e-07
+    1.592651878251177e-07
+     4.17318867184596e-07
+     5.25315913111887e-08
+    1.012052201982302e-07
+    4.173293739464556e-07
+    3.147217941853403e-08
+    5.258433710675084e-08
+    1.593022412199842e-07
+    4.212859360191254e-07
+ 2.36e+10    
+    4.217675050292189e-07
+    1.596118147304979e-07
+    4.176558403164258e-07
+    5.273563301640488e-08
+    1.014896623416282e-07
+    4.176658846663153e-07
+    3.163960448905445e-08
+     5.27911956316911e-08
+    1.596490074178741e-07
+    4.216832260927658e-07
+ 2.41e+10    
+    4.221688896779257e-07
+    1.599616005238287e-07
+    4.179955774378934e-07
+    5.294057306274836e-08
+    1.017757586285858e-07
+    4.180051549761028e-07
+    3.180473154129198e-08
+    5.299904557008362e-08
+    1.599989386631241e-07
+    4.220854315585079e-07
+ 2.46e+10    
+    4.225751793823257e-07
+     1.60314503112203e-07
+    4.183381241949921e-07
+    5.314670450358735e-08
+     1.02063526707406e-07
+    4.183472323467395e-07
+    3.196750457692533e-08
+    5.320814407491702e-08
+    1.603519901703584e-07
+    4.224925539310635e-07
+ 2.51e+10    
+    4.229863929984741e-07
+    1.606704995239022e-07
+    4.186835387142419e-07
+     5.33544496025201e-08
+    1.023530266599169e-07
+    4.186921775695953e-07
+    3.212791268744915e-08
+    5.341885870337351e-08
+    1.607081349186406e-07
+    4.229046062500027e-07
+ 2.56e+10    
+    4.234025643879747e-07
+    1.610295895940663e-07
+    4.190318942722184e-07
+    5.356439184211557e-08
+    1.026443701979766e-07
+    4.190400677655481e-07
+    3.228599928696617e-08
+    5.363169243726604e-08
+    1.610673668157664e-07
+    4.233216149544546e-07
+ 2.61e+10    
+    4.238237454658075e-07
+    1.613918005049485e-07
+    4.193832826079345e-07
+    5.377731490208892e-08
+    1.029377318189894e-07
+    4.193910001433745e-07
+     3.24418732744612e-08
+    5.384731353259105e-08
+    1.614297045563064e-07
+    4.237436222353339e-07
+ 2.66e+10    
+     4.24250009924995e-07
+    1.617571922320584e-07
+    4.197378178996007e-07
+    5.399424898699698e-08
+    1.032333620042165e-07
+    4.197450965479294e-07
+    3.259572221051933e-08
+      5.4066590217284e-08
+    1.617951961963308e-07
+    4.241706888757335e-07
+ 2.71e+10    
+    4.246814575953174e-07
+    1.621258638242852e-07
+    4.200956413357987e-07
+    5.421652381753518e-08
+    1.035316022399215e-07
+    4.201025087385018e-07
+    3.274782729243605e-08
+    5.429062941111237e-08
+    1.621639243598506e-07
+    4.246028975212745e-07
+ 2.76e+10    
+    4.251182192249768e-07
+    1.624979602001355e-07
+    4.204569260358989e-07
+    5.444582547561093e-08
+    1.038329010491991e-07
+    4.204634241363738e-07
+    3.289857932279412e-08
+    5.452081707566246e-08
+    1.625360117866976e-07
+    4.250403561929127e-07
+ 2.81e+10    
+    4.255604611635814e-07
+    1.628736786947655e-07
+    4.208218817611775e-07
+    5.468425045022054e-08
+    1.041378291683715e-07
+     4.20828071413094e-07
+    3.304849382052671e-08
+    5.475885511377815e-08
+     1.62911626568918e-07
+    4.254832016271449e-07
+ 2.86e+10    
+    4.260083889005236e-07
+    1.632532738440946e-07
+    4.211907583436071e-07
+    5.493434380006309e-08
+    1.044470902593187e-07
+    4.211967246746408e-07
+    3.319822169230429e-08
+    5.500678543084731e-08
+    1.632909858308647e-07
+    4.259316016579303e-07
+ 2.91e+10    
+    4.264622475962618e-07
+    1.636370577357886e-07
+    4.215638459750386e-07
+    5.519909846330862e-08
+    1.047615208968959e-07
+     4.21569704042995e-07
+    3.334854924683947e-08
+    5.526698538299203e-08
+    1.636743557132442e-07
+    4.263857552966125e-07
+ 2.96e+10    
+     4.26922316607849e-07
+    1.640253916619143e-07
+    4.219414694291785e-07
+    5.548187916727652e-08
+    1.050820699461121e-07
+    4.219473691155859e-07
+    3.350037773292606e-08
+    5.554211031385201e-08
+    1.640620443047716e-07
+    4.268458884083256e-07
+ 3.01e+10    
+    4.273888936903848e-07
+    1.644186629718517e-07
+    4.223239720557235e-07
+    5.578621899087896e-08
+    1.054097433178917e-07
+    4.223301002545217e-07
+    3.365466848111837e-08
+    5.583494935868002e-08
+    1.644543827771272e-07
+    4.273122420143778e-07
+ 3.06e+10    
+    4.278622635710847e-07
+     1.64817239682158e-07
+    4.227116844533709e-07
+     5.61154259679262e-08
+    1.057454971075116e-07
+     4.22718261513544e-07
+      3.3812336758554e-08
+    5.614815385649319e-08
+    1.648516889409233e-07
+    4.277850495842926e-07
+ 3.11e+10    
+    4.283426461088696e-07
+    1.652213961826965e-07
+    4.231048731054226e-07
+    5.647194558728553e-08
+    1.060900638828712e-07
+    4.231121395825238e-07
+    3.397407919060983e-08
+    5.648380140983255e-08
+    1.652542078991378e-07
+    4.282644999029013e-07
+ 3.16e+10    
+    4.288301231599814e-07
+    1.656312089094603e-07
+    4.235036676005025e-07
+    5.685647542902644e-08
+    1.064437091812221e-07
+    4.235118575716911e-07
+    3.414013180592145e-08
+    5.684278541524454e-08
+    1.656620282821889e-07
+    4.287506843302841e-07
+ 3.21e+10    
+    4.293245524653562e-07
+    1.660464337525616e-07
+    4.239079731024612e-07
+    5.726694228027963e-08
+     1.06805943933329e-07
+    4.239172729596621e-07
+    3.430998422704741e-08
+    5.722408308329525e-08
+    1.660749816672132e-07
+    4.292435327357961e-07
+ 3.26e+10    
+     4.29825491039773e-07
+     1.66466396786899e-07
+     4.24317387576558e-07
+    5.769762318730223e-08
+    1.071752629699324e-07
+    4.243278853366702e-07
+    3.448211968009512e-08
+    5.762405613309806e-08
+    1.664925473355882e-07
+    4.297427512911648e-07
+ 3.31e+10    
+    4.303321638545588e-07
+    1.668899486202335e-07
+    4.247311565931442e-07
+    5.813884558538051e-08
+    1.075490231433385e-07
+    4.247427952767247e-07
+    3.465389361464808e-08
+    5.803604677342999e-08
+     1.66913799700709e-07
+    4.302477849943978e-07
+ 3.36e+10    
+    4.308435139188722e-07
+    1.673155334533096e-07
+    4.251482022644744e-07
+     5.85776892552655e-08
+    1.079235805416139e-07
+    4.251607570809657e-07
+    3.482166967500509e-08
+    5.845057226377877e-08
+    1.673374402724581e-07
+     4.30757831630017e-07
+ 3.41e+10    
+    4.313583459604736e-07
+    1.677413911150681e-07
+    4.255672459619439e-07
+    5.899980484278347e-08
+    1.082947385006465e-07
+    4.255803420678323e-07
+    3.498126447971543e-08
+    5.885630438305699e-08
+     1.67761937315143e-07
+    4.312719238606538e-07
+ 3.46e+10    
+    4.318755320820003e-07
+     1.68165849248902e-07
+    4.259870065680929e-07
+    5.939192691016304e-08
+    1.086584232362141e-07
+    4.260001791901539e-07
+    3.512861867400585e-08
+    5.924172586759901e-08
+    1.681857535204748e-07
+    4.317890705388892e-07
+ 3.51e+10    
+    4.323942102929172e-07
+    1.685876093369657e-07
+    4.264064160254376e-07
+    5.974422423502529e-08
+    1.090113758633635e-07
+    4.264191947530432e-07
+    3.526048445701032e-08
+    5.959701300820572e-08
+    1.686075958685759e-07
+    4.323084184783165e-07
+ 3.56e+10    
+    4.329139056998198e-07
+    1.690059264398579e-07
+    4.268247801467911e-07
+     6.00516529633509e-08
+    1.093516242215083e-07
+    4.268367677753615e-07
+    3.537489451783195e-08
+     5.99155310861539e-08
+    1.690266046278426e-07
+    4.328293818276384e-07
+ 3.61e+10    
+    4.334345428996876e-07
+    1.694206350071211e-07
+    4.272418374971674e-07
+    6.031397670783722e-08
+    1.096786024804409e-07
+    4.272527589913547e-07
+    3.547128112126562e-08
+    6.019448649451973e-08
+    1.694424254876018e-07
+    4.333516997566946e-07
+ 3.66e+10    
+    4.339563682097064e-07
+    1.698320436495295e-07
+    4.276577157160869e-07
+    6.053472545311277e-08
+    1.099929470399207e-07
+    4.276674295325707e-07
+    3.555027356047084e-08
+    6.043465996663452e-08
+    1.698551620344498e-07
+    4.338754158054332e-07
+ 3.71e+10    
+    4.344798292072078e-07
+    1.702407645294364e-07
+    4.280728222366986e-07
+    6.071969114666587e-08
+    1.102961090528048e-07
+    4.280813020934348e-07
+    3.561331332410785e-08
+    6.063949793487126e-08
+    1.702652501034046e-07
+    4.344008023148775e-07
+ 3.76e+10    
+    4.350054573151791e-07
+    1.706475430596147e-07
+    4.284877171386714e-07
+    6.087550952395537e-08
+    1.105899405526593e-07
+    4.284950192168588e-07
+    3.566224292249868e-08
+    6.081397835264413e-08
+     1.70673309378216e-07
+    4.349282651809131e-07
+ 3.81e+10    
+    4.355337797619987e-07
+    1.710531274331001e-07
+    4.289030039084864e-07
+    6.100862756304528e-08
+    1.108763595544688e-07
+    4.289092327273412e-07
+    3.569897308362796e-08
+    6.096359278543807e-08
+    1.710800146236346e-07
+    4.354582578858738e-07
+ 3.86e+10    
+    4.360652671227319e-07
+    1.714581888360424e-07
+    4.293192540623255e-07
+    6.112471147049951e-08
+    1.111571324667829e-07
+    4.293245346695189e-07
+    3.572526644727418e-08
+     6.10936171761265e-08
+    1.714860060398141e-07
+    4.359912194964295e-07
+ 3.91e+10    
+    4.366003105043442e-07
+    1.718632850663462e-07
+    4.297369657383563e-07
+    6.122840984907261e-08
+    1.114337645691639e-07
+    4.297414246132854e-07
+    3.574262860690831e-08
+    6.120869321403619e-08
+     1.71891839475986e-07
+    4.365275386476878e-07
+ 3.96e+10    
+    4.371392184848469e-07
+    1.722688537857904e-07
+    4.301565483793381e-07
+    6.132334649263425e-08
+    1.117074686772246e-07
+    4.301603022646312e-07
+    3.575227683711157e-08
+    6.131265845482548e-08
+    1.722979675552693e-07
+       4.370675384561e-07
+ 4.01e+10    
+     4.37682224831216e-07
+    1.726752224083424e-07
+    4.305783239649116e-07
+     6.14122335288187e-08
+    1.119791805516037e-07
+    4.305814746024742e-07
+    3.575515527725322e-08
+    6.140853979336528e-08
+     1.72704740567808e-07
+      4.3761147527336e-07
+ 4.06e+10    
+    4.382295006544496e-07
+    1.730826251919383e-07
+    4.310025368692364e-07
+    6.149702997161737e-08
+    1.122495966934103e-07
+    4.310051695552466e-07
+    3.575197237447824e-08
+    6.149863552308543e-08
+    1.731124177644948e-07
+    4.381595450361498e-07
+ 4.11e+10    
+    4.387811672365181e-07
+    1.734912217926925e-07
+    4.314293669560734e-07
+    6.157910254715921e-08
+    1.125192188437759e-07
+     4.31431551265788e-07
+    3.574324500377908e-08
+    6.158463337030982e-08
+    1.735211826317588e-07
+    4.387118927908187e-07
+ 4.16e+10    
+     4.39337307651439e-07
+    1.739011143281287e-07
+    4.318589427809822e-07
+    6.165936821495197e-08
+    1.127883965849176e-07
+    4.318607343357209e-07
+    3.572934071451891e-08
+    6.166773298448494e-08
+    1.739311583895521e-07
+    4.392686227231322e-07
+ 4.21e+10    
+     4.39897976471095e-07
+     1.74312361765831e-07
+    4.322913533703693e-07
+    6.173841139109536e-08
+    1.130573641888556e-07
+    4.322927959571803e-07
+    3.571051427211287e-08
+    6.174875689629541e-08
+    1.743424218598145e-07
+    4.398298073208841e-07
+ 4.26e+10    
+    4.404632074767449e-07
+    1.747249914321606e-07
+    4.327266580286743e-07
+    6.181657597248435e-08
+    1.133262706348443e-07
+    4.327277856928742e-07
+    3.568693741931684e-08
+    6.182824374370542e-08
+    1.747550150282586e-07
+    4.403954951202266e-07
+ 4.31e+10    
+    4.410330195866095e-07
+    1.751390079011095e-07
+    4.331648941534634e-07
+    6.189403535193772e-08
+    1.135952031239448e-07
+    4.331657330818816e-07
+    3.565872218197118e-08
+    6.190652298141836e-08
+    1.751689542593745e-07
+    4.409657169460243e-07
+ 4.36e+10    
+    4.416074213080939e-07
+    1.755543996932723e-07
+    4.336060832811076e-07
+    6.197084451764835e-08
+    1.138642050082894e-07
+    4.336066534095668e-07
+    3.562593862889208e-08
+    6.198377286821595e-08
+    1.755842374197884e-07
+     4.41540490778985e-07
+ 4.41e+10    
+    4.421864140250802e-07
+    1.759711442333111e-07
+    4.340502356657002e-07
+    6.204697818060423e-08
+    1.141332891944117e-07
+    4.340505520062986e-07
+    3.558862813768555e-08
+    6.206006446060546e-08
+    1.760008492646173e-07
+    4.421198254656177e-07
+ 4.46e+10    
+    4.427699943929988e-07
+    1.763892114662852e-07
+    4.344973536932215e-07
+    6.212235830590135e-08
+    1.144024480119883e-07
+    4.344974274065354e-07
+    3.554681315046958e-08
+     6.21353944248743e-08
+    1.764187654432419e-07
+    4.427037234986563e-07
+ 4.51e+10    
+    4.433581560639776e-07
+    1.768085664631534e-07
+    4.349474343959536e-07
+    6.219687376035814e-08
+    1.146716603890999e-07
+    4.349472736442855e-07
+    3.550050425489337e-08
+    6.220970917916924e-08
+    1.768379554381362e-07
+    4.432921830730207e-07
+ 4.56e+10    
+    4.439508909162419e-07
+    1.772291712760379e-07
+    4.354004712849742e-07
+    6.227039417286182e-08
+    1.149408970099833e-07
+      4.3540008190477e-07
+    3.544970526145051e-08
+    6.228292245070786e-08
+    1.772583846957333e-07
+    4.438851995891584e-07
+ 4.61e+10    
+    4.445481899202897e-07
+    1.776509862428841e-07
+     4.35856455673199e-07
+    6.234277958988565e-08
+    1.152101239801208e-07
+    4.358558417007034e-07
+    3.539441679883075e-08
+    6.235492790508695e-08
+     1.77680016153268e-07
+    4.444827667408334e-07
+ 4.66e+10    
+    4.451500437410936e-07
+    1.780739708910145e-07
+    4.363153776207879e-07
+    6.241388709936813e-08
+    1.154793053973804e-07
+    4.363145417016453e-07
+    3.533463882255021e-08
+     6.24256081271697e-08
+    1.781028113194958e-07
+    4.450848772937389e-07
+ 4.71e+10    
+    4.457564431496953e-07
+    1.784980845514088e-07
+    4.367772266037533e-07
+    6.248357528423968e-08
+    1.157484051273345e-07
+    4.367761703104194e-07
+    3.527037233365076e-08
+    6.249484092422139e-08
+    1.785267310280102e-07
+    4.456915236362303e-07
+ 4.76e+10    
+    4.463673792979474e-07
+    1.789232867648724e-07
+    4.372419919800941e-07
+    6.255170713189505e-08
+    1.160173880035895e-07
+    4.372407160577033e-07
+    3.520162052642584e-08
+    6.256250367703922e-08
+    1.789517359523484e-07
+    4.463026981628374e-07
+ 4.81e+10    
+    4.469828438955726e-07
+    1.793495375400174e-07
+    4.377096633091157e-07
+    6.261815185342122e-08
+    1.162862206153061e-07
+    4.377081678653922e-07
+    3.512838952581516e-08
+    6.262847627749491e-08
+    1.793777869486099e-07
+     4.46918393536069e-07
+ 4.86e+10    
+    4.476028293179018e-07
+    1.797767975062902e-07
+    4.381802305647194e-07
+    6.268278593859135e-08
+    1.165548717998628e-07
+    4.381785152164743e-07
+    3.505068883287627e-08
+    6.269264304882472e-08
+    1.798048452742262e-07
+     4.47538602860028e-07
+ 4.91e+10    
+    4.482273286650277e-07
+     1.80205027993438e-07
+    4.386536842726018e-07
+    6.274549368140745e-08
+    1.168233129277997e-07
+    4.386517482587948e-07
+     3.49685315631408e-08
+    6.275489393897471e-08
+    1.802328727182777e-07
+    4.481633197904673e-07
+ 4.96e+10    
+    4.488563357869213e-07
+    1.806341910600983e-07
+    4.391300155931823e-07
+    6.280616734347207e-08
+    1.170915180412621e-07
+    4.391278578618788e-07
+    3.488193453989845e-08
+    6.281512519912019e-08
+    1.806618316693962e-07
+    4.487925385994441e-07
+ 5.01e+10    
+    4.494898452854083e-07
+    1.810642494874987e-07
+     4.39609216366251e-07
+    6.286470707455188e-08
+    1.173594638920059e-07
+    4.396068356414856e-07
+     3.47909182876818e-08
+    6.287323970105194e-08
+    1.810916851398894e-07
+    4.494262542077664e-07
+ 5.06e+10    
+    4.501278525004327e-07
+    1.814951667501698e-07
+    4.400912791287317e-07
+    6.292102067510792e-08
+    1.176271299108226e-07
+    4.400886739620526e-07
+    3.469550695744308e-08
+    6.292914700539646e-08
+    1.815223967600203e-07
+    4.500644621949101e-07
+ 5.11e+10    
+    4.507703534861982e-07
+    1.819269069719144e-07
+     4.40576197114246e-07
+    6.297502326020697e-08
+    1.178944981318597e-07
+    4.405733659239917e-07
+    3.459572820685534e-08
+     6.29827632609132e-08
+    1.819539307520385e-07
+    4.507071587933762e-07
+ 5.16e+10    
+     4.51417344980918e-07
+    1.823594348726874e-07
+    4.410639642400365e-07
+    6.302663686681303e-08
+    1.181615530883472e-07
+    4.410609053416546e-07
+    3.449161305214893e-08
+    6.303401099298168e-08
+    1.823862518911561e-07
+    4.513543408725804e-07
+ 5.21e+10    
+    4.520688243730226e-07
+    1.827927157108261e-07
+    4.415545750861097e-07
+     6.30757900333126e-08
+    1.184282816914118e-07
+    4.415512867150404e-07
+     3.43831957029452e-08
+    6.308281882231249e-08
+    1.828193254585466e-07
+    4.520060059159414e-07
+ 5.26e+10    
+    4.527247896656287e-07
+    1.832267152231374e-07
+    4.420480248691548e-07
+    6.312241737086566e-08
+    1.186946731002444e-07
+      4.4204450519848e-07
+    3.427051338837294e-08
+    6.312912114352403e-08
+    1.832531171899195e-07
+     4.52662151993843e-07
+ 5.31e+10    
+    4.533852394406322e-07
+    1.836613995651987e-07
+    4.425443094140029e-07
+    6.316645914002113e-08
+    1.189607185892852e-07
+    4.425405565675815e-07
+    3.415360618013717e-08
+    6.317285778386417e-08
+    1.836875932221394e-07
+    4.533227777341831e-07
+ 5.36e+10    
+    4.540501728233235e-07
+    1.840967352527773e-07
+    4.430434251234632e-07
+    6.320786084108256e-08
+    1.192264114164148e-07
+    4.430394371859569e-07
+    3.403251681622493e-08
+      6.3213973656597e-08
+    1.841227200397518e-07
+    4.539878822920305e-07
+ 5.41e+10    
+    4.547195894480929e-07
+    1.845326891055694e-07
+    4.435453689482459e-07
+    6.324657282348353e-08
+    1.194917466944288e-07
+    4.435411439726534e-07
+    3.390729052798684e-08
+    6.325241841846196e-08
+    1.845584644224403e-07
+    4.546574653192197e-07
+ 5.46e+10    
+    4.553934894255428e-07
+       1.849692281935e-07
+    4.440501383574103e-07
+    6.328254991729302e-08
+    1.197567212677207e-07
+    4.440456743704076e-07
+    3.377797487217439e-08
+    6.328814613779878e-08
+    1.849947933943448e-07
+    4.553315269344794e-07
+ 5.51e+10    
+    4.560718733114318e-07
+     1.85406319786054e-07
+     4.44557731309491e-07
+     6.33157510882154e-08
+    1.200213335950026e-07
+    4.445530263156591e-07
+     3.36446195689389e-08
+    6.332111497729856e-08
+    1.854316741755959e-07
+    4.560100676945536e-07
+ 5.56e+10    
+    4.567547420772454e-07
+    1.858439313046795e-07
+    4.450681462253242e-07
+    6.334613911643697e-08
+    1.202855836386848e-07
+    4.450631982098853e-07
+    3.350727634623661e-08
+    6.335128689373862e-08
+     1.85869074136447e-07
+    4.566930885666627e-07
+ 5.61e+10    
+    4.574420970827715e-07
+    1.862820302782734e-07
+    4.455813819619028e-07
+    6.337368029897449e-08
+    1.205494727608226e-07
+    4.455761888928985e-07
+    3.336599879113719e-08
+    6.337862735594197e-08
+    1.863069607540997e-07
+    4.573805909023231e-07
+ 5.66e+10    
+    4.581339400504176e-07
+    1.867205843018231e-07
+     4.46097437788076e-07
+    6.339834417464308e-08
+    1.208130036259498e-07
+    4.460919976175975e-07
+    3.322084220766099e-08
+    6.340310508119948e-08
+    1.867453015722167e-07
+    4.580725764126894e-07
+ 5.71e+10    
+    4.588302730413989e-07
+    1.871595609977945e-07
+    4.466163133615289e-07
+    6.342010327065118e-08
+     1.21076180110293e-07
+    4.466106240267139e-07
+    3.307186348151705e-08
+    6.342469179022812e-08
+    1.871840641631373e-07
+    4.587690471455242e-07
+ 5.76e+10    
+    4.595310984336461e-07
+    1.875989279806219e-07
+     4.47138008707326e-07
+     6.34389328693829e-08
+    1.213390072174774e-07
+    4.471320681308517e-07
+    3.291912095101215e-08
+    6.344336197984675e-08
+    1.876232160928277e-07
+    4.594700054636341e-07
+ 5.81e+10    
+     4.60236418901387e-07
+    1.880386528235169e-07
+    4.476625241980657e-07
+    6.345481079403147e-08
+    1.216014909998208e-07
+    4.476563302883192e-07
+    3.276267428438372e-08
+    6.345909271272979e-08
+    1.880627248881034e-07
+    4.601754540248965e-07
+ 5.86e+10    
+    4.609462373963232e-07
+    1.884787030280932e-07
+    4.481898605351254e-07
+    6.346771721191863e-08
+    1.218636384854739e-07
+    4.481834111863503e-07
+    3.260258436286991e-08
+    6.347186342325329e-08
+    1.885025580065412e-07
+    4.608853957637164e-07
+ 5.91e+10    
+    4.616605571303632e-07
+      1.8891904599615e-07
+    4.487200187314905e-07
+    6.347763445389579e-08
+    1.221254576106161e-07
+    4.487133118235802e-07
+    3.243891316957449e-08
+    6.348165573864446e-08
+    1.889426828083737e-07
+    4.615998338739886e-07
+ 5.96e+10    
+    4.623793815597523e-07
+    1.893596490037137e-07
+    4.492530000956172e-07
+    6.348454684887895e-08
+    1.223869571565371e-07
+    4.492460334939286e-07
+     3.22717236835421e-08
+    6.348845331403681e-08
+    1.893830665307361e-07
+    4.623187717933312e-07
+ 6.01e+10    
+     4.63102714370606e-07
+    1.898004791770979e-07
+     4.49788806216496e-07
+    6.348844057185472e-08
+    1.226481466910797e-07
+    4.497815777715972e-07
+    3.210107977913526e-08
+    6.349224168088524e-08
+     1.89823676263695e-07
+    4.630422131887558e-07
+ 6.06e+10    
+    4.638305594656874e-07
+    1.902415034709296e-07
+     4.50327438949951e-07
+    6.348930350482597e-08
+    1.229090365143286e-07
+    4.503199464971359e-07
+    3.192704613007829e-08
+    6.349300810737788e-08
+    1.902644789283352e-07
+    4.637701619434862e-07
+ 6.11e+10    
+    4.645629209524922e-07
+    1.906826886478663e-07
+    4.508689004055598e-07
+    6.348712510902403e-08
+    1.231696376080191e-07
+    4.508611417645351e-07
+    3.174968811829937e-08
+    6.349074147026312e-08
+    1.907054412564777e-07
+     4.64502622145009e-07
+ 6.16e+10    
+    4.652998031323768e-07
+     1.91124001259958e-07
+    4.514131929348294e-07
+    6.348189630799573e-08
+    1.234299615885435e-07
+    4.514051659092598e-07
+    3.156907174721779e-08
+    6.348543213694177e-08
+    1.911465297720469e-07
+    4.652395980743091e-07
+ 6.21e+10    
+    4.660412104909085e-07
+    1.915654076316888e-07
+    4.519603191201435e-07
+    6.347360938023927e-08
+    1.236900206629136e-07
+    4.519520214971422e-07
+    3.138526355907561e-08
+    6.347707185718634e-08
+    1.915877107739827e-07
+    4.659810941961189e-07
+ 6.26e+10    
+    4.667871476891546e-07
+    1.920068738442135e-07
+    4.525102817643385e-07
+    6.346225786082539e-08
+    1.239498275879928e-07
+     4.52501711314022e-07
+    3.119833055676536e-08
+     6.34656536636667e-08
+    1.920289503205232e-07
+    4.667271151502186e-07
+ 6.31e+10    
+    4.675376195560273e-07
+     1.92448365721144e-07
+    4.530630838813191e-07
+    6.344783645121006e-08
+    1.242093956323495e-07
+     4.53054238356256e-07
+     3.10083401292484e-08
+    6.345117178068172e-08
+    1.924702142148798e-07
+    4.674776657437633e-07
+ 6.36e+10    
+    4.682926310815326e-07
+     1.92889848815454e-07
+    4.536187286869856e-07
+    6.343034093651622e-08
+    1.244687385403219e-07
+    4.536096058216626e-07
+    3.081535998097376e-08
+    6.343362154021674e-08
+     1.92911467992045e-07
+     4.68232750944459e-07
+ 6.41e+10    
+    4.690521874109111e-07
+    1.933312883975042e-07
+    4.541772195912036e-07
+    6.340976810973274e-08
+    1.247278704987756e-07
+    4.541678171014427e-07
+    3.061945806500707e-08
+    6.341299930506042e-08
+    1.933526769069277e-07
+    4.689923758747532e-07
+ 6.46e+10    
+     4.69816293839709e-07
+    1.937726494443564e-07
+    4.547385601899807e-07
+    6.338611570225104e-08
+    1.249868061057717e-07
+    4.547288757724225e-07
+    3.042070251971347e-08
+    6.338930239815837e-08
+    1.937938059233821e-07
+    4.697565458067293e-07
+ 6.51e+10    
+    4.705849558095136e-07
+    1.942138966298145e-07
+    4.553027542585882e-07
+    6.335938232022936e-08
+    1.252455603410223e-07
+     4.55292785589928e-07
+    3.021916160893749e-08
+    6.336252903797518e-08
+    1.942348197043317e-07
+    4.705252661579073e-07
+ 6.56e+10    
+    4.713581789045692e-07
+    1.946549943156679e-07
+    4.558698057447918e-07
+    6.332956738629991e-08
+    1.255041485384332e-07
+    4.558595504812228e-07
+    3.001490366571381e-08
+    6.333267827905319e-08
+     1.94675682602901e-07
+    4.712985424878362e-07
+ 6.61e+10    
+    4.721359688491335e-07
+    1.950959065436645e-07
+    4.564397187630142e-07
+    6.329667108623994e-08
+    1.257625863599055e-07
+    4.564291745394347e-07
+    2.980799703918495e-08
+     6.32997499577695e-08
+    1.951163586543848e-07
+    4.720763804953339e-07
+ 6.66e+10    
+    4.729183315054562e-07
+    1.955365970283957e-07
+    4.570124975885169e-07
+    6.326069432027596e-08
+    1.260208897709707e-07
+    4.570016620179146e-07
+    2.959851004489603e-08
+    6.326374464264718e-08
+    1.955568115690624e-07
+    4.728587860165198e-07
+ 6.71e+10    
+    4.737052728725297e-07
+    1.959770291509627e-07
+    4.575881466524691e-07
+    6.322163865849946e-08
+    1.262790750175623e-07
+    4.575770173249934e-07
+    2.938651091815125e-08
+    6.322466358887715e-08
+    1.959970047257529e-07
+    4.736457650234546e-07
+ 6.76e+10    
+    4.744967990853764e-07
+    1.964171659533245e-07
+    4.581666705370296e-07
+    6.317950630024312e-08
+    1.265371586041086e-07
+    4.581552450192421e-07
+     2.91720677706936e-08
+    6.318250869691205e-08
+    1.964369011662015e-07
+    4.744373236234684e-07
+ 6.81e+10    
+    4.752929164150314e-07
+    1.968569701334272e-07
+    4.587480739710867e-07
+    6.313430003708079e-08
+    1.267951572729085e-07
+    4.587363498050417e-07
+    2.895524855015442e-08
+    6.313728247460993e-08
+    1.968764635901645e-07
+    4.752334680590529e-07
+ 6.86e+10    
+     4.76093631269031e-07
+    1.972964040409502e-07
+    4.593323618263808e-07
+    6.308602321921815e-08
+    1.270530879842889e-07
+    4.593203365286525e-07
+    2.873612100271773e-08
+     6.30889880029022e-08
+    1.973156543510535e-07
+    4.760342047083976e-07
+ 6.91e+10    
+    4.768989501925378e-07
+    1.977354296736328e-07
+    4.599195391137102e-07
+    6.303467972482778e-08
+    1.273109678980879e-07
+    4.599072101744262e-07
+    2.851475263863697e-08
+    6.303762890451383e-08
+    1.977544354523075e-07
+    4.768395400864257e-07
+ 6.96e+10    
+    4.777088798698839e-07
+    1.981740086742728e-07
+    4.605096109798786e-07
+    6.298027393249169e-08
+     1.27568814355696e-07
+    4.604969758616082e-07
+     2.82912107005001e-08
+    6.298320931568585e-08
+    1.981927685443202e-07
+    4.776494808463763e-07
+ 7.01e+10    
+     4.78523427126725e-07
+    1.986121023282055e-07
+    4.611025827046037e-07
+    6.292281069613992e-08
+    1.278266448632085e-07
+    4.610896388412807e-07
+    2.806556213427153e-08
+     6.29257338605632e-08
+    1.986306149218671e-07
+    4.784640337818768e-07
+ 7.06e+10    
+    4.793425989325754e-07
+    1.990496715613293e-07
+    4.616984596980774e-07
+    6.286229532261862e-08
+    1.280844770752071e-07
+    4.616852044937937e-07
+     2.78378735631241e-08
+    6.286520762824604e-08
+    1.990679355222215e-07
+    4.792832058295332e-07
+ 7.11e+10    
+    4.801664024038669e-07
+    1.994866769386382e-07
+    4.622972474985933e-07
+    6.279873355144173e-08
+    1.283423287791095e-07
+    4.622836783262803e-07
+    2.760821126368708e-08
+    6.280163615197412e-08
+    1.995046909234966e-07
+     4.80107004071876e-07
+ 7.16e+10    
+    4.809948448073282e-07
+    1.999230786631911e-07
+    4.628989517705344e-07
+    6.273213153681397e-08
+    1.286002178803329e-07
+    4.628850659706973e-07
+    2.737664114489556e-08
+    6.273502539073098e-08
+    1.999408413437668e-07
+    4.809354357408805e-07
+ 7.21e+10    
+    4.818279335639194e-07
+    2.003588365755411e-07
+    4.635035783027106e-07
+    6.266249583158627e-08
+    1.288581623880426e-07
+    4.634893731820489e-07
+    2.714322872932559e-08
+    6.266538171274643e-08
+     2.00376346640396e-07
+    4.817685082216946e-07
+ 7.26e+10    
+    4.826656762529744e-07
+    2.007939101535903e-07
+    4.641111330070321e-07
+    6.258983337309849e-08
+    1.291161804011879e-07
+    4.640966058368088e-07
+    2.690803913667111e-08
+    6.259271188092295e-08
+    2.008111663098606e-07
+    4.826062290569302e-07
+ 7.31e+10    
+    4.835080806168066e-07
+    2.012282585127945e-07
+    4.647216219171284e-07
+    6.251415147074885e-08
+    1.293742900953619e-07
+    4.647067699318417e-07
+     2.66711370696044e-08
+    6.251702304009125e-08
+    2.012452594880251e-07
+    4.834486059511797e-07
+ 7.36e+10    
+    4.843551545656167e-07
+    2.016618404067732e-07
+    4.653350511876404e-07
+    6.243545779519429e-08
+    1.296325097097412e-07
+    4.653198715833126e-07
+     2.64325868016787e-08
+    6.243832270582394e-08
+    2.016785849507077e-07
+    4.842956467759155e-07
+ 7.41e+10    
+    4.852069061826861e-07
+    2.020946142283079e-07
+    4.659514270936214e-07
+    6.235376036898329e-08
+    1.298908575346962e-07
+    4.659359170260778e-07
+    2.619245216724673e-08
+     6.23566187547428e-08
+    2.021111011146273e-07
+    4.851473595747244e-07
+ 7.46e+10    
+    4.860633437299098e-07
+    2.025265380105139e-07
+    4.665707560300008e-07
+    6.226906755867193e-08
+     1.30149351899479e-07
+    4.665549126132115e-07
+    2.595079655341199e-08
+     6.22719194163628e-08
+    2.025427660387044e-07
+    4.860037525687677e-07
+ 7.51e+10    
+    4.869244756535364e-07
+    2.029575694285623e-07
+    4.671930445115811e-07
+    6.218138806812397e-08
+    1.304080111605905e-07
+    4.671768648157587e-07
+    2.570768289357589e-08
+     6.21842332661718e-08
+    2.029735374256146e-07
+    4.868648341625371e-07
+ 7.56e+10    
+    4.877903105902093e-07
+    2.033876658014783e-07
+    4.678182991731293e-07
+    6.209073093309743e-08
+    1.306668536899653e-07
+    4.678017802228881e-07
+    2.546317366293401e-08
+    6.209356921984572e-08
+    2.034033726237291e-07
+    4.877306129499137e-07
+ 7.61e+10    
+     4.88660857373173e-07
+    2.038167840942873e-07
+    4.684465267695792e-07
+    6.199710551681459e-08
+    1.309258978637475e-07
+    4.684296655419772e-07
+    2.521733087528005e-08
+    6.199993652868543e-08
+    2.038322286292471e-07
+    4.886010977203119e-07
+ 7.66e+10    
+    4.895361250387722e-07
+    2.042448809205045e-07
+    4.690777341768294e-07
+    6.190052150667776e-08
+    1.311851620511272e-07
+    4.690605275992335e-07
+    2.497021608149045e-08
+    6.190334477607755e-08
+    2.042600620885542e-07
+    4.894762974652272e-07
+ 7.71e+10    
+    4.904161228330524e-07
+    2.046719125447074e-07
+    4.697119283922772e-07
+    6.180098891182515e-08
+    1.314446646034616e-07
+    4.696943733404596e-07
+    2.472189036931573e-08
+    6.180380387481828e-08
+    2.046868293010101e-07
+    4.903562213847808e-07
+ 7.76e+10    
+    4.913008602186204e-07
+    2.050978348854488e-07
+    4.703491165359243e-07
+    6.169851806156116e-08
+    1.317044238432633e-07
+    4.703312098317915e-07
+    2.447241436424856e-08
+    6.170132406540096e-08
+    2.051124862217198e-07
+    4.912408788946009e-07
+ 7.81e+10    
+    4.921903468815535e-07
+    2.055226035183617e-07
+    4.709893058516667e-07
+    6.159311960454734e-08
+    1.319644580537313e-07
+    4.709710442610114e-07
+    2.422184823178906e-08
+    6.159591591499849e-08
+    2.055369884647281e-07
+    4.921302796327026e-07
+ 7.86e+10    
+    4.930845927385754e-07
+    2.059461736794261e-07
+    4.716325037084824e-07
+    6.148480450876539e-08
+    1.322247854680301e-07
+    4.716138839388283e-07
+    2.397025168040676e-08
+    6.148759031727109e-08
+    2.059602913062386e-07
+    4.930244334666518e-07
+ 7.91e+10    
+    4.939836079442275e-07
+    2.063685002684432e-07
+    4.722787176022653e-07
+    6.137358406212491e-08
+    1.324854242587701e-07
+    4.722597363004205e-07
+     2.37176839656452e-08
+    6.137635849272896e-08
+      2.0638234968815e-07
+    4.939233505007658e-07
+ 7.96e+10    
+    4.948874028982451e-07
+     2.06789537852708e-07
+    4.729279551574714e-07
+    6.125946987351946e-08
+    1.327463925275711e-07
+    4.729086089071703e-07
+    2.346420389475226e-08
+    6.126223198976937e-08
+     2.06803118221712e-07
+     4.94827041083413e-07
+ 8.01e+10    
+    4.957959882529539e-07
+    2.072092406707532e-07
+    4.735802241291981e-07
+    6.114247387457408e-08
+    1.330077082945761e-07
+    4.735605094486881e-07
+    2.320986983220638e-08
+    6.114522268614241e-08
+    2.072225511913007e-07
+    4.957355158144637e-07
+ 8.06e+10    
+    4.967093749208332e-07
+    2.076275626363736e-07
+    4.742355324052827e-07
+    6.102260832176575e-08
+    1.332693894879729e-07
+    4.742154457448584e-07
+    2.295473970550039e-08
+    6.102534279099075e-08
+    2.076406025584742e-07
+     4.96648785552781e-07
+ 8.11e+10    
+    4.976275740820382e-07
+     2.08044457342672e-07
+    4.748938880087288e-07
+    6.089988579900343e-08
+    1.335314539336577e-07
+    4.748734257480897e-07
+    2.269887101170166e-08
+     6.09026048472821e-08
+    2.080572259659607e-07
+    4.975668614237658e-07
+ 8.16e+10    
+    4.985505971920248e-07
+    2.084598780662787e-07
+    4.755552991001947e-07
+    6.077431922047037e-08
+    1.337939193445502e-07
+    4.755344575459331e-07
+    2.244232082393413e-08
+    6.077702173448043e-08
+    2.084723747419763e-07
+    4.984897548269817e-07
+ 8.21e+10    
+    4.994784559892669e-07
+    2.088737777717202e-07
+    4.762197739806899e-07
+    6.064592183394936e-08
+    1.340568033101484e-07
+    4.761985493636649e-07
+    2.218514579837705e-08
+    6.064860667175249e-08
+    2.088860019045824e-07
+    4.994174774437922e-07
+ 8.26e+10    
+    5.004111625029005e-07
+    2.092861091158468e-07
+    4.768873210945123e-07
+    6.051470722423027e-08
+    1.343201232859092e-07
+    4.768657095671653e-07
+     2.19274021812275e-08
+    6.051737322118254e-08
+    2.092980601660958e-07
+    5.003500412450722e-07
+ 8.31e+10    
+    5.013487290604457e-07
+    2.096968244523809e-07
+    4.775579490321951e-07
+    6.038068931683557e-08
+    1.345838965824825e-07
+    4.775359466658305e-07
+    2.166914581573843e-08
+    6.038333529150603e-08
+    2.097085019377223e-07
+    5.012874584988613e-07
+ 8.36e+10    
+    5.022911682955583e-07
+    2.101058758365639e-07
+    4.782316665337164e-07
+    6.024388238192351e-08
+    1.348481403549779e-07
+    4.782092693158245e-07
+    2.141043214903975e-08
+    6.024650714169655e-08
+    2.101172793341561e-07
+    5.022297417780995e-07
+ 8.41e+10    
+    5.032384931557006e-07
+    2.105132150299125e-07
+    4.789084824918412e-07
+    6.010430103833312e-08
+      1.3511287159198e-07
+    4.788856863233319e-07
+    2.115131623891488e-08
+    6.010690338495252e-08
+     2.10524344178379e-07
+    5.031769039683123e-07
+ 8.46e+10    
+    5.041907169098924e-07
+    2.109187935050064e-07
+    4.795884059556939e-07
+    5.996196025768567e-08
+    1.353781071045494e-07
+    4.795652066480114e-07
+    2.089185276022469e-08
+    5.996453899267371e-08
+    2.109296480064653e-07
+    5.041289582752949e-07
+ 8.51e+10    
+    5.051478531563602e-07
+    2.113225624503849e-07
+     4.80271446134236e-07
+    5.981687536861632e-08
+    1.356438635149623e-07
+    4.802478394066779e-07
+    2.063209601095425e-08
+    5.981942929849895e-08
+    2.113331420725012e-07
+    5.050859182328031e-07
+ 8.56e+10    
+     5.06109915830233e-07
+    2.117244727755403e-07
+     4.80957612400209e-07
+    5.966906206100868e-08
+    1.359101572455285e-07
+    4.809335938770264e-07
+    2.037209991788764e-08
+    5.967159000241857e-08
+    2.117347773535492e-07
+    5.060477977101558e-07
+ 8.61e+10    
+    5.070769192111223e-07
+    2.121244751159163e-07
+    4.816469142939148e-07
+     5.95185363902324e-08
+    1.361770045069696e-07
+    4.816224795014617e-07
+    2.011191804168528e-08
+    5.952103717489218e-08
+    2.121345045547538e-07
+    5.070146109198781e-07
+ 8.66e+10    
+    5.080488779307585e-07
+    2.125225198379956e-07
+    4.823393615273761e-07
+    5.936531478140075e-08
+    1.364444212868083e-07
+    4.823145058912839e-07
+    1.985160358131507e-08
+    5.936778726087101e-08
+    2.125322741143211e-07
+    5.079863724252336e-07
+ 8.71e+10    
+    5.090258069804632e-07
+    2.129185570444571e-07
+    4.830349639884083e-07
+    5.920941403359259e-08
+    1.367124233375614e-07
+    4.830096828307407e-07
+    1.959120937804071e-08
+    5.921185708393179e-08
+    2.129280362088333e-07
+    5.089630971477318e-07
+ 8.76e+10    
+    5.100077217186837e-07
+    2.133125365794327e-07
+    4.837337317450054e-07
+    5.905085132390223e-08
+    1.369810261647494e-07
+    4.837080202813155e-07
+    1.933078791828975e-08
+     5.90532638501491e-08
+    2.133217407583845e-07
+    5.099448003746171e-07
+ 8.81e+10    
+    5.109946378783683e-07
+    2.137044080337003e-07
+    4.844356750496699e-07
+    5.888964421150698e-08
+    1.372502450146728e-07
+    4.844095283862251e-07
+    1.907039133618916e-08
+    5.889202515198742e-08
+    2.137133374318774e-07
+    5.109314977662322e-07
+ 8.86e+10    
+    5.119865715743394e-07
+    2.140941207500206e-07
+    4.851408043441018e-07
+      5.8725810641631e-08
+     1.37520094862033e-07
+    4.851142174749146e-07
+    1.881007141475146e-08
+    5.872815897210197e-08
+    2.141027756523289e-07
+    5.119232053633396e-07
+ 8.91e+10    
+    5.129835393105614e-07
+    2.144816238285292e-07
+    4.858491302636712e-07
+    5.855936894931932e-08
+    1.377905903973908e-07
+    4.858220980676891e-07
+     1.85498795865103e-08
+    5.856168368688451e-08
+    2.144900046022842e-07
+    5.129199395944026e-07
+ 8.96e+10    
+    5.139855579873496e-07
+     2.14866866132119e-07
+    4.865606636422884e-07
+    5.839033786308451e-08
+    1.380617460143887e-07
+    4.865331808805415e-07
+    1.828986693316945e-08
+    5.839261807005015e-08
+    2.148749732292271e-07
+    5.139217172827468e-07
+ 9.01e+10    
+    5.149926449084943e-07
+    2.152497962919102e-07
+    4.872754155172152e-07
+    5.821873650846345e-08
+    1.383335757968158e-07
+    4.872474768300125e-07
+    1.803008418395881e-08
+     5.82209812958961e-08
+    2.152576302510599e-07
+    5.149285556536755e-07
+ 9.06e+10    
+    5.160048177882946e-07
+    2.156303627127848e-07
+    4.879933971341011e-07
+    5.804458441132831e-08
+    1.386060935053532e-07
+    4.879649970380687e-07
+    1.777058171328107e-08
+    5.804679294242855e-08
+    2.156379241615757e-07
+    5.159404723414286e-07
+ 9.11e+10    
+     5.17022094758533e-07
+    2.160085135789341e-07
+    4.887146199519204e-07
+    5.786790150108226e-08
+    1.388793125643535e-07
+    4.886857528373769e-07
+    1.751140953705467e-08
+    5.787007299447242e-08
+    2.160158032361222e-07
+    5.169574853962138e-07
+ 9.16e+10    
+    5.180444943752729e-07
+    2.163841968594351e-07
+    4.894390956482124e-07
+    5.768870811362539e-08
+    1.391532460481876e-07
+     4.89409755776248e-07
+    1.725261730801464e-08
+    5.769084184629527e-08
+    2.163912155371388e-07
+    5.179796132909183e-07
+ 9.21e+10    
+    5.190720356257085e-07
+    2.167573603140072e-07
+    4.901668361243163e-07
+    5.750702499419354e-08
+     1.39427906667542e-07
+    4.901370176241591e-07
+    1.699425430993495e-08
+     5.75091203043328e-08
+    2.167641089199016e-07
+    5.190068749279363e-07
+ 9.26e+10    
+    5.201047379347512e-07
+    2.171279514986196e-07
+    4.908978535107346e-07
+    5.732287329992412e-08
+    1.397033067554325e-07
+    4.908675503768434e-07
+    1.673636945041815e-08
+    5.732492958952172e-08
+    2.171344310381328e-07
+    5.200392896457611e-07
+ 9.31e+10    
+    5.211426211716182e-07
+    2.174959177713426e-07
+     4.91632160172339e-07
+    5.713627460235371e-08
+    1.399794582532248e-07
+    4.916013662619068e-07
+    1.647901125292789e-08
+    5.713829133954653e-08
+    2.175021293499192e-07
+    5.210768772255309e-07
+ 9.36e+10    
+    5.221857056563098e-07
+    2.178612062981285e-07
+    4.923697687141344e-07
+    5.694725088950558e-08
+    1.402563726961829e-07
+    4.923384777442835e-07
+    1.622222784709698e-08
+    5.694922761082403e-08
+    2.178671511234119e-07
+    5.221196578974554e-07
+ 9.41e+10    
+    5.232340121659411e-07
+     2.18223764058752e-07
+    4.931106919865579e-07
+    5.675582456805693e-08
+    1.405340611990355e-07
+    4.930788975318221e-07
+    1.596606695822786e-08
+    5.675776088027388e-08
+    2.182294434427854e-07
+    5.231676523471446e-07
+ 9.46e+10    
+    5.242875619409363e-07
+    2.185835378526657e-07
+    4.938549430912454e-07
+    5.656201846505875e-08
+    1.408125344414497e-07
+    4.938226385809886e-07
+    1.571057589521686e-08
+    5.656391404696806e-08
+    2.185889532141875e-07
+    5.242208817218145e-07
+ 9.51e+10    
+    5.253463766912071e-07
+    2.189404743050938e-07
+    4.946025353866522e-07
+    5.636585582963604e-08
+    1.410918026530991e-07
+    4.945697141024819e-07
+    1.545580153757966e-08
+    5.636771043352602e-08
+    2.189456271717042e-07
+     5.25279367636381e-07
+ 9.56e+10    
+     5.26410478602136e-07
+    2.192945198730778e-07
+    4.953534824938297e-07
+    5.616736033440184e-08
+    1.413718755988118e-07
+    4.953201375671336e-07
+     1.52017903208015e-08
+    5.616917378727504e-08
+    2.192994118834685e-07
+    5.263431321794305e-07
+ 9.61e+10    
+    5.274798903404211e-07
+    2.196456208516019e-07
+     4.96107798302139e-07
+    5.596655607676082e-08
+     1.41652762563478e-07
+    4.960739227117532e-07
+    1.494858822079371e-08
+    5.596832828138401e-08
+     2.19650253757767e-07
+     5.27412197919073e-07
+ 9.66e+10    
+     5.28554635059872e-07
+    2.199937233798467e-07
+    4.968654969751383e-07
+    5.576346757993074e-08
+    1.419344723368498e-07
+    4.968310835448139e-07
+    1.469624073688565e-08
+    5.576519851562739e-08
+    2.199980990492801e-07
+    5.284865879086879e-07
+ 9.71e+10    
+    5.296347364069926e-07
+    2.203387734474354e-07
+    4.976265929564356e-07
+    5.555811979394527e-08
+     1.42217013198244e-07
+    4.975916343527102e-07
+    1.444479287360834e-08
+    5.555980951712394e-08
+    2.203428938654082e-07
+    5.295663256925155e-07
+ 9.76e+10    
+    5.307202185265325e-07
+     2.20680716900887e-07
+    4.983911009756717e-07
+    5.535053809643325e-08
+    1.425003929011015e-07
+    4.983555897054783e-07
+    1.419428912122544e-08
+    5.535218674083779e-08
+    2.206845841725136e-07
+    5.306514353111206e-07
+ 9.81e+10    
+    5.318111060667862e-07
+    2.210194994499568e-07
+    4.991590360543392e-07
+    5.514074829312242e-08
+    1.427846186575389e-07
+    4.991229644629249e-07
+    1.394477343501884e-08
+    5.514235606994607e-08
+    2.210231158024936e-07
+    5.317419413067324e-07
+ 9.86e+10    
+    5.329074241848308e-07
+    2.213550666742864e-07
+    4.999304135118924e-07
+    5.492877661846074e-08
+    1.430696971227429e-07
+    4.998937737806296e-07
+    1.369628921335212e-08
+    5.493034381608976e-08
+    2.213584344592317e-07
+    5.328378687284811e-07
+ 9.91e+10    
+       5.340091985516e-07
+    2.216873640299532e-07
+    5.007052489716636e-07
+    5.471464973585386e-08
+    1.433556343794134e-07
+    5.006680331160452e-07
+    1.344887927449681e-08
+    5.471617671950164e-08
+    2.216904857252425e-07
+    5.339392431373572e-07
+ 9.96e+10    
+    5.351164553568179e-07
+    2.220163368562281e-07
+    5.014835583668535e-07
+    5.449839473801795e-08
+    1.436424359220034e-07
+    5.014457582345049e-07
+    1.320258583226983e-08
+    5.449988194894629e-08
+    2.220192150683974e-07
+    5.350460906112408e-07
+ 1.001e+11   
+    5.362292213137547e-07
+    2.223419303823775e-07
+    5.022653579466317e-07
+    5.428003914704454e-08
+    1.439301066412048e-07
+    5.022269652154871e-07
+    1.295745047040049e-08
+    5.428148710169929e-08
+    2.223445678486575e-07
+    5.361584377495577e-07
+ 1.006e+11   
+    5.373475236638644e-07
+    2.226640897346053e-07
+    5.030506642821461e-07
+     5.40596109145039e-08
+    1.442186508080962e-07
+    5.030116704585026e-07
+     1.27135141158976e-08
+    5.406102020329327e-08
+    2.226664893250335e-07
+    5.372763116779634e-07
+ 1.011e+11   
+    5.384713901812241e-07
+    2.229827599429765e-07
+    5.038394942724238e-07
+    5.383713842138966e-08
+     1.44508072058598e-07
+    5.037998906893522e-07
+    1.247081701109096e-08
+     5.38385097072985e-08
+    2.229849246625468e-07
+    5.383997400527081e-07
+ 1.016e+11   
+    5.396008491768202e-07
+    2.232978859486402e-07
+    5.046318651505519e-07
+    5.361265047812915e-08
+    1.447983733777809e-07
+    5.045916429661489e-07
+    1.222939868467896e-08
+    5.361398449497734e-08
+    2.232998189393411e-07
+    5.395287510649834e-07
+ 1.021e+11   
+    5.407359295027138e-07
+    2.236094126110073e-07
+    5.054277944895901e-07
+    5.338617632437767e-08
+    1.450895570843651e-07
+    5.053869446854742e-07
+    1.198929792159602e-08
+    5.338747387497187e-08
+    2.236111171538735e-07
+    5.406633734450037e-07
+ 1.026e+11   
+    5.418766605558891e-07
+    2.239172847150472e-07
+    5.062273002085204e-07
+    5.315774562897893e-08
+    1.453816248152261e-07
+    5.061858135883791e-07
+    1.175055273184501e-08
+    5.315900758292118e-08
+    2.239187642322102e-07
+    5.418036364659222e-07
+ 1.031e+11   
+     5.43023072282133e-07
+    2.242214469787798e-07
+    5.070304005782467e-07
+    5.292738848973928e-08
+    1.456745775099378e-07
+    5.069882677663597e-07
+     1.15132003183437e-08
+    5.292861578107516e-08
+    2.242227050354453e-07
+    5.429495699476186e-07
+ 1.036e+11   
+    5.441751951794976e-07
+    2.245218440607469e-07
+    5.078371142274076e-07
+    5.269513543336646e-08
+    1.459684153955923e-07
+    5.077943256675454e-07
+    1.127727704362975e-08
+    5.269632905794538e-08
+    2.245228843672456e-07
+    5.441012042602484e-07
+ 1.041e+11   
+    5.453330603017614e-07
+    2.248184205677573e-07
+    5.086474601484002e-07
+    5.246101741536837e-08
+    1.462631379716244e-07
+    5.086040061025087e-07
+    1.104281839570717e-08
+     5.24621784279436e-08
+    2.248192469814212e-07
+    5.452585703276361e-07
+ 1.046e+11   
+    5.464966992615637e-07
+    2.251111210625644e-07
+    5.094614577030098e-07
+    5.222506581989114e-08
+    1.465587439948863e-07
+    5.094173282501979e-07
+    1.080985895298138e-08
+    5.222619533111604e-08
+    2.251117375897284e-07
+    5.464216996304201e-07
+ 1.051e+11   
+    5.476661442333946e-07
+    2.253998900718061e-07
+    5.102791266282955e-07
+    5.198731245981884e-08
+    1.468552314648759e-07
+    5.102343116638117e-07
+    1.057843234809137e-08
+    5.198841163292108e-08
+    2.254003008696494e-07
+    5.475906242090824e-07
+ 1.056e+11   
+    5.488414279563553e-07
+    2.256846720939342e-07
+    5.111004870421601e-07
+    5.174778957684885e-08
+    1.471525976092119e-07
+    5.110549762766326e-07
+    1.034857123117515e-08
+    5.174885962407467e-08
+    2.256848814723777e-07
+    5.487653766666519e-07
+ 1.061e+11   
+    5.500225837366978e-07
+    2.259654116073657e-07
+    5.119255594490762e-07
+    5.150652984157027e-08
+    1.474508388692946e-07
+    5.118793424076262e-07
+    1.012030723205291e-08
+    5.150757202052568e-08
+    2.259654240308769e-07
+    5.499459901713168e-07
+ 1.066e+11   
+    5.512096454501755e-07
+    2.262420530786142e-07
+    5.127543647454646e-07
+    5.126356635384196e-08
+    1.477499508862851e-07
+     5.12707430767193e-07
+     9.89367092171884e-09
+    5.126458196350553e-08
+    2.262418731680418e-07
+    5.511324984587056e-07
+ 1.071e+11   
+    5.524026475440666e-07
+    2.265145409706015e-07
+    5.135869242252657e-07
+    5.101893264315783e-08
+    1.480499284873678e-07
+    5.135392624626608e-07
+    9.668691773269475e-09
+    5.101992301977004e-08
+    2.265141735049469e-07
+    5.523249358340099e-07
+ 1.076e+11   
+    5.536016250391034e-07
+    2.267828197510699e-07
+    5.144232595852014e-07
+    5.077266266918738e-08
+    1.483507656722726e-07
+      5.1437485900375e-07
+    9.445398121711445e-09
+    5.077362918193086e-08
+    2.267822696691781e-07
+    5.535233371738349e-07
+ 1.081e+11   
+    5.548066135309913e-07
+    2.270468339010328e-07
+    5.152633929299447e-07
+     5.05247908225726e-08
+     1.48652455600208e-07
+    5.152142423078783e-07
+    9.223817123701148e-09
+    5.052573486904986e-08
+    2.270461063033059e-07
+    5.547277379278176e-07
+ 1.086e+11   
+    5.560176491918698e-07
+    2.273065279233773e-07
+    5.161073467773744e-07
+     5.02753519257527e-08
+    1.489549905771263e-07
+    5.160574347054474e-07
+    9.003974716132609e-09
+    5.027627492731963e-08
+    2.273056280734214e-07
+     5.55938174120019e-07
+ 1.091e+11   
+    5.572347687713194e-07
+    2.275618463514482e-07
+    5.169551440634057e-07
+     5.00243812341411e-08
+    1.492583620433367e-07
+    5.169044589449608e-07
+    8.785895574613147e-09
+    5.002528463099619e-08
+    2.275607796776574e-07
+    5.571546823500099e-07
+ 1.096e+11   
+    5.584580095972408e-07
+    2.278127337578384e-07
+    5.178068081469604e-07
+     4.97719144373915e-08
+    1.495625605616298e-07
+    5.177553381979029e-07
+    8.569603071111854e-09
+    4.977279968363423e-08
+    2.278115058549863e-07
+    5.583772997937673e-07
+ 1.101e+11   
+    5.596874095763983e-07
+     2.28059134763031e-07
+    5.186623628146025e-07
+    4.951798766102739e-08
+    1.498675758056972e-07
+    5.186100960637291e-07
+    8.355119231527864e-09
+    4.951885621938512e-08
+    2.280577513938311e-07
+     5.59606064204211e-07
+ 1.106e+11   
+    5.609230071947578e-07
+    2.283009940443544e-07
+    5.195218322851471e-07
+    4.926263746819517e-08
+    1.501733965491952e-07
+     5.19468756574476e-07
+     8.14246469243839e-09
+    4.926349080477142e-08
+    2.282994611408571e-07
+    5.608410139115788e-07
+ 1.111e+11   
+    5.621648415174341e-07
+    2.285382563447321e-07
+    5.203852412140558e-07
+     4.90059008617788e-08
+    1.504800106550547e-07
+    5.203313441993299e-07
+    7.931658657974457e-09
+    4.900674044055749e-08
+     2.28536580009805e-07
+    5.620821878234129e-07
+ 1.116e+11   
+    5.634129521884831e-07
+    2.287708664815691e-07
+    5.212526146977102e-07
+    4.874781528682199e-08
+    1.507874050655807e-07
+    5.211978838490411e-07
+    7.722718856045558e-09
+    4.874864256405156e-08
+    2.287690529902724e-07
+     5.63329625424359e-07
+ 1.121e+11   
+    5.646673794302947e-07
+    2.289987693556305e-07
+    5.221239782775424e-07
+    4.848841863315637e-08
+    1.510955657927939e-07
+    5.220684008801761e-07
+    7.515661494734642e-09
+    4.848923505165937e-08
+    2.289968251565487e-07
+     5.64583366775622e-07
+ 1.126e+11   
+    5.659281640427835e-07
+    2.292219099598453e-07
+    5.229993579438626e-07
+     4.82277492384111e-08
+    1.514044779095417e-07
+    5.229429210991297e-07
+    7.310501218094594e-09
+     4.82285562217636e-08
+    2.292198416763869e-07
+    5.658434525141403e-07
+ 1.131e+11   
+    5.671953474022018e-07
+    2.294402333881908e-07
+    5.238787801397138e-07
+    4.796584589145278e-08
+    1.517141255411002e-07
+    5.238214707660889e-07
+    7.107251062379865e-09
+    4.796664483802126e-08
+     2.29438047819792e-07
+    5.671099238514761e-07
+ 1.136e+11   
+    5.684689714597133e-07
+    2.296536848443207e-07
+    5.247622717643833e-07
+     4.77027478360428e-08
+     1.52024491857231e-07
+    5.247040765987442e-07
+    6.905922411831553e-09
+    4.770354011300288e-08
+    2.296513889676652e-07
+    5.683828225724252e-07
+ 1.141e+11   
+    5.697490787396729e-07
+    2.298622096503293e-07
+    5.256498601768168e-07
+    4.743849477497198e-08
+     1.52335559065132e-07
+    5.255907657757572e-07
+    6.706524954782569e-09
+    4.743928171213994e-08
+    2.298598106204351e-07
+    5.696621910333114e-07
+ 1.146e+11   
+    5.710357123375985e-07
+    2.300657532552477e-07
+    5.265415731988866e-07
+    4.717312687460933e-08
+    1.526473084027354e-07
+    5.264815659402891e-07
+    6.509066639832599e-09
+    4.717390975833506e-08
+    2.300632584065699e-07
+    5.709480721599938e-07
+ 1.151e+11   
+    5.723289159177892e-07
+     2.30264261243398e-07
+    5.274374391183299e-07
+    4.690668476984877e-08
+    1.529597201327182e-07
+    5.273765052030455e-07
+    6.313553632150037e-09
+    4.690746483671181e-08
+    2.302616780908367e-07
+     5.72240509445568e-07
+ 1.156e+11   
+    5.736287337107675e-07
+    2.304576793426913e-07
+    5.283374866917365e-07
+    4.663920956946486e-08
+    1.532727735373062e-07
+    5.282756121453635e-07
+    6.119990270141619e-09
+     4.66399880000317e-08
+    2.304550155825554e-07
+    5.735395469478031e-07
+ 1.161e+11   
+    5.749352105103574e-07
+    2.306459534325339e-07
+    5.292417451471473e-07
+    4.637074286211157e-08
+    1.535864469134715e-07
+    5.291789158221147e-07
+    5.928379022428824e-09
+    4.637152077456889e-08
+    2.306432169434389e-07
+    5.748452292862884e-07
+ 1.166e+11   
+    5.762483916704694e-07
+    2.308290295516306e-07
+     5.30150244186607e-07
+    4.610132672258093e-08
+    1.539007175689855e-07
+    5.300864457643118e-07
+    5.738720445180524e-09
+    4.610210516637722e-08
+     2.30826228395342e-07
+    5.761576016392735e-07
+ 1.171e+11   
+    5.775683231016824e-07
+    2.310068539053644e-07
+    5.310630139885725e-07
+    4.583100371883617e-08
+    1.542155618190737e-07
+    5.309982319816527e-07
+    5.551013140196742e-09
+    4.583178366827465e-08
+    2.310039963276008e-07
+    5.774767097402689e-07
+ 1.176e+11   
+    5.788950512675322e-07
+    2.311793728729056e-07
+    5.319800852101129e-07
+     4.55598169194149e-08
+    1.545309549836926e-07
+    5.319143049649497e-07
+    5.365253713207495e-09
+    4.556059926732204e-08
+    2.311764673040503e-07
+    5.788025998743976e-07
+ 1.181e+11   
+    5.802286231805147e-07
+    2.313465330139015e-07
+    5.329014889890572e-07
+    4.528780990155901e-08
+    1.548468713855559e-07
+     5.32834695688358e-07
+    5.181436733194308e-09
+     4.52885954528241e-08
+    2.313435880696697e-07
+    5.801353188744528e-07
+ 1.186e+11   
+    5.815690863979335e-07
+    2.315082810746433e-07
+     5.33827256945839e-07
+    4.501502675985618e-08
+    1.551632843487145e-07
+    5.337594356115684e-07
+    4.999554692154828e-09
+    4.501581622510664e-08
+    2.315053055567168e-07
+    5.814749141167648e-07
+ 1.191e+11   
+    5.829164890174782e-07
+    2.316645639937938e-07
+    5.347574211855836e-07
+    4.474151211565685e-08
+    1.554801661978696e-07
+    5.346885566818112e-07
+    4.819597966028314e-09
+    4.474230610487801e-08
+    2.316615668903481e-07
+    5.828214335168762e-07
+ 1.196e+11   
+    5.842708796726295e-07
+    2.318153289074936e-07
+    5.356920142998189e-07
+    4.446731112708415e-08
+    1.557974882582598e-07
+    5.356220913358426e-07
+    4.641554776164034e-09
+    4.446811014333617e-08
+    2.318123193936897e-07
+    5.841749255249539e-07
+ 1.201e+11   
+    5.856323075279416e-07
+    2.319605231537935e-07
+    5.366310693682733e-07
+    4.419246949987282e-08
+    1.561152208560682e-07
+    5.365600725019329e-07
+    4.465411152163636e-09
+    4.419327393300174e-08
+    2.319575105922051e-07
+    5.855354391211171e-07
+ 1.206e+11   
+    5.870008222741076e-07
+    2.321000942763395e-07
+    5.375746199607509e-07
+    4.391703349893125e-08
+    1.564333333196016e-07
+     5.37502533601831e-07
+    4.291150895503667e-09
+    4.391784361940654e-08
+    2.320970882173287e-07
+    5.869030238106239e-07
+ 1.211e+11   
+    5.883764741230202e-07
+    2.322339900272574e-07
+    5.385227001388454e-07
+    4.364104996081149e-08
+    1.567517939809076e-07
+    5.384495085527393e-07
+    4.118755544619028e-09
+    4.364186591359967e-08
+    2.322310002093126e-07
+    5.882777296188387e-07
+ 1.216e+11   
+    5.897593138027154e-07
+    2.323621583691388e-07
+    5.394753444580065e-07
+    4.336456630697789e-08
+     1.57070570177761e-07
+    5.394010317693321e-07
+    3.948204340998804e-09
+    4.336538810554644e-08
+    2.323591947190836e-07
+    5.896596070863585e-07
+ 1.221e+11   
+    5.911493925522896e-07
+    2.324845474759187e-07
+    5.404325879694297e-07
+    4.308763055812606e-08
+    1.573896282563344e-07
+    5.403571381660403e-07
+    3.779474196733527e-09
+    4.308845807848991e-08
+    2.324816201091771e-07
+     5.91048707263939e-07
+ 1.226e+11   
+    5.925467621169134e-07
+    2.326011057327394e-07
+     5.41394466222505e-07
+     4.28102913494704e-08
+    1.577089335741611e-07
+    5.413178631594414e-07
+    3.612539663665097e-09
+    4.281112432443336e-08
+    2.325982249534264e-07
+     5.92445081707473e-07
+ 1.231e+11   
+    5.939514747428587e-07
+    2.327117817345334e-07
+    5.423610152671755e-07
+    4.253259794708635e-08
+    1.580284505032718e-07
+    5.422832426708833e-07
+     3.44737290379659e-09
+    4.253343596060331e-08
+    2.327089580356025e-07
+    5.938487824731747e-07
+ 1.236e+11   
+    5.953635831727242e-07
+    2.328165242832193e-07
+    5.433322716569574e-07
+    4.225460026549214e-08
+    1.583481424338696e-07
+    5.432533131295465e-07
+    3.283943661405661e-09
+    4.225544274712617e-08
+    2.328137683464776e-07
+    5.952598621127702e-07
+ 1.241e+11   
+    5.967831406408742e-07
+    2.329152823834082e-07
+    5.443082724521132e-07
+    4.197634888641949e-08
+    1.586679717779748e-07
+    5.442281114758546e-07
+    3.122219237053418e-09
+    4.197719510604977e-08
+    2.329126050795845e-07
+    5.966783736689821e-07
+ 1.246e+11   
+    5.982102008691384e-07
+    2.330080052365509e-07
+    5.452890552236275e-07
+    4.169789507891765e-08
+     1.58987899973179e-07
+    5.452076751654425e-07
+    2.962164463069386e-09
+    4.169874414158174e-08
+    2.330054176252181e-07
+    5.981043706712737e-07
+ 1.251e+11   
+     5.99644818062907e-07
+    2.330946422331702e-07
+    5.462746580575788e-07
+    4.141929082090767e-08
+    1.593078874863059e-07
+    5.461920421737169e-07
+    2.803741681062067e-09
+    4.142014166187977e-08
+    2.330921555626713e-07
+    5.995379071319657e-07
+ 1.256e+11   
+    6.010870469077276e-07
+    2.331751429432323e-07
+    5.472651195603784e-07
+    4.114058882227164e-08
+    1.596278938169424e-07
+    5.471812510011926e-07
+    2.646910721350572e-09
+    4.114144020234788e-08
+    2.331727686506136e-07
+    6.009790375428489e-07
+ 1.261e+11   
+    6.025369425663777e-07
+    2.332494571043046e-07
+    5.482604788649746e-07
+    4.086184254958319e-08
+    1.599478775007001e-07
+    5.481753406797362e-07
+    2.491628884369252e-09
+    4.086269305064297e-08
+    2.332472068152351e-07
+    6.024278168723375e-07
+ 1.266e+11   
+    6.039945606767787e-07
+    2.333175346075058e-07
+    5.492607756379286e-07
+    4.058310625264738e-08
+    1.602677961118516e-07
+    5.491743507797732e-07
+    2.337850924178249e-09
+    4.058395427341569e-08
+    2.333154201360255e-07
+     6.03884300563239e-07
+ 1.271e+11   
+    6.054599573505137e-07
+      2.3337932548075e-07
+    5.502660500879013e-07
+    4.030443499288246e-08
+    1.605876062654582e-07
+    5.501783214187875e-07
+    2.185529034035563e-09
+    4.030527874504524e-08
+    2.333773588292455e-07
+     6.05348544531461e-07
+ 1.276e+11   
+    6.069331891724323e-07
+    2.334347798694007e-07
+    5.512763429752713e-07
+    4.002588467383349e-08
+    1.609072636184613e-07
+    5.511872932710017e-07
+    2.034612834256363e-09
+    4.002672217844712e-08
+    2.334329732283696e-07
+    6.068206051655028e-07
+ 1.281e+11   
+    6.084143132013007e-07
+    2.334838480138295e-07
+    5.522916956235893e-07
+    3.974751207387998e-08
+    1.612267228699798e-07
+    5.522013075789247e-07
+    1.885049362188813e-09
+     3.97483411580728e-08
+    2.334822137618002e-07
+    6.083005393271231e-07
+ 1.286e+11   
+    6.099033869716631e-07
+    2.335264802238008e-07
+    5.533121499327366e-07
+    3.946937488128384e-08
+    1.615459377599495e-07
+    5.532204061663775e-07
+    1.736783064560079e-09
+    3.947019317538228e-08
+    2.335250309271767e-07
+    6.097884043531854e-07
+ 1.291e+11   
+    6.114004684971462e-07
+    2.335626268492824e-07
+    5.543377483941132e-07
+    3.919153173190691e-08
+    1.618648610664504e-07
+    5.542446314537863e-07
+    1.589755792036671e-09
+    3.919233666687576e-08
+    2.335613752622723e-07
+    6.112842580589239e-07
+ 1.296e+11   
+    6.129056162753725e-07
+     2.33592238247547e-07
+    5.553685341082315e-07
+    3.891404224958294e-08
+    1.621834446010558e-07
+    5.552740264756945e-07
+     1.44390679617833e-09
+    3.891483105494807e-08
+    2.335911973120775e-07
+    6.127881587428331e-07
+ 1.301e+11   
+    6.144188892946412e-07
+    2.336152647459782e-07
+    5.564045508047657e-07
+    3.863696708958003e-08
+    1.625016392018398e-07
+    5.563086349007655e-07
+    1.299172728567653e-09
+    3.863773679171122e-08
+    2.336144475917445e-07
+    6.143001651932805e-07
+ 1.306e+11   
+    6.159403470427242e-07
+    2.336316566006506e-07
+    5.574458428657954e-07
+    3.836036798523889e-08
+     1.62819394724173e-07
+    5.573485010549339e-07
+    1.155487642415545e-09
+    3.836111540613674e-08
+    2.336310765451915e-07
+    6.158203366972273e-07
+ 1.311e+11   
+    6.174700495178609e-07
+    2.336413639499636e-07
+    5.584924553520948e-07
+    3.808430779810256e-08
+    1.631366600281716e-07
+    5.583936699475368e-07
+    1.012782996330288e-09
+    3.808502955468617e-08
+    2.336410344988128e-07
+     6.17348733051174e-07
+ 1.316e+11   
+    6.190080572422883e-07
+    2.336443367630719e-07
+    5.595444340331497e-07
+    3.780885057173322e-08
+    1.634533829630567e-07
+    5.594441873012423e-07
+     8.70987660308436e-10
+    3.780954307563232e-08
+    2.336442716100462e-07
+    6.188854145745641e-07
+ 1.321e+11   
+    6.205544312786653e-07
+    2.336405247828214e-07
+    5.606018254214346e-07
+     3.75340615896658e-08
+    1.637695103475925e-07
+     5.60500099586126e-07
+    7.300279239294891e-10
+    3.753472104753888e-08
+    2.336407378104585e-07
+     6.20430442126119e-07
+ 1.326e+11   
+    6.221092332495499e-07
+    2.336298774626158e-07
+    5.616646768110288e-07
+    3.726000743762693e-08
+     1.64084987946074e-07
+    5.615614540579586e-07
+     5.89827506649594e-10
+    3.726062985210782e-08
+    2.336303827426528e-07
+    6.219838771231321e-07
+ 1.331e+11   
+     6.23672525360317e-07
+    2.336123438966775e-07
+    5.627330363213045e-07
+     3.69867560704621e-08
+    1.643997604395695e-07
+    5.626282988017712e-07
+    4.503075699611869e-10
+    3.698733724171414e-08
+    2.336131556908636e-07
+    6.235457815642918e-07
+ 1.336e+11   
+    6.252443704259788e-07
+     2.33587872743505e-07
+    5.638069529463659e-07
+    3.671437688417107e-08
+    1.647137713916354e-07
+    5.637006827809139e-07
+    3.113867314803401e-10
+    3.671491241202183e-08
+    2.335890055044989e-07
+     6.25116218056285e-07
+ 1.341e+11   
+    6.268248319020521e-07
+     2.33556412141638e-07
+    5.648864766105075e-07
+    3.644294079328078e-08
+    1.650269632077974e-07
+    5.647786558921209e-07
+    1.729810806027803e-10
+    3.644342608012386e-08
+    2.335578805141787e-07
+    6.266952498445038e-07
+ 1.346e+11   
+    6.284139739201958e-07
+    2.335179096174227e-07
+     5.65971658230533e-07
+    3.617252031419001e-08
+     1.65339277088183e-07
+    5.658622690274065e-07
+    3.500419571504026e-11
+    3.617295056848256e-08
+    2.335197284397348e-07
+    6.282829408483751e-07
+ 1.351e+11   
+    6.300118613287214e-07
+    2.334723119840365e-07
+    5.670625497855744e-07
+     3.59031896547523e-08
+    1.656506529726621e-07
+    5.669515741434946e-07
+    -1.02632837495175e-10
+    3.590355989534137e-08
+    2.334744962895644e-07
+    6.298793557017116e-07
+ 1.356e+11   
+    6.316185597387848e-07
+    2.334195652311951e-07
+    5.681592043952403e-07
+    3.563502481069152e-08
+    1.659610294772833e-07
+    5.680466243393225e-07
+   -2.400214066813694e-10
+    3.563532987182679e-08
+     2.33422130250599e-07
+    6.314845597985164e-07
+ 1.361e+11   
+    6.332341355764549e-07
+    2.333596144048018e-07
+    5.692616764067195e-07
+    3.536810366935774e-08
+    1.662703438215989e-07
+     5.69147473942661e-07
+   -3.772553528481109e-10
+    3.536833820652936e-08
+    2.333625755684184e-07
+    6.330986193448185e-07
+ 1.366e+11   
+    6.348586561414994e-07
+    2.332924034758798e-07
+    5.703700214920182e-07
+    3.510250612133691e-08
+      1.6657853174547e-07
+    5.702541786065097e-07
+   -5.144309502358635e-10
+    3.510266461788608e-08
+    2.332957764164884e-07
+    6.347216014170455e-07
+ 1.371e+11   
+    6.364921896732417e-07
+    2.332178751979174e-07
+    5.714842967559225e-07
+    3.483831418051765e-08
+    1.668855274144809e-07
+    5.713667954164498e-07
+   -6.516468861050638e-10
+    3.483839095513566e-08
+     2.33221675754002e-07
+    6.363535740274813e-07
+ 1.376e+11   
+    6.381348054242508e-07
+    2.331359709518746e-07
+    5.726045608560299e-07
+    3.457561211344261e-08
+    1.671912633130503e-07
+    5.724853830098025e-07
+   -7.890042412469708e-10
+    3.457560132842334e-08
+    2.331402151713939e-07
+    6.379946061975336e-07
+ 1.381e+11   
+    6.397865737424883e-07
+    2.330466305779572e-07
+    5.737308741358465e-07
+       3.431448657823e-08
+    1.674956701234639e-07
+    5.736100017077617e-07
+   -9.266064716800373e-10
+    3.431438224872282e-08
+    2.330513347226127e-07
+     6.39644768039393e-07
+ 1.386e+11   
+    6.414475661626347e-07
+    2.329497921931544e-07
+    5.748632987720228e-07
+    3.405502677433035e-08
+    1.677986765901118e-07
+    5.747407136616926e-07
+   -1.064559391870796e-09
+    3.405482277833727e-08
+    2.329549727433338e-07
+    6.413041308468214e-07
+ 1.391e+11   
+    6.431178555073852e-07
+     2.32845391993678e-07
+    5.760018989373239e-07
+    3.379732460348872e-08
+    1.681002093671707e-07
+     5.75877583014909e-07
+   -1.202971160395807e-09
+    3.379701469283946e-08
+    2.328510656539834e-07
+    6.429727671958426e-07
+ 1.396e+11   
+    6.447975159994727e-07
+    2.327333640410928e-07
+    5.771467409803667e-07
+    3.354147484304517e-08
+    1.684001928482074e-07
+    5.770206760812165e-07
+   -1.341952268631716e-09
+    3.354105265518912e-08
+    2.327395477466043e-07
+    6.446507510561416e-07
+ 1.401e+11   
+    6.464866233853791e-07
+    2.326136400311545e-07
+    5.782978936239423e-07
+     3.32875753323148e-08
+    1.686985489763675e-07
+     5.78170061541929e-07
+   -1.481615533238131e-09
+    3.328703440306898e-08
+    2.326203509545159e-07
+    6.463381579140614e-07
+ 1.406e+11   
+    6.481852550715827e-07
+    2.324861490440802e-07
+    5.794554281832846e-07
+    3.303572717322699e-08
+    1.689951970330075e-07
+    5.793258106626794e-07
+   -1.622076093430146e-09
+    3.303506095030775e-08
+    2.324934046034036e-07
+    6.480350649080959e-07
+ 1.411e+11   
+    6.498934902743712e-07
+    2.323508172750574e-07
+    5.806194188062585e-07
+    3.278603494605462e-08
+    1.692900534031922e-07
+    5.804879975319583e-07
+   -1.763451413865667e-09
+    3.278523680355006e-08
+    2.323586351427678e-07
+    6.497415509778542e-07
+ 1.416e+11   
+    6.516114101842813e-07
+    2.322075677435993e-07
+    5.817899427370972e-07
+    3.253860694169207e-08
+    1.695830313160211e-07
+    5.816566993232086e-07
+   -1.905861294261549e-09
+    3.253767019529317e-08
+    2.322159658562805e-07
+    6.514576970275786e-07
+ 1.421e+11   
+    6.533390981462212e-07
+    2.320563199803726e-07
+    5.829670806057736e-07
+    3.229355541132556e-08
+    1.698740405574359e-07
+    5.828319965822932e-07
+   -2.049427886851062e-09
+    3.229247333442647e-08
+    2.320653165497215e-07
+    6.531835861053111e-07
+ 1.426e+11   
+    6.550766398565547e-07
+    2.318969896900536e-07
+    5.841509167452438e-07
+    3.205099683527248e-08
+    1.701629871536144e-07
+     5.84013973542765e-07
+   -2.194275723064084e-09
+    3.204976267571546e-08
+    2.319066032150108e-07
+    6.549193035988793e-07
+ 1.431e+11   
+    6.568241235783219e-07
+    2.317294883885661e-07
+    5.853415395386982e-07
+    3.181105221196111e-08
+    1.704497730221005e-07
+    5.852027184708252e-07
+   -2.340531750476273e-09
+    3.180965920957644e-08
+    2.317397376687026e-07
+    6.566649374499609e-07
+ 1.436e+11   
+    6.585816403759262e-07
+    2.315537230130384e-07
+    5.865390417992992e-07
+    3.157384736889379e-08
+     1.70734295588388e-07
+     5.86398324042895e-07
+   -2.488325382001161e-09
+    3.157228877360099e-08
+    2.315646271633734e-07
+    6.584205783875383e-07
+ 1.441e+11   
+    6.603492843707946e-07
+    2.313695955028469e-07
+    5.877435211851074e-07
+    3.133951329707946e-08
+    1.710164473651024e-07
+    5.876008877578632e-07
+   -2.637788558378653e-09
+    3.133778238763879e-08
+    2.313811739701205e-07
+    6.601863201821885e-07
+ 1.446e+11   
+    6.621271530193689e-07
+    2.311770023497596e-07
+    5.889550806519311e-07
+    3.110818651081022e-08
+     1.71296115490808e-07
+     5.88810512387262e-07
+    -2.78905582621918e-09
+    3.110627661389692e-08
+    2.311892749303218e-07
+    6.619622599226247e-07
+ 1.451e+11   
+    6.639153474150643e-07
+    2.309758341152971e-07
+    5.901738289469771e-07
+    3.088000943448068e-08
+    1.715731812254122e-07
+    5.900273064660616e-07
+   -2.942264432985628e-09
+    3.087791394427326e-08
+    2.309888209747737e-07
+    6.637484983160941e-07
+ 1.456e+11   
+    6.657139726158665e-07
+    2.307659749133644e-07
+      5.9139988114675e-07
+     3.06551308186615e-08
+    1.718475193988088e-07
+    5.912513848272863e-07
+   -3.097554441400233e-09
+    3.065284321659762e-08
+    2.307796966080861e-07
+    6.655451400142809e-07
+ 1.461e+11   
+    6.675231379992813e-07
+    2.305473018557738e-07
+    5.926333592421743e-07
+    3.043370618750271e-08
+    1.721189978092704e-07
+     5.92482869184024e-07
+   -3.255068865077019e-09
+    3.043122006221407e-08
+    2.305617793563339e-07
+    6.673522939664468e-07
+ 1.466e+11   
+    6.693429576464547e-07
+    2.303196844586904e-07
+     5.93874392775062e-07
+    3.021589831976881e-08
+    1.723874765679597e-07
+    5.937218887620474e-07
+   -3.414953828008907e-09
+    3.021320738700444e-08
+    2.303349391755595e-07
+    6.691700738016306e-07
+ 1.471e+11   
+    6.711735507574465e-07
+     2.30082984007368e-07
+    5.951231195291075e-07
+    3.000187776603593e-08
+    1.726528073855269e-07
+    5.949685809872251e-07
+   -3.577358750209916e-09
+    2.999897588841657e-08
+     2.30099037818909e-07
+    6.709985982418409e-07
+ 1.476e+11   
+    6.730150420996462e-07
+    2.298370528769178e-07
+    5.963796862801508e-07
+    2.979182340468394e-08
+    1.729148327967716e-07
+      5.9622309223157e-07
+   -3.742436562265469e-09
+    2.978870461115949e-08
+    2.298539281598339e-07
+    6.728379915482457e-07
+ 1.481e+11   
+    6.748675624914615e-07
+     2.29581733806373e-07
+    5.976442496094318e-07
+    2.958592303945538e-08
+    1.731733853188903e-07
+    5.974855786221675e-07
+   -3.910343951790671e-09
+    2.958258154432062e-08
+    2.295994534688388e-07
+    6.746883840024911e-07
+ 1.486e+11   
+    6.767312493234941e-07
+    2.293168591233737e-07
+    5.989169767847532e-07
+    2.938437404178327e-08
+    1.734282865388733e-07
+    5.987562069178195e-07
+   -4.081241644670686e-09
+    2.938080426294031e-08
+    2.293354466410598e-07
+     6.76549912425372e-07
+ 1.491e+11   
+    6.786062471195527e-07
+    2.290422499166322e-07
+    6.001980467141984e-07
+    2.918738404084155e-08
+    1.736793461249563e-07
+    6.000351554577613e-07
+   -4.255294724520585e-09
+    2.918358061726017e-08
+    2.290617293717822e-07
+    6.784227207351298e-07
+ 1.496e+11   
+    6.804927081398944e-07
+    2.287577151532679e-07
+    6.014876509776448e-07
+    2.899517166496681e-08
+    1.739263607573421e-07
+    6.013226151880153e-07
+   -4.432672993691421e-09
+    2.899112947309109e-08
+    2.287781112770838e-07
+    6.803069605478573e-07
+ 1.501e+11   
+     6.82390793029273e-07
+    2.284630507378058e-07
+    6.027859949412349e-07
+    2.880796733798452e-08
+    1.741691129725483e-07
+    6.026187907703945e-07
+   -4.613551379770992e-09
+    2.880368150685025e-08
+     2.28484388956375e-07
+    6.822027918224666e-07
+ 1.506e+11   
+    6.843006715123705e-07
+    2.281580385097395e-07
+    6.040932989608026e-07
+    2.862601413438713e-08
+     1.74407369915966e-07
+    6.039239017800314e-07
+   -4.798110391233575e-09
+    2.862148005918372e-08
+    2.281803449937027e-07
+    6.841103835529216e-07
+ 1.511e+11   
+    6.862225231394052e-07
+    2.278424451761834e-07
+    6.054097996798551e-07
+     2.84495686972814e-08
+    1.746408819966435e-07
+    6.052381839972943e-07
+   -4.986536626572332e-09
+    2.844478205134725e-08
+    2.278657468945498e-07
+    6.860299145104058e-07
+ 1.516e+11   
+    6.881565380847195e-07
+     2.27516021176296e-07
+    6.067357514287448e-07
+    2.827890222370348e-08
+    1.748693814381209e-07
+    6.065618908003869e-07
+   -5.179023341318339e-09
+    2.827385896843531e-08
+    2.275403459545207e-07
+    6.879615740382741e-07
+ 1.521e+11   
+    6.901029180013264e-07
+    2.271784994736525e-07
+    6.080714277314679e-07
+    2.811430152160652e-08
+    1.750925807190446e-07
+    6.078952946653198e-07
+   -5.375771077626023e-09
+    2.810899791429988e-08
+    2.272038760564062e-07
+    6.899055629027734e-07
+ 1.526e+11   
+    6.920618769344547e-07
+    2.268295942730093e-07
+    6.094171229268744e-07
+    2.795607014352361e-08
+    1.753101708965088e-07
+     6.09238688779953e-07
+   -5.576988361142989e-09
+     2.79505027427715e-08
+    2.268560523918912e-07
+    6.918620942025031e-07
+ 1.531e+11   
+    6.940336422971886e-07
+    2.264689996573793e-07
+    6.107731539120002e-07
+    2.780452960186482e-08
+    1.755218198054825e-07
+    6.105923887796805e-07
+   -5.782892470610382e-09
+    2.779869527037456e-08
+    2.264965701040404e-07
+    6.938313943398049e-07
+ 1.536e+11   
+    6.960184559115692e-07
+    2.260963881416294e-07
+    6.121398620146085e-07
+    2.766002067124945e-08
+    1.757271701267789e-07
+    6.119567346120437e-07
+   -5.993710285447988e-09
+     2.76539165758332e-08
+    2.261251028464383e-07
+    6.958137040572837e-07
+ 1.541e+11   
+    6.980165751183709e-07
+    2.257114091381717e-07
+    6.135176150031785e-07
+    2.752290478333271e-08
+    1.759258373159927e-07
+    6.133320925383009e-07
+   -6.209679217025445e-09
+    2.751652839181298e-08
+    2.257413012551241e-07
+    6.978092795428713e-07
+ 1.546e+11   
+    7.000282739590507e-07
+    2.253136873307111e-07
+    6.149068092425383e-07
+    2.739356552000557e-08
+    1.761174073857451e-07
+    6.147188572804464e-07
+   -6.431048229686301e-09
+    2.738691459493932e-08
+    2.253447913287104e-07
+    6.998183936067117e-07
+ 1.551e+11   
+    7.020538444334024e-07
+    2.249028209514179e-07
+    6.163078720037825e-07
+     2.72724102110186e-08
+    1.763014345327207e-07
+    6.161174543217549e-07
+    -6.65807895759044e-09
+    2.726548279995006e-08
+    2.249351727125895e-07
+     7.01841336933556e-07
+ 1.556e+11   
+    7.040935978364553e-07
+    2.244783799571638e-07
+     6.17721263937396e-07
+    2.715987164229153e-08
+    1.764774386014144e-07
+    6.175283423704243e-07
+   -6.891046923868675e-09
+    2.715266606442614e-08
+    2.245120168824732e-07
+    7.038784194140881e-07
+ 1.561e+11   
+    7.061478661783817e-07
+    2.240399040999492e-07
+    6.191474817188558e-07
+    2.705640988142737e-08
+    1.766449023755817e-07
+    6.189520159951434e-07
+   -7.130242869024127e-09
+    2.704892471052082e-08
+    2.240748652227842e-07
+    7.059299715589828e-07
+ 1.566e+11   
+    7.082170036910526e-07
+    2.235869008868545e-07
+    6.205870608764009e-07
+    2.696251422719069e-08
+    1.768032686885988e-07
+    6.203890084423724e-07
+   -7.375974195110895e-09
+    2.695474827057692e-08
+    2.236232269949885e-07
+    7.079963459993539e-07
+ 1.571e+11   
+     7.10301388425166e-07
+     2.23118843424544e-07
+    6.220405788109561e-07
+    2.687870528984084e-08
+    1.769519373433542e-07
+    6.218398946453759e-07
+   -7.628566533287592e-09
+    2.687065756336784e-08
+    2.231565771910388e-07
+    7.100779190774119e-07
+ 1.576e+11   
+    7.124014239417178e-07
+    2.226351681432862e-07
+    6.235086580183234e-07
+     2.68055372094478e-08
+    1.770902618322439e-07
+    6.233052944350269e-07
+   -7.888365441810039e-09
+    2.679720690837024e-08
+    2.226743542669049e-07
+    7.121750925311806e-07
+ 1.581e+11   
+    7.145175411017688e-07
+    2.221352723952698e-07
+    6.249919695243148e-07
+    2.674360001959747e-08
+    1.772175458474634e-07
+    6.247858759631778e-07
+   -8.155738242177689e-09
+    2.673498648513508e-08
+    2.221759577510157e-07
+    7.142882952771763e-07
+ 1.586e+11   
+    7.166501999584588e-07
+    2.216185119220786e-07
+    6.264912365437733e-07
+    2.669352216368518e-08
+    1.773330395718259e-07
+    6.262823593492855e-07
+   -8.431076000942765e-09
+    2.668462484547194e-08
+    2.216607457224413e-07
+    7.164179852949577e-07
+ 1.591e+11   
+    7.187998917551932e-07
+    2.210841981858122e-07
+    6.280072383743467e-07
+    2.665597317161307e-08
+    1.774359357397156e-07
+    6.277955205615191e-07
+   -8.714795665211032e-09
+    2.664679158565851e-08
+    2.211280321534196e-07
+    7.185646516175214e-07
+ 1.596e+11   
+     7.20967141034064e-07
+    2.205315955585576e-07
+    6.295408145366412e-07
+    2.663166650438741e-08
+    1.775253654580257e-07
+    6.293261955435683e-07
+   -9.007342359405386e-09
+    2.662220018683683e-08
+    2.205770841108392e-07
+    7.207288164314953e-07
+ 1.601e+11   
+    7.231525078583756e-07
+     2.19959918364455e-07
+    6.310928691721932e-07
+    2.662136257435926e-08
+    1.776003937767089e-07
+    6.308752845989056e-07
+   -9.309191851318906e-09
+    2.661161103088593e-08
+       2.200071188111e-07
+    7.229110372910792e-07
+ 1.606e+11   
+    7.253565901533822e-07
+    2.193683277690008e-07
+    6.326643757110205e-07
+    2.662587194896134e-08
+     1.77660014998113e-07
+     6.32443757044054e-07
+   -9.620853195146898e-09
+    2.661583459981055e-08
+    2.194173005228014e-07
+    7.251119094497069e-07
+ 1.611e+11   
+    7.275800261690346e-07
+    2.187559285096357e-07
+    6.342563818206926e-07
+     2.66460587454934e-08
+    1.777031477147525e-07
+    6.340326561428737e-07
+   -9.942871559198266e-09
+    2.663573486631349e-08
+     2.18806737311596e-07
+    7.273320683133222e-07
+ 1.616e+11   
+    7.298234970687426e-07
+    2.181217654620114e-07
+    6.358700146488946e-07
+     2.66828442249093e-08
+    1.777286295647055e-07
+    6.356431043338438e-07
+   -1.027583124570323e-08
+    2.667223288327815e-08
+    2.181744776213765e-07
+    7.295721920191021e-07
+ 1.621e+11   
+    7.320877296479156e-07
+    2.174648200361607e-07
+    6.375064863716411e-07
+    2.673721059194444e-08
+    1.777352116940056e-07
+    6.372763087624031e-07
+   -1.062035890977308e-08
+    2.672631057983179e-08
+    2.175195066861873e-07
+    7.318330041434999e-07
+ 1.626e+11   
+    7.343734991860234e-07
+     2.16784006396655e-07
+    6.391671000589778e-07
+    2.681020500929648e-08
+    1.777215529154963e-07
+    6.389335671302063e-07
+   -1.097712698432637e-08
+    2.679901477134904e-08
+    2.168407427668894e-07
+    7.341152765432173e-07
+ 1.631e+11   
+    7.366816324358241e-07
+    2.160781675009442e-07
+    6.408532558702701e-07
+    2.690294383298459e-08
+    1.776862135536909e-07
+    6.406162738735015e-07
+   -1.134685731708722e-08
+    2.689146139084941e-08
+    2.161370332068111e-07
+    7.364198323327348e-07
+ 1.636e+11   
+     7.39013010753204e-07
+    2.153460709500637e-07
+    6.425664575909795e-07
+     2.70166170759976e-08
+    1.776276489654175e-07
+    6.423259266822623e-07
+   -1.173032502513668e-08
+    2.700483994869872e-08
+    2.154071503006069e-07
+    7.387475490018178e-07
+ 1.641e+11   
+    7.413685733709284e-07
+     2.14586404645879e-07
+    6.443083195222329e-07
+    2.715249310696473e-08
+    1.775442027261527e-07
+    6.440641333715694e-07
+   -1.212836257180117e-08
+    2.714041822738759e-08
+    2.146497869704124e-07
+     7.41099361676268e-07
+ 1.646e+11   
+    7.437493208194566e-07
+    2.137977722490983e-07
+     6.46080573734674e-07
+    2.731192359017196e-08
+    1.774340994727163e-07
+    6.458326191166603e-07
+   -1.254186406943096e-08
+    2.729954721781705e-08
+    2.138635522436153e-07
+    7.434762665249433e-07
+ 1.651e+11   
+    7.461563184975438e-07
+    2.129786884323846e-07
+    6.478850776973239e-07
+    2.749634867287808e-08
+    1.772954373928503e-07
+    6.476332340621897e-07
+   -1.297178981092784e-08
+     2.74836663028432e-08
+    2.130469665265328e-07
+    7.458793243158387e-07
+ 1.656e+11   
+    7.485907003952483e-07
+    2.121275739229805e-07
+    6.497238222914447e-07
+    2.770730242525886e-08
+    1.771261803532914e-07
+    6.494679613159836e-07
+      -1.341917103106e-08
+    2.769430869355005e-08
+      2.1219845666841e-07
+    7.483096641236834e-07
+ 1.661e+11   
+    7.510536729714936e-07
+    2.112427503295265e-07
+    6.515989402192113e-07
+    2.794641853783312e-08
+       1.769241496584e-07
+    6.513389253367046e-07
+   -1.388511489747605e-08
+    2.793310712302324e-08
+    2.113163508104029e-07
+    7.507684871912243e-07
+ 1.666e+11   
+    7.535465191878613e-07
+     2.10322434747782e-07
+    6.535127148155047e-07
+    2.821543628031605e-08
+    1.766870154322265e-07
+    6.532484007238884e-07
+   -1.437080972954089e-08
+    2.820179980151035e-08
+    2.103988730142437e-07
+    7.532570709458003e-07
+ 1.671e+11   
+    7.560706026999773e-07
+    2.093647341404794e-07
+    6.554675892704384e-07
+    2.851620672515209e-08
+    1.764122876178789e-07
+    6.551988214180095e-07
+   -1.487753044106486e-08
+    2.850223663629281e-08
+    2.094441376658179e-07
+    7.557767731724743e-07
+ 1.676e+11   
+    7.586273722069951e-07
+    2.083676394867003e-07
+    6.574661762688655e-07
+    2.885069923803391e-08
+      1.7609730658928e-07
+    6.571927903164996e-07
+   -1.540664420117798e-08
+    2.883638571841921e-08
+    2.084501436489995e-07
+     7.58329036344302e-07
+ 1.681e+11   
+    7.612183659593047e-07
+    2.073290196967721e-07
+    6.595112680514027e-07
+    2.922100823647745e-08
+    1.757392333716549e-07
+    6.592330893105073e-07
+   -1.595961630499022e-08
+    2.920634007742793e-08
+    2.074147682856969e-07
+    7.609153921096586e-07
+ 1.686e+11   
+    7.638452164235241e-07
+    2.062466152891471e-07
+    6.616058469000167e-07
+    2.962936021646826e-08
+    1.753350394686523e-07
+    6.613226897451687e-07
+   -1.653801624337013e-08
+    2.961432470394372e-08
+    2.063357610386121e-07
+     7.63537465935791e-07
+ 1.691e+11   
+    7.665096551031327e-07
+    2.051180318265459e-07
+    6.637530960487994e-07
+    3.007812104556999e-08
+    1.748814962958621e-07
+    6.634647633040901e-07
+   -1.714352395837751e-08
+    3.006270383858018e-08
+    2.052107369738556e-07
+    7.661969819068547e-07
+ 1.696e+11   
+    7.692135175118947e-07
+    2.039407331094435e-07
+    6.659564110183481e-07
+    3.056980351947471e-08
+     1.74375164222612e-07
+    6.656626933164126e-07
+    -1.77779362679158e-08
+    3.055398852396282e-08
+     2.04037169981562e-07
+    7.688957676735944e-07
+ 1.701e+11   
+    7.719587482961455e-07
+    2.027120341260801e-07
+    6.682194113692105e-07
+    3.110707517690205e-08
+    1.738123812261177e-07
+    6.679200864816766e-07
+   -1.844317344025936e-08
+    3.109084441483307e-08
+    2.028123857535532e-07
+    7.716357595507273e-07
+ 1.706e+11   
+    7.747474065005188e-07
+    2.014290937594788e-07
+    6.705459528666344e-07
+    3.169276636591859e-08
+     1.73189251165122e-07
+    6.702407850049673e-07
+   -1.914128589562563e-08
+    3.167609983906744e-08
+    2.015335545185534e-07
+    7.744190077566295e-07
+ 1.711e+11   
+     7.77581670970207e-07
+    2.000889072535452e-07
+    6.729401400452245e-07
+    3.232987855219835e-08
+    1.725016316830624e-07
+    6.726288791306963e-07
+    -1.98744610087838e-08
+    3.231275410021983e-08
+    2.001976835368807e-07
+    7.772476817884616e-07
+ 1.716e+11   
+    7.804638458810408e-07
+    1.986882984420575e-07
+    6.754063391577887e-07
+    3.302159285715979e-08
+    1.717451217545071e-07
+    6.750887200592617e-07
+    -2.06450299831911e-08
+    3.300398600932768e-08
+     1.98801609358506e-07
+    7.801240759240379e-07
+ 1.721e+11   
+    7.833963663867065e-07
+    1.972239117468109e-07
+    6.779491914879622e-07
+    3.377127881108971e-08
+    1.709150488926226e-07
+    6.776249332262234e-07
+   -2.145547476339563e-08
+    3.375316263094804e-08
+    1.973419898505139e-07
+    7.830506148398491e-07
+ 1.726e+11   
+    7.863818043701211e-07
+    1.956922039534887e-07
+    6.805736270008363e-07
+    3.458250330275349e-08
+    1.700064560400944e-07
+    6.802424319182101e-07
+   -2.230843494919328e-08
+    3.456384822486267e-08
+    1.958152960025816e-07
+    7.860298593323257e-07
+ 1.731e+11   
+    7.894228742836046e-07
+    1.940894357771156e-07
+    6.832848782996654e-07
+    3.545903970361184e-08
+    1.690140881709881e-07
+    6.829464311935227e-07
+    -2.32067146712201e-08
+    3.543981336137186e-08
+    1.942178035222121e-07
+    7.890645121271302e-07
+ 1.736e+11   
+    7.925224390596553e-07
+     1.92411663232394e-07
+    6.860884948503227e-07
+     3.64048771404019e-08
+    1.679323786370259e-07
+    6.857424620692572e-07
+    -2.41532893841769e-08
+    3.638504418374484e-08
+    1.925455842348835e-07
+    7.921574237583464e-07
+ 1.741e+11   
+    7.956835160711744e-07
+    1.906547288282165e-07
+    6.889903574274822e-07
+    3.742422988556636e-08
+    1.667554352980725e-07
+     6.88636385928834e-07
+   -2.515131253069773e-08
+    3.740375178709467e-08
+     1.90794497308389e-07
+    7.953115984965911e-07
+ 1.746e+11   
+    7.989092831166272e-07
+    1.888142526104261e-07
+    6.919966927285008e-07
+    3.852154682987238e-08
+    1.654770264839102e-07
+    6.916344090961657e-07
+   -2.620412202536627e-08
+    3.850038167769019e-08
+    1.889601803252475e-07
+    7.985302003017073e-07
+ 1.751e+11   
+    8.022030844021694e-07
+    1.868856230820251e-07
+    6.951140880922192e-07
+    3.970152099634246e-08
+    1.640905668423187e-07
+    6.947430975135977e-07
+   -2.731524650566248e-08
+    3.967962327155229e-08
+    1.870380402323229e-07
+    8.018165587721778e-07
+ 1.756e+11   
+    8.055684364887684e-07
+    1.848639880359618e-07
+    6.983495062500146e-07
+    4.096909904868568e-08
+    1.625891031371769e-07
+    6.979693914513073e-07
+   -2.848841129374985e-08
+    4.094641938508984e-08
+    1.850232442025782e-07
+    8.051741750595392e-07
+ 1.761e+11   
+    8.090090341684876e-07
+    1.827442453422001e-07
+     7.01710300026373e-07
+    4.232949074134269e-08
+    1.609653000697311e-07
+    7.013206201656261e-07
+   -2.972754401076845e-08
+    4.230597566429498e-08
+    1.829107104505454e-07
+    8.086067277120305e-07
+ 1.766e+11   
+     8.12528756229562e-07
+     1.80521033737837e-07
+    7.052042268951354e-07
+    4.378817825143051e-08
+    1.592114262064838e-07
+    7.048045164126089e-07
+   -3.103677978327863e-08
+    4.376376989227724e-08
+    1.806950990501121e-07
+    8.121180784073841e-07
+ 1.771e+11   
+    8.161316710656067e-07
+    1.781887236769845e-07
+    7.088394632859666e-07
+     4.53509253260644e-08
+    1.573193401079259e-07
+    7.084292307120111e-07
+   -3.242046598016278e-08
+    4.532556110778162e-08
+    1.783708028110942e-07
+    8.157122775301196e-07
+ 1.776e+11   
+    8.198220420795371e-07
+    1.757414083054213e-07
+    7.126246185236074e-07
+    4.702378617101777e-08
+    1.552804767640283e-07
+    7.122033452445471e-07
+   -3.388316641722152e-08
+    4.699739845976927e-08
+     1.75931938279418e-07
+    8.193935695441342e-07
+ 1.781e+11   
+    8.236043328281792e-07
+    1.731728946338389e-07
+    7.165687482699676e-07
+    4.881311399899675e-08
+    1.530858344543117e-07
+    7.161358872531522e-07
+   -3.542966496661103e-08
+    4.878562971537453e-08
+    1.733723369345727e-07
+    8.231663981065419e-07
+ 1.786e+11   
+    8.274832118487563e-07
+    1.704766949929702e-07
+    7.206813673265277e-07
+    5.072556914761207e-08
+    1.507259621627386e-07
+    7.202363418065283e-07
+   -3.706496850837927e-08
+    5.069690933019551e-08
+    1.706855366672824e-07
+    8.270354108640164e-07
+ 1.791e+11   
+    8.314635571038547e-07
+    1.676460188630774e-07
+    7.249724616419256e-07
+    5.276812666822061e-08
+    1.481909476901238e-07
+      7.2451466377055e-07
+   -3.879430916283911e-08
+    5.273820598118581e-08
+    1.678647736298108e-07
+    8.310054638681675e-07
+ 1.796e+11   
+    8.355504599769168e-07
+    1.646737651800721e-07
+    7.294524993571857e-07
+    5.494808327679872e-08
+    1.454704066189601e-07
+    7.289812888211717e-07
+   -4.062314574428073e-08
+    5.491680945278163e-08
+    1.649029745609644e-07
+     8.35081625541853e-07
+ 1.801e+11   
+    8.397492287458568e-07
+    1.615525152295995e-07
+    7.341324407091604e-07
+    5.727306354565382e-08
+    1.425534722972684e-07
+    7.336471433204165e-07
+   -4.255716437979553e-08
+    5.724033675593801e-08
+      1.6179274969724e-07
+    8.392691801240142e-07
+ 1.806e+11   
+    8.440653914580858e-07
+    1.582745262493254e-07
+    7.390237466014235e-07
+    5.975102519800274e-08
+    1.394287870185344e-07
+    7.385236528658048e-07
+   -4.460227824125519e-08
+    5.971673734576875e-08
+    1.585263863906901e-07
+    8.435736305162281e-07
+ 1.811e+11   
+    8.485046981254043e-07
+    1.548317258675401e-07
+    7.441383856411847e-07
+    6.239026334213186e-08
+    1.360844945834007e-07
+     7.43622749312685e-07
+   -4.676462634438383e-08
+    6.235429728438579e-08
+    1.550958435626439e-07
+    8.480007004500013e-07
+ 1.816e+11   
+    8.530731221513887e-07
+    1.512157075128063e-07
+     7.49488839430748e-07
+     6.51994134391923e-08
+    1.325082344345155e-07
+    7.489568760577294e-07
+   -4.905057137698255e-08
+    6.516164216567576e-08
+    1.514927471302207e-07
+    8.525563358890829e-07
+ 1.821e+11   
+    8.577768608947818e-07
+    1.474177269346062e-07
+    7.550881058913375e-07
+    6.818745272277943e-08
+    1.286871375574619e-07
+    7.545389913591753e-07
+   -5.146669652937125e-08
+    6.814773856897481e-08
+    1.477083865500624e-07
+    8.572467055746915e-07
+ 1.826e+11   
+    8.626223352560912e-07
+    1.434286999782038e-07
+    7.609497003843186e-07
+    7.136369964594552e-08
+    1.246078243355153e-07
+    7.603825694507376e-07
+   -5.401980131570939e-08
+    7.132189371967467e-08
+    1.437337126314602e-07
+    8.620782006115532e-07
+ 1.831e+11   
+    8.676161881418181e-07
+    1.392392017590986e-07
+    7.670876543747207e-07
+    7.473781065629609e-08
+    1.202564045309261e-07
+    7.665015991738511e-07
+   -5.671689639734479e-08
+     7.46937528701006e-08
+    1.395593367817386e-07
+     8.67057432973554e-07
+ 1.836e+11   
+    8.727652815924929e-07
+    1.348394673851604e-07
+    7.735165113449924e-07
+    7.831977305679123e-08
+    1.156184795350002e-07
+    7.729105797879858e-07
+   -5.956519745304121e-08
+    7.827329360048255e-08
+    1.351755318664493e-07
+    8.721912327698345e-07
+ 1.841e+11   
+     8.78076692214471e-07
+    1.302193943839123e-07
+    7.802513195914675e-07
+    8.211989161670554e-08
+    1.106791469739239e-07
+    7.796245134809872e-07
+   -6.257211819219425e-08
+    8.207081563046762e-08
+    1.305722349102501e-07
+    8.774866440331269e-07
+ 1.846e+11   
+    8.835577042396302e-07
+    1.253685470251623e-07
+    7.873076213770011e-07
+    8.614876436323833e-08
+    1.054230076638201e-07
+     7.86658893801831e-07
+   -6.574526268564758e-08
+    8.609692352845435e-08
+     1.25739051965638e-07
+    8.829509186258536e-07
+ 1.851e+11   
+     8.89215798848808e-07
+     1.20276162829902e-07
+    7.947014375734931e-07
+    9.041723837347644e-08
+    9.983417475805985e-08
+    7.940296885804001e-07
+   -6.909241730311184e-08
+    9.036249730115296e-08
+    1.206652657155936e-07
+     8.88591507506514e-07
+ 1.856e+11   
+    8.950586368987736e-07
+    1.149311618439751e-07
+    8.024492462035059e-07
+    9.493632690685766e-08
+     9.38962847161227e-08
+    8.017533144604842e-07
+   -7.262154268487003e-08
+      9.4878641024348e-08
+    1.153398469348379e-07
+    8.944160478476586e-07
+ 1.861e+11   
+    9.010940290226666e-07
+    1.093221600453223e-07
+     8.10567951766695e-07
+    9.971705043775728e-08
+    8.759250952759246e-08
+    8.098465971097331e-07
+   -7.634076622073174e-08
+    9.965659016268624e-08
+    1.097514722053213e-07
+    9.004323429119323e-07
+ 1.866e+11   
+    9.073298809415979e-07
+    1.034374903600251e-07
+    8.190748391832382e-07
+    1.047701315189637e-07
+    8.090556993531285e-08
+    8.183267052202554e-07
+   -8.025837492048031e-08
+    1.047075406283784e-07
+    1.038885529695424e-07
+    9.066483283807882e-07
+ 1.871e+11   
+    9.137740933124387e-07
+    9.726524004374097e-08
+    8.279875008921277e-07
+    1.101054414734488e-07
+     7.38177522235707e-08
+    8.272110380914762e-07
+    -8.43828053457982e-08
+    1.100423364179146e-07
+    9.773928555582408e-08
+     9.13072013109776e-07
+ 1.876e+11   
+    9.204344014724529e-07
+    9.079332413895754e-08
+     8.37323720682656e-07
+    1.157311971556331e-07
+    6.631094294507074e-08
+    8.365170521977166e-07
+   -8.872261556676759e-08
+    1.156709453405441e-07
+    9.129173357096649e-08
+    9.197113762938789e-07
+ 1.881e+11   
+    9.273182463983024e-07
+     8.40096231563262e-08
+     8.47101314809298e-07
+    1.216536825273382e-07
+    5.836672913793849e-08
+    8.462621145731309e-07
+   -9.328639465513032e-08
+    1.216018225292305e-07
+    8.453392347276542e-08
+     9.26574218619707e-07
+ 1.886e+11   
+    9.344331478727327e-07
+    7.690214372712826e-08
+    8.573380531176134e-07
+    1.278805359638849e-07
+     4.99666452763203e-08
+    8.564638409098742e-07
+   -9.808254610559086e-08
+    1.278421194162506e-07
+    7.745379853822575e-08
+     9.33668091674967e-07
+ 1.891e+11   
+    9.417882144305653e-07
+    6.945884590246722e-08
+    8.680521103361831e-07
+    1.344304102833719e-07
+    4.109247724882816e-08
+    8.671415442596359e-07
+   -1.031190659161936e-07
+     1.34401523740956e-07
+    7.003875906264082e-08
+    9.410007860760945e-07
+ 1.896e+11   
+    9.493951366648265e-07
+     6.16667101684373e-08
+    8.792633969632605e-07
+    1.413364908400771e-07
+     3.17260411155915e-08
+    8.783171962923908e-07
+   -1.084038576853427e-07
+    1.413005525502479e-07
+    6.227518739076295e-08
+     9.48581770637761e-07
+ 1.901e+11   
+    9.572655696205798e-07
+    5.351124826114939e-08
+    8.909939963924309e-07
+    1.486275982421156e-07
+    2.184832824465308e-08
+     8.90012848684725e-07
+   -1.139455481932466e-07
+    1.485706204213071e-07
+    5.414901104954466e-08
+    9.564226987503761e-07
+ 1.906e+11   
+      9.6540860125344e-07
+    4.497790425653486e-08
+    9.032656582477658e-07
+    1.563148912687416e-07
+     1.14393470934055e-08
+    9.022480972922899e-07
+    -1.19753522556027e-07
+    1.562369122421916e-07
+    4.564657433329424e-08
+    9.645348049689719e-07
+ 1.911e+11   
+    9.738318984356201e-07
+    3.605319346862024e-08
+    9.160979231635364e-07
+    1.644020580162084e-07
+    4.789127232215754e-10
+    9.150411704489182e-07
+   -1.258371490028785e-07
+    1.643097700975347e-07
+    3.675471915568593e-08
+    9.729269788069135e-07
+ 1.916e+11   
+    9.825432530395329e-07
+    2.672426180662692e-08
+    9.295091873037154e-07
+    1.728951021962064e-07
+   -1.105282875552107e-08
+    9.284104317320924e-07
+   -1.322053745347131e-07
+    1.727939920708518e-07
+    2.746049602022468e-08
+    9.816069151025023e-07
+ 1.921e+11   
+    9.915509045015817e-07
+    1.697829024940932e-08
+     9.43517927599024e-07
+    1.818035847989234e-07
+     -2.3175406458484e-08
+    9.423746654230577e-07
+   -1.388668165340951e-07
+    1.816964886285685e-07
+    1.775096481091728e-08
+    9.905824221440738e-07
+ 1.926e+11   
+    1.000863364729629e-06
+    6.802359012792865e-09
+    9.581429245121716e-07
+    1.911391387723028e-07
+   -3.590813472500382e-08
+    9.569528652026777e-07
+   -1.458299118003548e-07
+    1.910271569416353e-07
+    7.613160834986454e-09
+    9.998616865503888e-07
+ 1.931e+11   
+    1.010489231913908e-06
+   -3.816480467872668e-09
+    9.734030760400187e-07
+    2.009142642222146e-07
+   -4.927014532205891e-08
+    9.721640140441688e-07
+    -1.53102976689742e-07
+    2.007976374952109e-07
+    -2.96585554593408e-09
+    1.009453116251022e-06
+ 1.936e+11   
+    1.020437074219921e-06
+   -1.489111137731241e-08
+    9.893171986296497e-07
+    2.111416981756057e-07
+   -6.328035910706581e-08
+    9.880269349342892e-07
+   -1.606942099023222e-07
+    2.110202905719502e-07
+   -1.399893322832899e-08
+    1.019365170952356e-06
+ 1.941e+11   
+    1.030715361554273e-06
+   -2.643427653893088e-08
+    1.005903886891299e-06
+    2.218341187821454e-07
+   -7.795743321598432e-08
+    1.004560189743629e-06
+   -1.686116746850641e-07
+    2.217076433243451e-07
+   -2.549877083016532e-08
+    1.029606253444386e-06
+ 1.946e+11   
+    1.041332422024108e-06
+   -3.845852026735747e-08
+    1.023181415992554e-06
+     2.33004004220117e-07
+   -9.331970158209429e-08
+    1.021782002935789e-06
+   -1.768632763859099e-07
+    2.328721211945972e-07
+   -3.747786539248884e-08
+    1.040184644488663e-06
+ 1.951e+11   
+    1.052296410263728e-06
+   -5.097614032985783e-08
+    1.041167667318533e-06
+    2.446635579914262e-07
+   -1.093851153480671e-07
+    1.039710197688343e-06
+   -1.854567404146611e-07
+    2.445259155707984e-07
+   -4.994846716966933e-08
+    1.051108460829105e-06
+ 1.956e+11   
+    1.063615281650801e-06
+   -6.399914581898825e-08
+    1.059880066455539e-06
+    2.568246621591738e-07
+   -1.261711853984289e-07
+     1.05836213887787e-06
+   -1.943995918611503e-07
+    2.566809119669403e-07
+   -6.292253864760016e-08
+    1.062385624683148e-06
+ 1.961e+11   
+    1.075296769815287e-06
+   -7.753921891332307e-08
+      1.0793355284186e-06
+    2.694988425861873e-07
+   -1.436949278470639e-07
+    1.077754680719448e-06
+   -2.036991369401708e-07
+    2.693486446771324e-07
+   -7.641171677835169e-08
+    1.074023839145688e-06
+ 1.966e+11   
+    1.087348366382269e-06
+    -9.16076797013124e-08
+    1.099550408024403e-06
+    2.826972398004124e-07
+   -1.619728129230001e-07
+    1.097904118340987e-06
+   -2.133624462021028e-07
+    2.825402633686311e-07
+   -9.042727801889123e-08
+    1.086030567032131e-06
+ 1.971e+11   
+    1.099777302568439e-06
+    -1.06215453825529e-07
+    1.120540454683944e-06
+    2.964305830957075e-07
+   -1.810207176028374e-07
+    1.118826143209264e-06
+   -2.233963394422866e-07
+    2.962665056277346e-07
+   -1.049801060941856e-07
+    1.098413012125241e-06
+ 1.976e+11   
+    1.112590532543916e-06
+   -1.213730429679885e-07
+    1.142320771487459e-06
+    3.107091671092858e-07
+   -2.008538823130658e-07
+    1.140535802577744e-06
+   -2.338073722768695e-07
+    3.105376731251238e-07
+   -1.200806625677272e-07
+    1.111178102435147e-06
+ 1.981e+11   
+    1.125794718589609e-06
+   -1.370904983041759e-07
+    1.164905778694659e-06
+     3.25542830764442e-07
+   -2.214868720047052e-07
+    1.163047463207271e-06
+   -2.446018243816599e-07
+    3.253636106013359e-07
+   -1.357389603691643e-07
+    1.124332475362493e-06
+ 1.986e+11   
+    1.139396218120016e-06
+   -1.533773970834709e-07
+    1.188309181818747e-06
+    3.409409387001699e-07
+   -2.429335418704616e-07
+    1.186374779612164e-06
+   -2.557856894058925e-07
+    3.407536874964186e-07
+    -1.51964540443249e-07
+    1.137882464769228e-06
+ 1.991e+11   
+    1.153401072644937e-06
+   -1.702428224854165e-07
+    1.212543944491584e-06
+    3.569123653683942e-07
+    -2.65207007930312e-07
+    1.210530667048515e-06
+   -2.673646665768836e-07
+    3.567167822794086e-07
+   -1.687664516700507e-07
+    1.151834089999923e-06
+ 1.996e+11   
+    1.167814998730256e-06
+   -1.876953468734018e-07
+    1.237622266260104e-06
+    3.734654819669533e-07
+   -2.883196226577956e-07
+    1.235527279407998e-06
+   -2.793441540075413e-07
+    3.732612695967371e-07
+   -1.861532341767112e-07
+    1.166193046899737e-06
+ 2.001e+11   
+    1.182643380997053e-06
+    -2.05743018529581e-07
+    1.263555565409992e-06
+    3.906081463357249e-07
+   -3.122829557593733e-07
+    1.261375992118761e-06
+    -2.91729243709571e-07
+    3.903950103510357e-07
+    -2.04132906122754e-07
+    1.180964700861915e-06
+ 2.006e+11   
+     1.19789126717421e-06
+   -2.243933519124175e-07
+    1.290354466851732e-06
+    4.083476958934774e-07
+   -3.371077801562649e-07
+    1.288087390090639e-06
+   -3.045247183028907e-07
+    4.081253447858421e-07
+   -2.227129539987433e-07
+    1.196154081917499e-06
+ 2.011e+11   
+    1.213563365194836e-06
+   -2.436533214341966e-07
+    1.318028795041314e-06
+    4.266909436421009e-07
+    -3.62804063154209e-07
+    1.315671260677529e-06
+   -3.177350493978201e-07
+    4.264590886060613e-07
+   -2.419003264343608e-07
+    1.211765881856751e-06
+ 2.016e+11   
+     1.22966404230235e-06
+   -2.635293587121525e-07
+    1.346587571846297e-06
+    4.456441772162784e-07
+    -3.89380962723822e-07
+    1.344136591567723e-06
+   -3.313643976118628e-07
+    4.454025321170282e-07
+   -2.617014314686313e-07
+    1.227804453348267e-06
+ 2.021e+11   
+    1.246197326109115e-06
+   -2.840273532051261e-07
+    1.376039019209807e-06
+    4.652131609122297e-07
+   -4.168468287543034e-07
+    1.373491573454738e-06
+   -3.454166141683701e-07
+    4.649614423205823e-07
+   -2.821221371936479e-07
+    1.244273810999096e-06
+ 2.026e+11   
+    1.263166907529168e-06
+   -3.051526561086336e-07
+    1.406390566411448e-06
+    4.854031405891968e-07
+   -4.452092090875741e-07
+    1.403743607287702e-06
+   -3.598952440103232e-07
+    4.851410678660853e-07
+     -3.0316777564441e-07
+    1.261177634278143e-06
+ 2.031e+11   
+    1.280576145487582e-06
+    -3.26910087345916e-07
+    1.437648861676133e-06
+    5.062188513023572e-07
+   -4.744748600893033e-07
+     1.43489931585265e-06
+   -3.748035303494908e-07
+    5.059461467186482e-07
+   -3.248431497723507e-07
+    1.278519272206141e-06
+ 2.036e+11   
+    1.298428073292436e-06
+   -3.493039454614748e-07
+    1.469819787840339e-06
+     5.27664527496051e-07
+   -5.046497614691064e-07
+    1.466964559394796e-06
+    -3.90144420559619e-07
+    5.273809163763394e-07
+   -3.471525433092971e-07
+    1.296301749698968e-06
+ 2.041e+11   
+    1.316725406541362e-06
+   -3.723380201971238e-07
+    1.502908481750504e-06
+     5.49743915561312e-07
+   -5.357391350244526e-07
+    1.499944454957246e-06
+   -4.059205733121622e-07
+    5.494491264427343e-07
+   -3.700997333023345e-07
+    1.314527775437121e-06
+ 2.046e+11   
+    1.335470552423384e-06
+   -3.960156075090335e-07
+     1.53691935704052e-06
+    5.724602885419699e-07
+   -5.677474669522783e-07
+    1.533843399084122e-06
+   -4.221343668447311e-07
+    5.721540533409496e-07
+   -3.936880050786287e-07
+    1.333199751122896e-06
+ 2.051e+11   
+    1.354665620268197e-06
+   -4.203395267676779e-07
+    1.571856129914699e-06
+    5.958164627587101e-07
+   -6.006785333490347e-07
+    1.568665093515622e-06
+   -4.387879082458213e-07
+    5.954985169400763e-07
+   -4.179201693829014e-07
+      1.3523197819783e-06
+ 2.056e+11   
+    1.374312433189228e-06
+   -4.453121398710423e-07
+    1.607721847548906e-06
+    6.198148161103568e-07
+   -6.345354285037338e-07
+    1.604412573489064e-06
+   -4.558830436346818e-07
+    6.194848988544614e-07
+   -4.427985814187455e-07
+    1.371889688330814e-06
+ 2.061e+11   
+    1.394412540663477e-06
+   -4.709353719947332e-07
+    1.644518918715724e-06
+    6.444573078059589e-07
+   -6.693205955795641e-07
+    1.641088238253105e-06
+   -4.734213691122716e-07
+    6.441151621704479e-07
+   -4.683251615183718e-07
+     1.39191101813091e-06
+ 2.066e+11   
+    1.414967231890355e-06
+   -4.972107337004705e-07
+    1.682249146238801e-06
+     6.69745499279797e-07
+   -7.050358592770991e-07
+    1.678693883401873e-06
+   -4.914042423581356e-07
+    6.693908723534239e-07
+   -4.945014171633188e-07
+    1.412385060244329e-06
+ 2.071e+11   
+    1.435977549773162e-06
+   -5.241393441266795e-07
+     1.72091376088692e-06
+    6.956805760436843e-07
+   -7.416824600759839e-07
+    1.717230734640972e-06
+   -5.098327947486045e-07
+    6.953132190902771e-07
+   -5.213284660808629e-07
+    1.433312858363564e-06
+ 2.076e+11   
+    1.457444305370395e-06
+   -5.517219549909792e-07
+    1.760513456328709e-06
+    7.222633702368222e-07
+   -7.792610896613401e-07
+    1.756699482607937e-06
+   -5.287079438739237e-07
+    7.218830388279697e-07
+   -5.488070601470533e-07
+    1.454695225386537e-06
+ 2.081e+11   
+    1.479368092669332e-06
+   -5.799589751438797e-07
+    1.801048424784093e-06
+    7.494943836420685e-07
+   -8.177719271554103e-07
+    1.797100318384652e-06
+   -5.480304063354329e-07
+    7.491008377775864e-07
+    -5.76937609836742e-07
+    1.476532758115675e-06
+ 2.086e+11   
+    1.501749303541364e-06
+    -6.08850495425571e-07
+    1.842518393027559e-06
+    7.773738109489565e-07
+   -8.572146757936528e-07
+    1.838432969358345e-06
+   -5.678007107088482e-07
+    7.769668151645099e-07
+    -6.05720208973611e-07
+    1.498825852137531e-06
+ 2.091e+11   
+    1.524588142746737e-06
+   -6.383963135927715e-07
+    1.884922658420652e-06
+    8.059015630572367e-07
+   -8.975885997067136e-07
+    1.880696735110011e-06
+   -5.880192105656467e-07
+    8.054808865188087e-07
+   -6.351546595482085e-07
+    1.521574716751323e-06
+ 2.096e+11   
+    1.547884642865678e-06
+   -6.685959590996156e-07
+    1.928260124675863e-06
+    8.350772902298681e-07
+   -9.388925604946519e-07
+    1.923890523033761e-06
+   -6.086860974514084e-07
+    8.346427068149923e-07
+   -6.652404963889735e-07
+    1.544779389824013e-06
+ 2.101e+11   
+    1.571638679043108e-06
+   -6.994487175351991e-07
+    1.972529337080893e-06
+    8.649004049209049e-07
+   -9.811250533070748e-07
+    1.968012883417307e-06
+   -6.298014137276346e-07
+    8.644516932867902e-07
+   -6.959770114898775e-07
+    1.568439752459656e-06
+ 2.106e+11   
+    1.595849983444806e-06
+   -7.309536545400795e-07
+    2.017728516940161e-06
+    8.953701041210705e-07
+   -1.024284242171487e-06
+    2.013062043741682e-06
+    -6.51365065191725e-07
+    8.949070477598716e-07
+   -7.273632778178357e-07
+    1.592555543381482e-06
+ 2.111e+11   
+    1.620518159334068e-06
+   -7.631096390443122e-07
+    2.063855595019115e-06
+    9.264853910816111e-07
+   -1.068367994341669e-06
+    2.059035941986728e-06
+   -6.733768333983402e-07
+    9.260077783632758e-07
+   -7.593981724433266e-07
+    1.617126372936153e-06
+ 2.116e+11   
+    1.645642694689048e-06
+   -7.959153656901214e-07
+    2.110908243805663e-06
+    9.582450962951489e-07
+   -1.113373913467689e-06
+    2.105932258757668e-06
+   -6.958363876142015e-07
+    9.577527204983109e-07
+    -7.92080398858102e-07
+    1.642151736640926e-06
+ 2.121e+11   
+    1.671222975292334e-06
+   -8.293693763227774e-07
+    2.158883908431452e-06
+    9.906478976300454e-07
+   -1.159299371418752e-06
+    2.153748448076279e-06
+   -7.187432963471905e-07
+    9.901405569615702e-07
+    -8.25408508364195e-07
+    1.667631028205526e-06
+ 2.126e+11   
+    1.697258297235221e-06
+   -8.634700804532043e-07
+     2.20777983612349e-06
+    1.023692339532394e-06
+   -1.206141538618984e-06
+    2.202481766707828e-06
+   -7.420970383994425e-07
+    1.023169837136195e-06
+   -8.593809204383742e-07
+    1.693563551971591e-06
+ 2.131e+11   
+    1.723747878789849e-06
+   -8.982157746150742e-07
+    2.257593104083026e-06
+    1.057376851226525e-06
+   -1.253897412783993e-06
+    2.252129301921377e-06
+   -7.658970134026839e-07
+    1.056838995182337e-06
+   -8.939959419953285e-07
+    1.719948534723104e-06
+ 2.136e+11   
+     1.75069087161261e-06
+   -9.336046605575347e-07
+    2.308320645713898e-06
+    1.091699763861028e-06
+   -1.302563845972561e-06
+    2.302687997606003e-06
+    -7.90142551802379e-07
+    1.091146367173836e-06
+   -9.292517854911288e-07
+    1.746785136831418e-06
+ 2.141e+11   
+    1.778086371251878e-06
+   -9.696348622319607e-07
+    2.359959275146142e-06
+    1.126659326562405e-06
+   -1.352137569892659e-06
+    2.354154678689226e-06
+   -8.148329242652164e-07
+    1.126090207143264e-06
+   -9.651465858257542e-07
+    1.774072462708129e-06
+ 2.146e+11   
+    1.805933426942099e-06
+   -1.006304441547029e-06
+    2.412505710022336e-06
+    1.162253721372427e-06
+   -1.402615219423839e-06
+    2.406526073825274e-06
+   -8.399673504918578e-07
+    1.161668702011378e-06
+   -1.001678416019216e-06
+    1.801809570547921e-06
+ 2.151e+11   
+    1.834231050674602e-06
+   -1.043611412881125e-06
+     2.46595659253408e-06
+    1.198481077058131e-06
+   -1.453993354339224e-06
+    2.459798836340839e-06
+   -8.655450074238725e-07
+    1.197879985389955e-06
+   -1.038845301650524e-06
+    1.829995481351858e-06
+ 2.156e+11   
+    1.862978225543148e-06
+   -1.081553756354348e-06
+    2.520308508714056e-06
+    1.235339481795174e-06
+   -1.506268479229324e-06
+    2.513969563443815e-06
+   -8.915650368402333e-07
+    1.234722150258678e-06
+   -1.076645234061888e-06
+    1.858629187229163e-06
+ 2.161e+11   
+    1.892173913368923e-06
+   -1.120129429874075e-06
+    2.575558006004803e-06
+    1.272826994735411e-06
+   -1.559437061646706e-06
+    2.569034813716154e-06
+   -9.180265523444502e-07
+     1.27219326052697e-06
+   -1.115076182342152e-06
+    1.887709658982194e-06
+ 2.166e+11   
+    1.921817061615914e-06
+   -1.159336379978573e-06
+    2.631701609139568e-06
+    1.310941656479075e-06
+   -1.613495548505636e-06
+    2.624991122926145e-06
+   -9.449286457488173e-07
+    1.310291361501077e-06
+   -1.154136104114018e-06
+    1.917235852985543e-06
+ 2.171e+11   
+    1.951906609612764e-06
+   -1.199172551511956e-06
+    2.688735834382383e-06
+    1.349681498479603e-06
+   -1.668440380783463e-06
+    2.681835018207154e-06
+   -9.722703928667383e-07
+     1.34901448928446e-06
+   -1.193822955158261e-06
+    1.947206717375286e-06
+ 2.176e+11   
+    1.982441494101953e-06
+   -1.239635896171562e-06
+    2.746657202184926e-06
+    1.389044551416211e-06
+   -1.724268006581638e-06
+    2.739563030660174e-06
+   -1.000050858728282e-06
+     1.38836067914656e-06
+   -1.234134697915932e-06
+    1.977621197569134e-06
+ 2.181e+11   
+    2.013420654140826e-06
+   -1.280724379974945e-06
+     2.80546224832591e-06
+     1.42902885257478e-06
+   -1.780974892613079e-06
+    2.798171706445694e-06
+   -1.028269102237483e-06
+    1.428327972900469e-06
+   -1.275069308915625e-06
+    2.008478241141953e-06
+ 2.186e+11   
+    2.044843035382382e-06
+   -1.322435989698881e-06
+     2.86514753360562e-06
+     1.46963245228239e-06
+   -1.838557534190101e-06
+    2.857657616437297e-06
+     -1.0569241802929e-06
+     1.46891442533479e-06
+   -1.316624785178022e-06
+    2.039776802084351e-06
+ 2.191e+11   
+    2.076707593766169e-06
+   -1.364768738346719e-06
+    2.925709652173442e-06
+    1.510853419444399e-06
+   -1.897012463792683e-06
+    2.918017364514438e-06
+   -1.086015151395354e-06
+    1.510118109748597e-06
+   -1.358799149653837e-06
+    2.071515844474654e-06
+ 2.196e+11   
+    2.109013298651652e-06
+   -1.407720669703181e-06
+    2.987145238569875e-06
+    1.552689846235655e-06
+   -1.956336258300996e-06
+    2.979247594575645e-06
+   -1.115541078768591e-06
+    1.551937122640994e-06
+   -1.401590455754042e-06
+    2.103694345596352e-06
+ 2.201e+11   
+    2.141759135427831e-06
+   -1.451289862037737e-06
+    3.049450973567164e-06
+    1.595139851999352e-06
+   -2.016525544979022e-06
+    3.041344996355898e-06
+   -1.145501033020169e-06
+     1.59436958760879e-06
+   -1.444996791033284e-06
+    2.136311298534757e-06
+ 2.206e+11   
+    2.174944107633896e-06
+   -1.495474431018757e-06
+    3.112623588893995e-06
+    1.638201586408176e-06
+   -2.077577006297624e-06
+    3.104306310133285e-06
+   -1.175894094370832e-06
+    1.637413658506884e-06
+   -1.489016280088342e-06
+    2.169365714287388e-06
+ 2.211e+11   
+    2.208567238626081e-06
+   -1.540272531900822e-06
+    3.176659870930018e-06
+    1.681873231942775e-06
+   -2.139487383685893e-06
+    3.168128330410311e-06
+   -1.206719354481307e-06
+    1.681067521926362e-06
+   -1.533647086733847e-06
+    2.202856623423118e-06
+ 2.216e+11   
+    2.242627572826057e-06
+    -1.58568236104729e-06
+    3.241556663455338e-06
+    1.726153005742486e-06
+   -2.202253480299149e-06
+    3.232807908654656e-06
+    -1.23797591790571e-06
+    1.725329399045208e-06
+   -1.578887415516966e-06
+    2.236783077325251e-06
+ 2.221e+11   
+    2.277124176586009e-06
+   -1.631702156849284e-06
+    3.307310869538983e-06
+    1.771039160882672e-06
+   -2.265872162890868e-06
+    3.298341955183003e-06
+   -1.269662903200852e-06
+    1.770197546905941e-06
+   -1.624735512632002e-06
+    2.271144149053414e-06
+ 2.226e+11   
+    2.312056138704762e-06
+   -1.678330200100642e-06
+    3.373919452648024e-06
+    1.816529987131706e-06
+    -2.33034036287341e-06
+    3.364727440269255e-06
+   -1.301779443720293e-06
+    1.815670259173204e-06
+   -1.671189666294121e-06
+    2.305938933858588e-06
+ 2.231e+11   
+    2.347422570628838e-06
+   -1.725564813886723e-06
+    3.441379437056844e-06
+    1.862623811239447e-06
+   -2.395655076650363e-06
+    3.431961394556261e-06
+   -1.334324688121647e-06
+    1.861745866423088e-06
+   -1.718248206629831e-06
+    2.341166549384836e-06
+ 2.236e+11   
+    2.383222606371018e-06
+   -1.773404363042538e-06
+    3.509687907632728e-06
+    1.909318996807003e-06
+   -2.461813365299802e-06
+    3.500040908846911e-06
+   -1.367297800614812e-06
+    1.908422736013997e-06
+   -1.765909505139394e-06
+    2.376826135590214e-06
+ 2.241e+11   
+    2.419455402177908e-06
+   -1.821847253233364e-06
+    3.578842009070888e-06
+    1.956613943785745e-06
+   -2.528812353684632e-06
+     3.56896313334731e-06
+   -1.400697960977971e-06
+     1.95569927158693e-06
+   -1.814171973784025e-06
+    2.412916854418166e-06
+ 2.246e+11   
+    2.456120135976648e-06
+   -1.870891929708146e-06
+    3.648838944648117e-06
+    2.004507087651143e-06
+   -2.596649229062267e-06
+    3.638725276430983e-06
+   -1.434524364367188e-06
+    2.003573912240804e-06
+   -1.863034063747977e-06
+    2.449437889249387e-06
+ 2.251e+11   
+    2.493216006629377e-06
+   -1.920536875773257e-06
+    3.719675974560636e-06
+    2.052996898294688e-06
+    -2.66532123926193e-06
+    3.709324602989287e-06
+   -1.468776220944256e-06
+    2.052045131425988e-06
+   -1.912494263922739e-06
+    2.486388444162581e-06
+ 2.256e+11   
+    2.530742233022639e-06
+   -1.970780611031212e-06
+    3.791350413907735e-06
+     2.10208187867472e-06
+   -2.734825690493957e-06
+    3.780758432429378e-06
+   -1.503452755346313e-06
+    2.101111435596869e-06
+   -1.962551099157766e-06
+    2.523767743031196e-06
+ 2.261e+11   
+    2.568698053017158e-06
+   -2.021621689425853e-06
+    3.863859630378549e-06
+     2.15176056326428e-06
+   -2.805159944850917e-06
+    3.853024136376813e-06
+   -1.538553206019388e-06
+    2.150771362661566e-06
+   -2.013203128318997e-06
+    2.561575028481349e-06
+ 2.266e+11   
+    2.607082722281866e-06
+   -2.073058697132616e-06
+    3.937201041695576e-06
+    2.202031516331679e-06
+   -2.876321417556569e-06
+     3.92611913613608e-06
+   -1.574076824436736e-06
+    2.201023480264429e-06
+   -2.064448942193528e-06
+    2.599809560734787e-06
+ 2.271e+11   
+    2.645895513034466e-06
+   -2.125090250329357e-06
+    4.011372112864197e-06
+    2.252893330086776e-06
+   -2.948307574014063e-06
+      4.0000408999581e-06
+   -1.610022874221529e-06
+    2.251866383934313e-06
+   -2.116287161275744e-06
+    2.638470616358901e-06
+ 2.276e+11   
+    2.685135712709004e-06
+   -2.177714992880391e-06
+    4.086370353273732e-06
+    2.304344622723484e-06
+   -3.021115926700995e-06
+    4.074786940160038e-06
+   -1.646390630192041e-06
+    2.303298695129135e-06
+   -2.168716433467328e-06
+    2.677557486944297e-06
+ 2.281e+11   
+     2.72480262256942e-06
+   -2.230931593963263e-06
+    4.162193313691344e-06
+    2.356384036386346e-06
+   -3.094744031954496e-06
+    4.150354810138479e-06
+   -1.683179377346133e-06
+    2.355319059204528e-06
+   -2.221735431720545e-06
+    2.717069477728671e-06
+ 2.286e+11   
+    2.764895556286491e-06
+   -2.284738745665343e-06
+     4.23883858318684e-06
+    2.409010235086854e-06
+   -3.169189486686048e-06
+    4.226742101313859e-06
+   -1.720388409800597e-06
+    2.407926143332253e-06
+   -2.275342851651636e-06
+    2.757005906184335e-06
+ 2.291e+11   
+    2.805413838493823e-06
+    -2.33913516057414e-06
+     4.31630378602211e-06
+    2.462221902592431e-06
+   -3.244449925061358e-06
+    4.303946440039696e-06
+   -1.758017029699431e-06
+    2.461118634391271e-06
+   -2.329537409148157e-06
+    2.797366100584961e-06
+ 2.296e+11   
+    2.846356803337289e-06
+    -2.39411956938309e-06
+    4.394586578536106e-06
+    2.516017740309054e-06
+   -3.320523015177527e-06
+    4.381965484507355e-06
+   -1.796064546104062e-06
+    2.514895236852468e-06
+    -2.38431783799182e-06
+    2.838149398565861e-06
+ 2.301e+11   
+    2.887723793030675e-06
+   -2.449690718531811e-06
+    4.473684646052388e-06
+    2.570396465176073e-06
+    -3.39740645576583e-06
+    4.460796921673302e-06
+   -1.834530273877101e-06
+    2.569254670675515e-06
+   -2.439682887515687e-06
+    2.879355145690436e-06
+ 2.306e+11   
+    2.929514156429069e-06
+   -2.505847367897641e-06
+    4.553595699833574e-06
+    2.625356807589865e-06
+   -3.475097972945474e-06
+    4.540438464232966e-06
+    -1.87341353257024e-06
+     2.62419566923457e-06
+   -2.495631320312494e-06
+    2.920982694034314e-06
+ 2.311e+11   
+    2.971727247630043e-06
+   -2.562588288552957e-06
+    4.634317474103697e-06
+    2.680897509370816e-06
+   -3.553595317050284e-06
+    4.620887847662144e-06
+   -1.912713645325552e-06
+    2.679716977287245e-06
+   -2.552161910008428e-06
+    2.963031400797134e-06
+ 2.316e+11   
+    3.014362424611569e-06
+   -2.619912260600809e-06
+    4.715847723156828e-06
+    2.737017321786412e-06
+   -3.632896259547566e-06
+    4.702142827344184e-06
+   -1.952429937798526e-06
+    2.735817348999649e-06
+   -2.609273439114813e-06
+    3.005500626950857e-06
+ 2.321e+11   
+    3.057419047914453e-06
+   -2.677818071099503e-06
+    4.798184218567854e-06
+    2.793715003641489e-06
+   -3.712998590065657e-06
+     4.78420117579882e-06
+   -1.992561737110197e-06
+    2.792495546038513e-06
+   -2.666964696968307e-06
+    3.048389735932349e-06
+ 2.326e+11   
+    3.100896479375803e-06
+   -2.736304512084817e-06
+    4.881324746518546e-06
+    2.850989319444871e-06
+   -3.793900113543941e-06
+    4.867060680025606e-06
+   -2.033108370834561e-06
+    2.849750335739663e-06
+   -2.725234477768162e-06
+    3.091698092386688e-06
+ 2.331e+11   
+    3.144794080919174e-06
+   -2.795370378697047e-06
+    4.965267105250039e-06
+    2.908839037660306e-06
+   -3.875598647516937e-06
+    4.950719138973095e-06
+   -2.074069166026748e-06
+    2.907580489360717e-06
+   -2.784081578717736e-06
+    3.135425060966819e-06
+ 2.336e+11   
+    3.189111213406097e-06
+   -2.855014467418604e-06
+    5.050009102650878e-06
+    2.967262929048219e-06
+   -3.958092019541938e-06
+    5.035174361142825e-06
+   -2.115443448296617e-06
+    2.965984780424536e-06
+   -2.843504798275901e-06
+    3.179570005194242e-06
+ 2.341e+11   
+    3.233847235552677e-06
+   -2.915235574426286e-06
+    5.135548553987477e-06
+    3.026259765103311e-06
+   -4.041378064777469e-06
+    5.120424162334935e-06
+   -2.157230540931427e-06
+    3.024961983158423e-06
+   -2.903502934522431e-06
+     3.22413228638431e-06
+ 2.346e+11   
+    3.279001502914178e-06
+   -2.976032494061228e-06
+    5.221883279782403e-06
+    3.085828316592001e-06
+   -4.125454623718122e-06
+    5.206466363540798e-06
+   -2.199429764070755e-06
+    3.084510871033124e-06
+   -2.964074783640374e-06
+    3.269111262639177e-06
+ 2.351e+11   
+    3.324573366939912e-06
+   -3.037404017418491e-06
+    5.309011103844458e-06
+    3.145967352192689e-06
+    -4.21031954008986e-06
+    5.293298788986533e-06
+   -2.242040433936061e-06
+    3.144630215404553e-06
+     -3.0252191385173e-06
+    3.314506287910531e-06
+ 2.356e+11   
+    3.370562174099809e-06
+   -3.099348931056959e-06
+    5.396929851452531e-06
+    3.206675637240605e-06
+   -4.295970658907984e-06
+    5.380919264329536e-06
+   -2.285061862116657e-06
+    3.205318784260022e-06
+   -3.086934787466123e-06
+    3.360316711133622e-06
+ 2.361e+11   
+    3.416967265083693e-06
+   -3.161866015829544e-06
+    5.485637347694563e-06
+    3.267951932578346e-06
+   -4.382405824698942e-06
+    5.469325615009129e-06
+   -2.328493354913354e-06
+    3.266575341070075e-06
+   -3.149220513065429e-06
+    3.406541875433456e-06
+ 2.366e+11   
+    3.463787974073382e-06
+    -3.22495404583265e-06
+    5.575131415961234e-06
+    3.329794993512182e-06
+   -4.469622879885724e-06
+    5.558515664751096e-06
+   -2.372334212740463e-06
+     3.32839864374604e-06
+   -3.212075091118328e-06
+    3.453181117403439e-06
+ 2.371e+11   
+    3.511023628087737e-06
+   -3.288611787473404e-06
+    5.665409876593431e-06
+    3.392203568873816e-06
+   -4.557619663335792e-06
+    5.648487234225186e-06
+   -2.416583729586484e-06
+    3.390787443702908e-06
+    -3.27549728972828e-06
+    3.500233766456397e-06
+ 2.376e+11   
+    3.558673546399719e-06
+   -3.352837998652194e-06
+    5.756470545681277e-06
+    3.455176400186176e-06
+   -4.646394009069074e-06
+    5.739238139853147e-06
+    -2.46124119253326e-06
+    3.453740485026217e-06
+   -3.339485868489485e-06
+    3.547699144247208e-06
+ 2.381e+11   
+    3.606737040024604e-06
+   -3.417631428057754e-06
+    5.848311234011805e-06
+     3.51871222093172e-06
+   -4.735943745123203e-06
+    5.830766192764722e-06
+   -2.506305881333086e-06
+    3.517256503741308e-06
+   -3.404039577789032e-06
+    3.595576564166083e-06
+ 2.386e+11   
+    3.655213411277887e-06
+   -3.482990814571445e-06
+    5.940929746161786e-06
+     3.58280975592088e-06
+   -4.826266692572083e-06
+    5.923069197897836e-06
+   -2.551777068042956e-06
+    3.581334227182723e-06
+   -3.469157158217545e-06
+    3.643865330901092e-06
+ 2.391e+11   
+    3.704101953401237e-06
+   -3.548914886777022e-06
+    6.034323879731516e-06
+    3.647467720758131e-06
+   -4.917360664693511e-06
+    6.016144953238944e-06
+    -2.59765401671476e-06
+    3.645972373461075e-06
+   -3.534837340084584e-06
+    3.692564740068251e-06
+ 2.396e+11   
+     3.75340195025436e-06
+   -3.615402362571735e-06
+    6.128491424714632e-06
+    3.712684821402427e-06
+    -5.00922346628065e-06
+    6.109991249198617e-06
+   -2.643935983139996e-06
+    3.711169651024261e-06
+   -3.601078843034645e-06
+    3.741674077907132e-06
+ 2.401e+11   
+    3.803112676070819e-06
+   -3.682451948874547e-06
+    6.223430162999171e-06
+    3.778459753818962e-06
+   -5.101852893092346e-06
+    6.204605868117604e-06
+   -2.690622214647469e-06
+    3.776924758309903e-06
+   -3.667880375759652e-06
+    3.791192621039911e-06
+ 2.406e+11   
+    3.853233395275125e-06
+   -3.750062341426737e-06
+    6.319137867993952e-06
+    3.844791203718303e-06
+   -5.195246731436027e-06
+    6.299986583897451e-06
+   -2.737711949952049e-06
+    3.843236383485118e-06
+   -3.735240635803166e-06
+    3.841119636291359e-06
+ 2.411e+11   
+    3.903763362358696e-06
+   -3.818232224680239e-06
+    6.415612304374766e-06
+    3.911677846379286e-06
+   -5.289402757877448e-06
+    6.396131161750206e-06
+   -2.785204419052537e-06
+    3.910103204269954e-06
+   -3.803158309451683e-06
+    3.891454380567224e-06
+ 2.416e+11   
+    3.954701821811983e-06
+   -3.886960271768861e-06
+    6.512851227944292e-06
+    3.979118346551614e-06
+    -5.38431873907085e-06
+    6.493037358061162e-06
+   -2.833098843176595e-06
+     3.97752388784049e-06
+   -3.871632071708239e-06
+    3.942196100788393e-06
+ 2.421e+11   
+    4.006048008109795e-06
+   -3.956245144557274e-06
+    6.610852385599288e-06
+    4.047111358433922e-06
+    -5.47999243170289e-06
+    6.590702920358262e-06
+   -2.881394434770392e-06
+    4.045497090807343e-06
+   -3.940660586343247e-06
+    3.993344033877942e-06
+ 2.426e+11   
+    4.057801145747132e-06
+   -4.026085493762978e-06
+    6.709613515399147e-06
+    4.115655525723186e-06
+   -5.576421582543942e-06
+    6.689125587382201e-06
+   -2.930090397530769e-06
+    4.114021459265429e-06
+   -4.010242506017712e-06
+    4.044897406798254e-06
+ 2.431e+11   
+    4.109960449322384e-06
+   -4.096479959145997e-06
+     6.80913234672899e-06
+    4.184749481731025e-06
+   -5.673603928599761e-06
+    6.788303089250477e-06
+   -2.979185926477439e-06
+    4.183095628910607e-06
+   -4.080376472473738e-06
+    4.096855436635215e-06
+ 2.436e+11   
+    4.162525123665065e-06
+   -4.167427169761474e-06
+    6.909406600551169e-06
+    4.254391849562695e-06
+   -5.771537197357102e-06
+     6.88823314770937e-06
+   -3.028680208062915e-06
+    4.252718225218935e-06
+   -4.151061116787447e-06
+    4.149217330726603e-06
+ 2.441e+11   
+     4.21549436400497e-06
+   -4.238925744270122e-06
+    7.010433989738626e-06
+     4.32458124235427e-06
+   -5.870219107116226e-06
+    6.988913476467178e-06
+   -3.078572420317609e-06
+    4.322887863684087e-06
+   -4.222295059679297e-06
+    4.201982286831631e-06
+ 2.446e+11   
+    4.268867356179766e-06
+   -4.310974291301572e-06
+    7.112212219483664e-06
+    4.395316263563741e-06
+    -5.96964736740379e-06
+    7.090341781602458e-06
+   -3.128861733027655e-06
+    4.393603150108592e-06
+   -4.294076911876917e-06
+    4.255149493338578e-06
+ 2.451e+11   
+    4.322643276878104e-06
+   -4.383571409865988e-06
+    7.214738987776024e-06
+    4.466595507311713e-06
+   -6.069819679459483e-06
+    7.192515762041079e-06
+     -3.1795473079431e-06
+    4.464862680944734e-06
+    -4.36640527452584e-06
+    4.308718129507752e-06
+ 2.456e+11   
+    4.376821293915189e-06
+   -4.456715689809022e-06
+     7.31801198594381e-06
+    4.538417558767427e-06
+   -6.170733736789797e-06
+     7.29543311009576e-06
+   -3.230628299013831e-06
+    4.536665043680601e-06
+   -4.439278739643226e-06
+    4.362687365746611e-06
+ 2.461e+11   
+    4.431400566537926e-06
+   -4.530405712305661e-06
+    7.422028899251278e-06
+    4.610780994575854e-06
+    -6.27238722578254e-06
+    7.399091512062081e-06
+   -3.282103852650945e-06
+    4.609008817267298e-06
+   -4.512695890610165e-06
+    4.417056363914268e-06
+ 2.466e+11   
+    4.486380245756848e-06
+   -4.604640050388521e-06
+    7.526787407547634e-06
+    4.683684383321934e-06
+   -6.374777826376006e-06
+    7.503488648865158e-06
+    -3.33397310801115e-06
+    4.681892572583175e-06
+   -4.586655302698157e-06
+    4.471824277652547e-06
+ 2.471e+11   
+     4.54175947470189e-06
+   -4.679417269506182e-06
+    7.632285185960839e-06
+    4.757126286027734e-06
+   -6.477903212776444e-06
+    7.608622196751025e-06
+   -3.386235197301817e-06
+    4.755314872931032e-06
+   -4.661155543625414e-06
+    4.526990252740744e-06
+ 2.476e+11   
+    4.597537388999401e-06
+    -4.75473592810748e-06
+    7.738519905630909e-06
+    4.831105256678769e-06
+   -6.581761054218101e-06
+    7.714489828017256e-06
+   -3.438889246104386e-06
+    4.829274274564374e-06
+   -4.736195174138822e-06
+    4.582553427471369e-06
+ 2.481e+11   
+    4.653713117167658e-06
+   -4.830594578247752e-06
+    7.845489234477315e-06
+    4.905619842775694e-06
+   -6.686349015760112e-06
+     7.82108921177748e-06
+   -3.491934373713962e-06
+    4.903769327239087e-06
+   -4.811772748617792e-06
+    4.638512933044363e-06
+ 2.486e+11   
+    4.710285781028358e-06
+   -4.906991766213223e-06
+    7.953190837995156e-06
+    4.980668585907656e-06
+     -6.7916647591146e-06
+    7.928418014754336e-06
+   -3.545369693492841e-06
+    4.978798574786689e-06
+   -4.887886815695929e-06
+    4.694867893977042e-06
+ 2.491e+11   
+    4.767254496131579e-06
+   -4.983926033159786e-06
+    8.061622380075028e-06
+    5.056250022343823e-06
+   -6.897705943500791e-06
+    8.036473902096107e-06
+   -3.599194313235932e-06
+    5.054360555705826e-06
+   -4.964535918897136e-06
+    4.751617428527482e-06
+ 2.496e+11   
+    4.824618372191829e-06
+   -5.061395915762822e-06
+    8.170781523841883e-06
+    5.132362683639701e-06
+   -7.004470226520005e-06
+    8.145254538212116e-06
+   -3.653407335545995e-06
+    5.130453803768439e-06
+   -5.041718597282499e-06
+    4.808760649128833e-06
+ 2.501e+11   
+     4.88237651353293e-06
+   -5.139399946874694e-06
+    8.280665932508234e-06
+    5.209005097255042e-06
+   -7.111955265046717e-06
+    8.254757587622322e-06
+   -3.708007858216828e-06
+    5.207076848637583e-06
+   -5.119433386104843e-06
+     4.86629666283242e-06
+ 2.506e+11   
+    4.940528019539453e-06
+   -5.217936656186726e-06
+    8.391273270237142e-06
+     5.28617578718014e-06
+   -7.220158716130914e-06
+    8.364980715816643e-06
+   -3.762994974622435e-06
+    5.284228216493597e-06
+   -5.197678817467678e-06
+    4.924224571757312e-06
+ 2.511e+11   
+    4.999071985112684e-06
+   -5.297004570892795e-06
+    8.502601203010987e-06
+    5.363873274567647e-06
+   -7.329078237907468e-06
+    8.475921590120038e-06
+   -3.818367774110445e-06
+    5.361906430665787e-06
+   -5.276453420985724e-06
+    4.982543473544384e-06
+ 2.516e+11   
+    5.058007501129159e-06
+   -5.376602216351752e-06
+    8.614647399502055e-06
+    5.442096078367118e-06
+   -7.438711490508324e-06
+    8.587577880559237e-06
+   -3.874125342398098e-06
+    5.440110012266851e-06
+   -5.355755724444249e-06
+    5.041252461812878e-06
+ 2.521e+11   
+    5.117333654899741e-06
+   -5.456728116745992e-06
+     8.72740953194109e-06
+    5.520842715959593e-06
+   -7.549056136973489e-06
+    8.699947260727541e-06
+   -3.930266761969117e-06
+    5.518837480827265e-06
+   -5.435584254454522e-06
+    5.100350626617526e-06
+ 2.526e+11   
+    5.177049530627623e-06
+   -5.537380795733765e-06
+    8.840885276980247e-06
+    5.600111703789609e-06
+   -7.660109844157019e-06
+    8.813027408643941e-06
+   -3.986791112469975e-06
+    5.598087354927245e-06
+   -5.515937537103079e-06
+    5.159837054904527e-06
+ 2.531e+11   
+    5.237154209863444e-06
+   -5.618558777093064e-06
+    8.955072316547495e-06
+    5.679901557992588e-06
+    -7.77187028362486e-06
+    8.926816007603751e-06
+   -4.043697471104115e-06
+    5.677858152823902e-06
+   -5.596814098592515e-06
+    5.219710830964704e-06
+ 2.536e+11   
+    5.297646771956003e-06
+   -5.700260585354747e-06
+    9.069968338688794e-06
+     5.76021079501498e-06
+   -7.884335132540699e-06
+    9.041310747017035e-06
+     -4.1009849130227e-06
+    5.758148393071295e-06
+   -5.678212465871654e-06
+    5.279971036882204e-06
+ 2.541e+11   
+    5.358526294497066e-06
+   -5.782484746423224e-06
+    9.185571038395783e-06
+    5.841037932225408e-06
+   -7.997502074537319e-06
+    9.156509323232552e-06
+   -4.158652511710694e-06
+    5.838956595131429e-06
+    -5.76013116725325e-06
+    5.340616752977354e-06
+ 2.546e+11   
+    5.419791853758866e-06
+   -5.865229788182654e-06
+    9.301878118415722e-06
+    5.922381488514711e-06
+   -8.111368800570167e-06
+    9.272409440344176e-06
+   -4.216699339366985e-06
+    5.920281279974161e-06
+   -5.842568733017343e-06
+    5.401647058242217e-06
+ 2.551e+11   
+    5.481442525123028e-06
+   -5.948494241087225e-06
+    9.418887290041723e-06
+    6.004239984883182e-06
+   -8.225933009750849e-06
+    9.389008810977517e-06
+   -4.275124467277513e-06
+    6.002120970664299e-06
+   -5.925523695998759e-06
+    5.463061030767655e-06
+ 2.556e+11   
+    5.543477383499758e-06
+   -6.032276638733886e-06
+    9.536596273880624e-06
+    6.086611945013255e-06
+   -8.341192410157806e-06
+     9.50630515705436e-06
+   -4.333926966180327e-06
+    6.084474192934201e-06
+    -6.00899459215713e-06
+    5.524857748160624e-06
+ 2.561e+11   
+    5.605895503736103e-06
+   -6.116575518416179e-06
+    9.655002800596533e-06
+     6.16949589582617e-06
+   -8.457144719622163e-06
+    9.624296210532935e-06
+   -4.393105906621544e-06
+    6.167339475740289e-06
+   -6.092979961128169e-06
+    5.587036287950663e-06
+ 2.566e+11   
+     5.66869596101235e-06
+   -6.201389421658048e-06
+    9.774104611628196e-06
+    6.252890368021209e-06
+    -8.57378766648657e-06
+    9.742979714122081e-06
+   -4.452660359301496e-06
+    6.250715351802205e-06
+   -6.177478346755008e-06
+     5.64959572798458e-06
+ 2.571e+11   
+    5.731877831225638e-06
+   -6.286716894726421e-06
+    9.893899459878388e-06
+    6.336793896596205e-06
+   -8.691118990335285e-06
+    9.862353421967556e-06
+   -4.512589395410064e-06
+    6.334600358123221e-06
+   -6.262488297598425e-06
+    5.712535146808376e-06
+ 2.576e+11   
+    5.795440191359875e-06
+   -6.372556489121618e-06
+    1.001438511037374e-05
+    6.421205021348126e-06
+   -8.809136442693645e-06
+    9.982415100308969e-06
+   -4.572892086950569e-06
+    6.418993036490737e-06
+   -6.348008367425058e-06
+    5.775853624035595e-06
+ 2.581e+11   
+    5.859382119841299e-06
+   -6.458906762044828e-06
+    1.013555934089372e-05
+    6.506122287352807e-06
+   -8.927837787695661e-06
+      1.0103162528106e-05
+   -4.633567507051543e-06
+    6.503891933955954e-06
+   -6.434037115672779e-06
+     5.83955024070138e-06
+ 2.586e+11   
+    5.923702696878913e-06
+   -6.545766276841746e-06
+    1.025741994256738e-05
+    6.591544245422735e-06
+   -9.047220802718106e-06
+    1.022459349763255e-05
+   -4.694614730265726e-06
+    6.589295603291582e-06
+   -6.520573107892415e-06
+    5.903624079601479e-06
+ 2.591e+11   
+    5.988401004789245e-06
+   -6.633133603421878e-06
+    1.037996472043691e-05
+    6.677469452542172e-06
+   -9.167283278980165e-06
+    1.034670581503787e-05
+   -4.756032832855782e-06
+    6.675202603426926e-06
+   -6.607614916165242e-06
+    5.968074225615675e-06
+ 2.596e+11   
+    6.053476128304904e-06
+   -6.721007318652986e-06
+    1.050319149398705e-05
+    6.763896472278884e-06
+   -9.288023022107532e-06
+    1.046949730087373e-05
+   -4.817820893066296e-06
+    6.761611499859582e-06
+   -6.695161119495779e-06
+     6.03289976601512e-06
+ 2.601e+11   
+    6.118927154866405e-06
+   -6.809386006730063e-06
+    1.062709809763945e-05
+    6.850823875171744e-06
+   -9.409437852659921e-06
+    1.059296579058667e-05
+   -4.879977991381517e-06
+    6.848520865043008e-06
+   -6.783210304179284e-06
+    6.098099790752994e-06
+ 2.606e+11   
+    6.184753174896991e-06
+   -6.898268259518795e-06
+     1.07516823812115e-05
+    6.938250239093808e-06
+   -9.531525606621539e-06
+    1.071710913497494e-05
+   -4.942503210768642e-06
+      6.9359292787496e-06
+   -6.871761064143832e-06
+    6.163673392738294e-06
+ 2.611e+11   
+    6.250953282059955e-06
+   -6.987652676872903e-06
+    1.087694221033882e-05
+    7.026174149590286e-06
+   -9.654284135853586e-06
+    1.084192520060932e-05
+   -5.005395636906171e-06
+    7.023835328408682e-06
+   -6.960812001266495e-06
+     6.22961966809222e-06
+ 2.616e+11   
+    6.317526573498362e-06
+    -7.07753786692551e-06
+    1.100287546686136e-05
+    7.114594200191172e-06
+   -9.777711308508561e-06
+    1.096741187021762e-05
+    -5.06865435839723e-06
+    7.112237609419116e-06
+   -7.050361725663653e-06
+    6.295937716387029e-06
+ 2.621e+11   
+    6.384472150056824e-06
+   -7.167922446354234e-06
+    1.112948004917243e-05
+    7.203508992698133e-06
+   -9.901805009405855e-06
+    1.109356704303244e-05
+   -5.132278466967533e-06
+    7.201134725436268e-06
+    -7.14040885595519e-06
+    6.362626640867092e-06
+ 2.626e+11   
+    6.451789116485219e-06
+   -7.258805040619996e-06
+    1.125675387253061e-05
+    7.292917137445494e-06
+   -1.002656314036836e-05
+     1.12203886351019e-05
+   -5.196267057647875e-06
+    7.290525288633012e-06
+   -7.230952019502579e-06
+    6.429685548651964e-06
+ 2.631e+11   
+    6.519476581624246e-06
+   -7.350184284179677e-06
+    1.138469486933463e-05
+    7.382817253535197e-06
+   -1.015198362052007e-05
+    1.134787457956353e-05
+   -5.260619228941053e-06
+     7.38040791993475e-06
+   -7.321989852620932e-06
+    6.497113550921414e-06
+ 2.636e+11   
+    6.587533658572775e-06
+   -7.442058820672645e-06
+    1.151330098936081e-05
+    7.473207969045673e-06
+    -1.02780643865445e-05
+    1.147602282688103e-05
+   -5.325334082973125e-06
+    7.470781249228358e-06
+   -7.413521000765118e-06
+    6.564909763082351e-06
+ 2.641e+11   
+    6.655959464836882e-06
+   -7.534427303081288e-06
+    1.164257019996349e-05
+     7.56408792121448e-06
+   -1.040480339290393e-05
+    1.160483134504397e-05
+   -5.390410725628907e-06
+    7.561643915544928e-06
+   -7.505544118689966e-06
+    6.633073304917502e-06
+ 2.646e+11   
+    6.724753122460758e-06
+   -7.627288393865839e-06
+    1.177250048623843e-05
+    7.655455756595045e-06
+   -1.053219861201989e-05
+    1.173429811973097e-05
+   -5.455848266671869e-06
+    7.652994567216575e-06
+   -7.598057870584985e-06
+    6.701603300716135e-06
+ 2.651e+11   
+    6.793913758139341e-06
+   -7.720640765073654e-06
+    1.190308985114955e-05
+    7.747310131187267e-06
+    -1.06602480344146e-05
+    1.186442115443603e-05
+   -5.521645819848265e-06
+    7.744831862007179e-06
+   -7.691060930183621e-06
+     6.77049887938656e-06
+ 2.656e+11   
+    6.863440503312987e-06
+   -7.814483098423329e-06
+     1.20343363156191e-05
+     7.83964971054241e-06
+   -1.078894966881418e-05
+    1.199519847055883e-05
+   -5.587802502975701e-06
+    7.837154467217368e-06
+   -7.784551980847506e-06
+    6.839759174550767e-06
+ 2.661e+11   
+    6.933332494244164e-06
+   -7.908814085363936e-06
+     1.21662379185819e-05
+    7.932473169842356e-06
+   -1.091830154221357e-05
+    1.212662810745906e-05
+   -5.654317438016211e-06
+    7.929961059763948e-06
+   -7.878529715625989e-06
+    6.909383324621219e-06
+ 2.666e+11   
+    7.003588872076432e-06
+   -8.003632427109819e-06
+    1.229879271700404e-05
+    8.025779193953538e-06
+   -1.104830169990389e-05
+    1.225870812247537e-05
+   -5.721189751133925e-06
+     8.02325032623395e-06
+   -7.972992837291309e-06
+    6.979370472860009e-06
+ 2.671e+11   
+    7.074208782875838e-06
+    -8.09893683465126e-06
+    1.243199878586625e-05
+     8.11956647745576e-06
+   -1.117894820546246e-05
+    1.239143659090932e-05
+    -5.78841857273751e-06
+    8.117020962913612e-06
+   -8.067940058349807e-06
+    7.049719767420501e-06
+ 2.676e+11   
+    7.145191377654981e-06
+   -8.194726028741546e-06
+    1.256585421811287e-05
+    8.213833724646318e-06
+   -1.131023914070624e-05
+    1.252481160597499e-05
+   -5.856003037507555e-06
+    8.211271675792672e-06
+   -8.163370101029667e-06
+    7.120430361371793e-06
+ 2.681e+11   
+    7.216535812380005e-06
+   -8.290998739860901e-06
+    1.270035712456683e-05
+    8.308579649519744e-06
+   -1.144217260560915e-05
+     1.26588312787148e-05
+   -5.923942284409089e-06
+    8.306001180544299e-06
+   -8.259281697245627e-06
+    7.191501412706181e-06
+ 2.686e+11   
+    7.288241247960811e-06
+   -8.387753708157772e-06
+    1.283550563381134e-05
+    8.403802975723604e-06
+   -1.157474671818398e-05
+    1.279349373788208e-05
+   -5.992235456689462e-06
+    8.401208202481043e-06
+   -8.355673588541097e-06
+    7.262932084329863e-06
+ 2.691e+11   
+    7.360306850224654e-06
+   -8.484989683367822e-06
+    1.297129789203872e-05
+    8.499502436490668e-06
+   -1.170795961432942e-05
+    1.292879712979121e-05
+   -6.060881701861756e-06
+    8.496891476487223e-06
+    -8.45254452600828e-06
+    7.334721544037246e-06
+ 2.696e+11   
+    7.432731789873698e-06
+   -8.582705424711568e-06
+    1.310773206286764e-05
+     8.59567677454807e-06
+    -1.18418094476432e-05
+    1.306473961813596e-05
+   -6.129880171674146e-06
+    8.593049746928311e-06
+   -8.549893270186805e-06
+    7.406868964469158e-06
+ 2.701e+11   
+    7.505515242426517e-06
+   -8.680899700770709e-06
+    1.324480632712881e-05
+    8.692324742003817e-06
+   -1.197629438920184e-05
+    1.320131938377678e-05
+    -6.19923002206522e-06
+    8.689681767537625e-06
+   -8.647718590941358e-06
+    7.479373523055204e-06
+ 2.706e+11   
+    7.578656388144218e-06
+    -8.77957128934409e-06
+    1.338251888262047e-05
+    8.789445100211152e-06
+   -1.211141262730787e-05
+    1.333853462449781e-05
+   -6.268930413105773e-06
+    8.786786301280895e-06
+   -8.746019267318917e-06
+     7.55223440194072e-06
+ 2.711e+11   
+    7.652154411941264e-06
+   -8.878718977283719e-06
+    1.352086794383419e-05
+    8.887036619611297e-06
+   -1.224716236720537e-05
+    1.347638355473427e-05
+   -6.338980508927243e-06
+    8.884362120199297e-06
+   -8.844794087386193e-06
+    7.625450787898598e-06
+ 2.716e+11   
+    7.726008503281582e-06
+   -8.978341560311445e-06
+    1.365985174165182e-05
+    8.985098079555184e-06
+   -1.238354183076466e-05
+    1.361486440527141e-05
+   -6.409379477637116e-06
+    8.982408005231358e-06
+   -8.944041848047804e-06
+    7.699021872226405e-06
+ 2.721e+11   
+    7.800217856060211e-06
+   -9.078437842816863e-06
+    1.379946852301444e-05
+    9.083628268104573e-06
+   -1.252054925613691e-05
+    1.375397542291541e-05
+   -6.480126491221583e-06
+    9.080922746014316e-06
+   -9.043761354845789e-06
+    7.772946850629108e-06
+ 2.726e+11   
+    7.874781668470885e-06
+   -9.179006637637159e-06
+    1.393971655056433e-05
+    9.182625981813236e-06
+   -1.265818289737963e-05
+    1.389371487013729e-05
+   -6.551220725435872e-06
+    9.179905140665578e-06
+   -9.143951421741067e-06
+    7.847224923087885e-06
+ 2.731e+11   
+    7.949699142860026e-06
+   -9.280046765819311e-06
+    1.408059410226043e-05
+    9.282090025488695e-06
+   -1.279644102405389e-05
+    1.403408102469072e-05
+   -6.622661359682413e-06
+      9.2793539955447e-06
+    -9.24461087087742e-06
+    7.921855293715291e-06
+ 2.736e+11   
+    8.024969485567451e-06
+   -9.381557056365483e-06
+    1.422209947096867e-05
+    9.382019211935202e-06
+   -1.293532192079419e-05
+    1.417507217920455e-05
+   -6.694447576877344e-06
+    9.379268124996611e-06
+    -9.34573853232866e-06
+    7.996837170597285e-06
+ 2.741e+11   
+    8.100591906754251e-06
+   -9.483536345961919e-06
+    1.436423096402745e-05
+    9.482412361678351e-06
+   -1.307482388685174e-05
+    1.431668664075075e-05
+   -6.766578563305531e-06
+    9.479646351076495e-06
+   -9.447333243829451e-06
+     8.07216976562246e-06
+ 2.746e+11   
+    8.176565620218281e-06
+   -9.585983478692345e-06
+    1.450698690278986e-05
+    9.583268302672195e-06
+   -1.321494523561244e-05
+    1.445892273038913e-05
+   -6.839053508464606e-06
+    9.580487503257143e-06
+    -9.54939385049059e-06
+    8.147852294298945e-06
+ 2.751e+11   
+     8.25288984319758e-06
+   -9.688897305736063e-06
+     1.46503656221428e-05
+    9.684585869989129e-06
+   -1.335568429408992e-05
+    1.460177878268902e-05
+   -6.911871604898197e-06
+    9.681790418119129e-06
+   -9.651919204499112e-06
+    8.223883975559255e-06
+ 2.756e+11   
+    8.329563796162227e-06
+   -9.792276685051622e-06
+    1.479436547000448e-05
+    9.786363905493391e-06
+   -1.349703940239507e-05
+    1.474525314522945e-05
+   -6.985032048018835e-06
+    9.783553939024593e-06
+   -9.754908164804049e-06
+    8.300264031553679e-06
+ 2.761e+11   
+    8.406586702595014e-06
+   -9.896120481046641e-06
+    1.493898480680086e-05
+    9.888601257498746e-06
+   -1.363900891318278e-05
+     1.48893441780784e-05
+   -7.058534035920846e-06
+    9.885776915775153e-06
+   -9.858359596788284e-06
+    8.376991687432534e-06
+ 2.766e+11   
+    8.483957788761339e-06
+   -1.000042756423416e-05
+    1.508422200492192e-05
+    9.991296780410761e-06
+   -1.378159119107662e-05
+    1.503405025325185e-05
+   -7.132376769183475e-06
+    9.988458204254458e-06
+   -9.962272371927069e-06
+    8.454066171117577e-06
+ 2.771e+11   
+    8.561676283468743e-06
+   -1.010519681087638e-05
+     1.52300754481588e-05
+    1.009444933435447e-05
+   -1.392478461207271e-05
+    1.517936975415386e-05
+   -7.206559450664752e-06
+    1.009159666605617e-05
+     -1.0066645367434e-05
+    8.531486713063253e-06
+ 2.776e+11   
+    8.639741417816513e-06
+   -1.021042710261631e-05
+     1.53765435311227e-05
+    1.019805778478797e-05
+   -1.406858756292357e-05
+    1.532530107499837e-05
+    -7.28108128528633e-06
+     1.01951911680978e-05
+   -1.017147746589475e-05
+    8.609252546007949e-06
+ 2.781e+11   
+    8.718152424935765e-06
+   -1.031611732609768e-05
+    1.552362465864605e-05
+    1.030212100210257e-05
+   -1.421299844050275e-05
+    1.547184262021354e-05
+   -7.355941479809702e-06
+    1.029924058222109e-05
+   -1.027676755488937e-05
+    8.687362904715759e-06
+ 2.786e+11   
+     8.79690853972037e-06
+   -1.042226637257396e-05
+    1.567131724516732e-05
+    1.040663786120981e-05
+   -1.435801565115117e-05
+     1.56189928038295e-05
+   -7.431139242604066e-06
+    1.040374378477943e-05
+   -1.038251452660355e-05
+    8.765817025709203e-06
+ 2.791e+11   
+    8.876008998549201e-06
+   -1.052887313750698e-05
+    1.581961971409991e-05
+    1.051160724111642e-05
+   -1.450363761000623e-05
+    1.576675004885043e-05
+   -7.506673783406264e-06
+    1.050869965621297e-05
+   -1.048871727742946e-05
+    8.844614146993188e-06
+ 2.796e+11   
+    8.955453039000006e-06
+   -1.063593652015559e-05
+     1.59685304971863e-05
+    1.061702802448743e-05
+   -1.464986274031445e-05
+    1.591511278661191e-05
+   -7.582544313073102e-06
+    1.061410708061203e-05
+   -1.059537470755685e-05
+    8.923753507770736e-06
+ 2.801e+11   
+    9.035239899555415e-06
+    -1.07434554231549e-05
+    1.611804803383784e-05
+    1.072289909719797e-05
+    -1.47966894727283e-05
+    1.606407945612387e-05
+   -7.658750043326313e-06
+    1.071996494526922e-05
+   -1.070248572055459e-05
+     9.00323434815075e-06
+ 2.806e+11   
+    9.115368819301365e-06
+   -1.085142875208693e-05
+    1.626817077046151e-05
+    1.082921934787461e-05
+   -1.494411624458859e-05
+    1.621364850340072e-05
+    -7.73529018649063e-06
+    1.082627214022104e-05
+   -1.081004922294362e-05
+    9.083055908848336e-06
+ 2.811e+11   
+    9.195839037618388e-06
+   -1.095985541504266e-05
+    1.641889715977414e-05
+    1.093598766742662e-05
+   -1.509214149919276e-05
+     1.63638183807787e-05
+   -7.812163955225197e-06
+    1.093302755777937e-05
+   -1.091806412376155e-05
+    9.163217430877929e-06
+ 2.816e+11   
+    9.276649793866154e-06
+   -1.106873432217662e-05
+    1.657022566010495e-05
+    1.104320294856763e-05
+    -1.52407636850502e-05
+    1.651458754622183e-05
+   -7.889370562248636e-06
+    1.104023009205344e-05
+   -1.102652933411938e-05
+    9.243718155239694e-06
+ 2.821e+11   
+    9.357800327061553e-06
+   -1.117806438525385e-05
+    1.672215473468711e-05
+    1.115086408532835e-05
+   -1.538998125512524e-05
+    1.666595446261681e-05
+   -7.966909220058128e-06
+    1.114787863846278e-05
+   -1.113544376675111e-05
+    9.324557322599536e-06
+ 2.826e+11   
+    9.439289875550788e-06
+   -1.128784451719038e-05
+    1.687468285093931e-05
+    1.125896997256083e-05
+   -1.553979266606887e-05
+    1.681791759705788e-05
+    -8.04477914064284e-06
+    1.125597209324181e-05
+    -1.12448063355564e-05
+    9.405734172963088e-06
+ 2.831e+11   
+     9.52111767667583e-06
+   -1.139807363158716e-05
+    1.702780847973788e-05
+    1.136751950543487e-05
+   -1.569019637743967e-05
+     1.69704754201224e-05
+   -8.122979535191938e-06
+    1.136450935293644e-05
+   -1.135461595513705e-05
+    9.487247945344058e-06
+ 2.836e+11   
+     9.60328296643544e-06
+   -1.150875064225823e-05
+    1.718153009468014e-05
+    1.147651157892682e-05
+   -1.584119085091485e-05
+    1.712362640513748e-05
+     -8.2015096137975e-06
+    1.147348931389317e-05
+   -1.146487154032747e-05
+    9.569097877427178e-06
+ 2.841e+11   
+    9.685784979141324e-06
+   -1.161987446275353e-05
+    1.733584617134009e-05
+    1.158594508730173e-05
+   -1.599277454949244e-05
+    1.727736902743912e-05
+   -8.280368585152746e-06
+    1.158291087174149e-05
+   -1.157557200571993e-05
+    9.651283205226353e-06
+ 2.846e+11   
+    9.768622947069651e-06
+   -1.173144400587668e-05
+    1.749075518651656e-05
+     1.16958189235888e-05
+   -1.614494593668479e-05
+    1.743170176362375e-05
+   -8.359555656245626e-06
+     1.16927729208696e-05
+    -1.16867162651847e-05
+    9.733803162737978e-06
+ 2.851e+11   
+     9.85179610010818e-06
+   -1.184345818319827e-05
+      1.7646255617475e-05
+    1.180613197905109e-05
+   -1.629770347570465e-05
+    1.758662309079332e-05
+   -8.439070032048345e-06
+    1.180307435389433e-05
+   -1.179830323138568e-05
+    9.816656981590118e-06
+ 2.856e+11   
+    9.935303665399471e-06
+   -1.195591590456503e-05
+    1.780234594118323e-05
+    1.191688314264966e-05
+    -1.64510456286443e-05
+    1.774213148579463e-05
+   -8.518910915202872e-06
+    1.191381406112555e-05
+   -1.191033181529206e-05
+    9.899843890687606e-06
+ 2.861e+11   
+    1.001914486698048e-05
+   -1.206881607760542e-05
+    1.795902463354224e-05
+    1.202807130050271e-05
+   -1.660497085564842e-05
+    1.789822542445328e-05
+    -8.59907750570287e-06
+    1.202499093002561e-05
+   -1.202280092568613e-05
+    9.983363115853581e-06
+ 2.866e+11   
+    1.010331892541868e-05
+   -1.218215760723175e-05
+    1.811629016861201e-05
+    1.213969533534018e-05
+   -1.675947761408136e-05
+    1.805490338080299e-05
+   -8.679569000572134e-06
+    1.213660384466405e-05
+   -1.213570946866778e-05
+    1.006721387946753e-05
+ 2.871e+11   
+    1.018782505744534e-05
+    -1.22959393951396e-05
+    1.827414101783368e-05
+    1.225175412595423e-05
+   -1.691456435768982e-05
+    1.821216382631117e-05
+   -8.760384593540072e-06
+    1.224865168516845e-05
+   -1.224905634715628e-05
+    1.015139540010045e-05
+ 2.876e+11   
+    1.027266247558579e-05
+   -1.241016033930458e-05
+    1.843257564924821e-05
+      1.2364246546646e-05
+   -1.707022953576087e-05
+    1.837000522910074e-05
+   -8.841523474714155e-06
+    1.236113332717133e-05
+   -1.236284046038929e-05
+    1.023590689214714e-05
+ 2.881e+11   
+    1.035783038778746e-05
+   -1.252481933347697e-05
+    1.859159252671218e-05
+    1.247717146666913e-05
+   -1.722647159227668e-05
+    1.852842605316946e-05
+   -8.922984830249888e-06
+      1.2474047641254e-05
+   -1.247706070341988e-05
+    1.032074756545605e-05
+ 2.886e+11   
+    1.044332799704565e-05
+   -1.263991526667466e-05
+    1.875119010911161e-05
+    1.259052774967044e-05
+   -1.738328896506629e-05
+    1.868742475760692e-05
+   -9.004767842018338e-06
+    1.258739349238729e-05
+   -1.259171596661158e-05
+    1.040591662495696e-05
+ 2.891e+11   
+    1.052915450102737e-05
+   -1.275544702267452e-05
+    1.891136684957387e-05
+    1.270431425312807e-05
+    -1.75406800849547e-05
+    1.884699979580978e-05
+     -9.0868716872716e-06
+    1.270116973937012e-05
+   -1.270680513513218e-05
+    1.049141327028677e-05
+ 2.896e+11   
+    1.061530909169359e-05
+   -1.287141347950279e-05
+    1.907212119467864e-05
+    1.281852982778767e-05
+   -1.769864337491054e-05
+    1.900714961469596e-05
+   -9.169295538306345e-06
+    1.281537523426577e-05
+   -1.282232708844615e-05
+    1.057723669541358e-05
+ 2.901e+11   
+    1.070179095492016e-05
+   -1.298781350892454e-05
+    1.923345158366826e-05
+    1.293317331709682e-05
+   -1.785717724919219e-05
+    1.916787265391823e-05
+   -9.252038562125729e-06
+    1.293000882183654e-05
+   -1.293828069980646e-05
+    1.066338608825948e-05
+ 2.906e+11   
+    1.078859927011752e-05
+    -1.31046459759329e-05
+    1.939535644765793e-05
+    1.304824355663819e-05
+   -1.801628011249345e-05
+    1.932916734507761e-05
+   -9.335099920099914e-06
+    1.304506933897713e-05
+    -1.30546648357459e-05
+    1.074986063032213e-05
+ 2.911e+11   
+    1.087573320984969e-05
+   -1.322190973823793e-05
+    1.955783420884646e-05
+    1.316373937356177e-05
+   -1.817595035908902e-05
+    1.949103211093728e-05
+   -9.418478767625333e-06
+    1.316055561414705e-05
+   -1.317147835556808e-05
+    1.083665949629554e-05
+ 2.916e+11   
+    1.096319193945249e-05
+   -1.333960364575586e-05
+    1.972088327972784e-05
+    1.327965958601644e-05
+   -1.833618637198026e-05
+    1.965346536463723e-05
+   -9.502174253783067e-06
+    1.327646646680242e-05
+   -1.328872011083884e-05
+    1.092378185369021e-05
+ 2.921e+11   
+    1.105097461665154e-05
+   -1.345772654009859e-05
+    1.988450206230416e-05
+    1.339600300258134e-05
+   -1.849698652204198e-05
+    1.981646550891038e-05
+   -9.586185520996393e-06
+    1.339280070682753e-05
+   -1.340638894487778e-05
+     1.10112268624528e-05
+ 2.926e+11   
+    1.113908039118011e-05
+   -1.357627725406419e-05
+    2.004868894730059e-05
+    1.351276842169747e-05
+   -1.865834916717069e-05
+    1.998003093530049e-05
+   -9.670511704687888e-06
+    1.350955713396661e-05
+   -1.352448369225088e-05
+    1.109899367458584e-05
+ 2.931e+11   
+    1.122750840439697e-05
+   -1.369525461112825e-05
+    2.021344231338232e-05
+    1.362995463109955e-05
+   -1.882027265143456e-05
+    2.014416002338222e-05
+   -9.755151932936134e-06
+    1.362673453725585e-05
+   -1.364300317826378e-05
+    1.118708143376734e-05
+ 2.936e+11   
+    1.131625778890466e-05
+   -1.381465742493669e-05
+    2.037876052637457e-05
+    1.374756040724878e-05
+   -1.898275530422595e-05
+    2.030885113998408e-05
+   -9.840105326132374e-06
+    1.374433169445639e-05
+   -1.376194621845672e-05
+    1.127548927497083e-05
+ 2.941e+11   
+    1.140532766816849e-05
+   -1.393448449880015e-05
+    2.054464193848563e-05
+    1.386558451476671e-05
+   -1.914579543941671e-05
+    2.047410263841431e-05
+   -9.925370996637315e-06
+    1.386234737148835e-05
+   -1.388131161810073e-05
+    1.136421632408593e-05
+ 2.946e+11   
+    1.149471715613599e-05
+   -1.405473462519027e-05
+    2.071108488753335e-05
+    1.398402570587054e-05
+   -1.930939135451684e-05
+    2.063991285769049e-05
+   -1.001094804843825e-05
+    1.398078032186627e-05
+   -1.400109817169602e-05
+    1.145326169753978e-05
+ 2.951e+11   
+    1.158442535685779e-05
+   -1.417540658523816e-05
+    2.087808769617599e-05
+    1.410288271981012e-05
+   -1.947354132983681e-05
+    2.080628012177296e-05
+   -1.009683557680674e-05
+    1.409962928613634e-05
+   -1.412130466247219e-05
+     1.15426245019193e-05
+ 2.956e+11   
+    1.167445136410949e-05
+   -1.429649914823537e-05
+     2.10456486711472e-05
+    1.422215428230723e-05
+   -1.963824362765433e-05
+    2.097320273880277e-05
+   -1.018303266795711e-05
+    1.421889299131575e-05
+   -1.424192986189111e-05
+    1.163230383359492e-05
+ 2.961e+11   
+    1.176479426101522e-05
+   -1.441801107113746e-05
+    2.121376610249597e-05
+    1.434183910499704e-05
+   -1.980349649138558e-05
+    2.114067900034434e-05
+   -1.026953839870597e-05
+     1.43385701503344e-05
+   -1.436297252915241e-05
+     1.17222987783457e-05
+ 2.966e+11   
+    1.185545311967284e-05
+   -1.453994109807079e-05
+    2.138243826283181e-05
+    1.446193588487257e-05
+   -1.996929814476168e-05
+    2.130870718063334e-05
+   -1.035635183613305e-05
+    1.445865946147941e-05
+    -1.44844314107019e-05
+    1.181260841098611e-05
+ 2.971e+11   
+    1.194642700078123e-05
+   -1.466228795984238e-05
+    2.155166340657551e-05
+    1.458244330373197e-05
+   -2.013564679101067e-05
+     2.14772855358301e-05
+   -1.044347203724347e-05
+    1.457915960784269e-05
+   -1.460630523974338e-05
+    1.190323179499497e-05
+ 2.976e+11   
+    1.203771495326976e-05
+   -1.478505037345372e-05
+    2.172143976921631e-05
+    1.470336002762953e-05
+   -2.030254061204562e-05
+    2.164641230327932e-05
+   -1.053089804863195e-05
+    1.470006925677193e-05
+   -1.472859273575395e-05
+    1.199416798214642e-05
+ 2.981e+11   
+     1.21293160139303e-05
+   -1.490822704161801e-05
+    2.189176556657484e-05
+    1.482468470633016e-05
+   -2.046997776765898e-05
+    2.181608570077573e-05
+   -1.061862890614885e-05
+    1.482138705932534e-05
+   -1.485129260400313e-05
+    1.208541601214345e-05
+ 2.986e+11   
+    1.222122920705201e-05
+    -1.50318166522821e-05
+    2.206263899407386e-05
+    1.494641597276818e-05
+   -2.063795639472409e-05
+    2.198630392583708e-05
+   -1.070666363456877e-05
+     1.49431116497305e-05
+   -1.497440353507629e-05
+    1.217697491225428e-05
+ 2.991e+11   
+    1.231345354405926e-05
+   -1.515581787815263e-05
+    2.223405822601559e-05
+    1.506855244251059e-05
+    -2.08064746064039e-05
+    2.215706515498415e-05
+   -1.079500124726167e-05
+    1.506524164484784e-05
+   -1.509792420440258e-05
+    1.226884369695162e-05
+ 2.996e+11   
+     1.24059880231526e-05
+   -1.528022937622716e-05
+     2.24060214148671e-05
+      1.5191092713225e-05
+   -2.097553049136751e-05
+    2.232836754302833e-05
+   -1.088364074586691e-05
+    1.518777564363861e-05
+    -1.52218532717874e-05
+    1.236102136755522e-05
* NOTE: Solution at 1e+08 Hz used as DC point.

.model g_m4lines_veryHighFreq_W_1 sp N=4 SPACING=nonuniform VALTYPE=real
+ INTERPOLATION=spline
+ DATA = 600
+ 0           
+    0.0008372886865442828
+   -0.0001520534244311461
+    0.0008425035763071074
+    -1.11451287389565e-06
+    -6.51938693519595e-05
+    0.0008425809538453706
+    1.957382798713116e-07
+   -1.109984968214201e-06
+   -0.0001518854387848884
+    0.0008368313165360179
+ 6e+08       
+     0.005017429006462109
+   -0.0009102275738481465
+     0.005047620513083435
+    -5.96414866986188e-06
+    -0.000389842589887871
+     0.005048094220217097
+    1.720131935089803e-06
+   -5.937072758294419e-06
+   -0.0009092211555692379
+     0.005014657661523924
+ 1.1e+09     
+     0.009231259066633437
+    -0.001672946937706703
+     0.009288783068475271
+   -1.408516479823834e-05
+   -0.0007601735624753161
+     0.009289785739288977
+    1.267267674869101e-05
+   -1.420106735990252e-05
+     -0.00167099743698179
+     0.009225565537327944
+ 1.6e+09     
+      0.01388183092182172
+     -0.00261413343005164
+      0.01398828367929343
+   -4.570866771569296e-05
+    -0.001341321612042763
+      0.01399027612764042
+    7.040530545532857e-05
+   -4.646334567797041e-05
+    -0.002611003570629392
+      0.01387132212559672
+ 2.1e+09     
+      0.01846275620235228
+    -0.003557545617716117
+      0.01862346679971199
+   -6.980629173446245e-05
+     -0.00185663344663722
+      0.01862605352812627
+     0.000126942243648171
+   -7.079154627076474e-05
+    -0.003553592650184061
+      0.01844914712846281
+ 2.6e+09     
+      0.02274415220558276
+    -0.004378653737072533
+      0.02294898890064436
+   -7.572565455140502e-05
+    -0.002263541985113521
+      0.02295189925236723
+    0.0001644531333437698
+   -7.664562510057273e-05
+    -0.004374072130385609
+      0.02272859401886124
+ 3.1e+09     
+      0.02676542251240051
+    -0.005078966974221465
+      0.02699802384499997
+   -6.331666305307608e-05
+    -0.002565091637736418
+       0.0270011488933545
+    0.0001792365465325354
+    -6.40100693668909e-05
+     -0.00507381504920826
+      0.02674846513617401
+ 3.6e+09     
+      0.03063113775183874
+    -0.005696536020416429
+      0.03087420295566512
+   -3.729804765281809e-05
+    -0.002774078226201437
+      0.03087752556851506
+     0.000174493398282612
+   -3.770604687527589e-05
+    -0.005690774599708458
+      0.03061293849699746
+ 4.1e+09     
+      0.03443591231756821
+    -0.006271108552200909
+      0.03467395228178168
+   -4.017375257590585e-06
+    -0.002905749619019002
+      0.03467748797494859
+     0.000156058687344952
+    -4.15942575611645e-06
+    -0.006264629142537411
+      0.03441639887073633
+ 4.6e+09     
+      0.03824708820927396
+    -0.006834653980901202
+      0.03846954685070398
+    3.140230988594127e-05
+    -0.002988136068041495
+      0.03847331555814577
+    0.0001302458064925781
+    3.144937569407678e-05
+    -0.006827309457401775
+      0.03822606307974626
+ 5.1e+09     
+      0.04210608119601462
+    -0.007410821249631128
+      0.04231168904605392
+    6.716246157536436e-05
+     -0.00307403130091158
+      0.04231571079826513
+    0.0001028651041723187
+    6.728894749661023e-05
+    -0.007402469768077833
+      0.04208329549471781
+ 5.6e+09     
+      0.04603392748102114
+     -0.00801689300522768
+      0.04623230626274735
+    0.0001026423886249491
+    -0.003225919234809818
+      0.04623661193798145
+    7.930137619249821e-05
+    0.0001027373582985654
+    -0.008007457149260887
+      0.04600913995142671
+ 6.1e+09     
+      0.05003658596075131
+    -0.008665695360401324
+      0.05024307671288552
+    0.0001324903796813312
+    -0.003474753345168177
+      0.05024772482426081
+    6.520346477844881e-05
+    0.0001324809566780312
+    -0.008655224181567712
+      0.05000961016659303
+ 6.6e+09     
+      0.05410862028112171
+    -0.009365936640167534
+      0.05433655963792931
+    0.0001449296243598803
+    -0.003804247252793194
+      0.05434164588313539
+    6.631225610654289e-05
+    0.0001448251538656005
+    -0.009354635091254613
+      0.05407935236168192
+ 7.1e+09     
+      0.05823498314311745
+     -0.01011996910110526
+      0.05849189319439291
+    0.0001266560004372804
+    -0.004175079355469174
+      0.05849753435426665
+    8.687234681585749e-05
+    0.0001265869247548445
+     -0.01010813885991339
+      0.05820339556851926
+ 7.6e+09     
+      0.06239125685367097
+     -0.01091896617854336
+      0.06267906561333804
+    6.889184255690447e-05
+    -0.004550162862706617
+      0.06268534626031727
+    0.0001273009406432047
+    6.912199579832108e-05
+     -0.01090682446340261
+      0.06235735072293934
+ 8.1e+09     
+      0.06654317572912596
+     -0.01173747904963121
+       0.0668596590341612
+   -2.730773404163532e-05
+    -0.004903016876284065
+      0.06686656387375793
+    0.0001812687371952656
+   -2.642836129310112e-05
+     -0.01172493557784155
+      0.06650691916561259
+ 8.6e+09     
+      0.07064686563006596
+     -0.01253192479927963
+      0.07098687379553814
+   -0.0001439980619740714
+    -0.005217758856897627
+      0.07099427411505103
+    0.0002317086307430996
+   -0.0001421876333677712
+     -0.01251854773848204
+      0.07060819248615738
+ 9.1e+09     
+      0.07465120552198629
+     -0.01324761290521459
+      0.07500759502275109
+   -0.0002350392141447361
+     -0.00548918698455297
+      0.07501534451474913
+    0.0002452178724712535
+   -0.0002324139925888708
+     -0.01323297292429239
+       0.0746101372524085
+ 9.6e+09     
+      0.07850211109772084
+     -0.01383348022223335
+      0.07886667920613133
+   -0.0002099711828582218
+    -0.005725427126900605
+      0.07887476721372332
+    0.0001644125974194315
+    -0.000207614715455543
+     -0.01381770942950047
+      0.07845895723966811
+ 1.01e+10    
+      0.08213055153890718
+     -0.01424381175819639
+      0.08247611796412826
+    -8.53355249128278e-05
+     -0.00590030384862779
+      0.08248369099069057
+   -2.145452667109667e-05
+   -8.615023813690354e-05
+     -0.01422667671249471
+      0.08208223148041646
+ 1.06e+10    
+      0.08562533781652901
+     -0.01452984134426513
+      0.08587113169450593
+   -0.0004995845417002863
+    -0.005862235344548972
+      0.08587392339023879
+     1.27152429057675e-05
+   -0.0005057239312725821
+     -0.01450691157619158
+      0.08555693129048912
+ 1.11e+10    
+      0.08915683819997459
+     -0.01480936723046265
+      0.08930015584617992
+   -0.0009419628603787482
+    -0.005807140524195209
+      0.08929791080677461
+    4.976927765046411e-05
+   -0.0009535087675901222
+     -0.01478063747888523
+      0.08906850177412109
+ 1.16e+10    
+      0.09271864638888699
+     -0.01508264904130751
+      0.09275662038915893
+    -0.001413831474320986
+    -0.005734785784600298
+      0.09274913368566977
+    9.012925422136812e-05
+    -0.001430823813075277
+     -0.01504818574047084
+      0.09261082759499721
+ 1.21e+10    
+      0.09630518562331167
+      -0.0153501654430053
+      0.09623487377568399
+    -0.001916676818664999
+    -0.005645088897282627
+      0.09622199139077357
+    0.0001342820486317617
+    -0.001939105259351426
+      -0.0153100973026296
+      0.09617857364422859
+ 1.26e+10    
+      0.09991164178546752
+     -0.01561257813050679
+      0.09973011826272279
+    -0.002452124630482755
+    -0.005538097362818522
+      0.09971173676676513
+    0.0001827842566167488
+     -0.00247991893229036
+     -0.01556708693914122
+      0.09976711957066871
+ 1.31e+10    
+       0.1035338952812455
+     -0.01587069625736051
+       0.1032383397966483
+    -0.003021955903845223
+    -0.005413965067384677
+       0.1032144054477505
+    0.0002362670768569853
+    -0.003054974660104309
+      -0.0158200082579578
+       0.1033724945830518
+ 1.36e+10    
+       0.1071684534300963
+     -0.01612544201152277
+       0.1067562351512043
+    -0.003628125240802591
+    -0.005272927695473875
+       0.1067267425935404
+    0.0002954416667949025
+    -0.003666142746506406
+     -0.01606982009343472
+       0.1069913137067099
+ 1.41e+10    
+        0.110812384711673
+     -0.01637781785739949
+       0.1102811385409657
+    -0.004272781948621231
+    -0.005115277251717652
+       0.1102461292635837
+    0.0003611050931343134
+    -0.004315472834032531
+     -0.01631755472543422
+       0.1106207164066132
+ 1.46e+10    
+       0.1144632558915581
+     -0.01662887580111912
+       0.1138109494870875
+    -0.004958294289658968
+    -0.004941335945414099
+       0.1137705101944037
+     0.000434147012993051
+    -0.005005215486894555
+     -0.01656428821954166
+       0.1142583082637681
+ 1.51e+10    
+       0.1181190727724138
+     -0.01687968889276868
+       0.1173440633062171
+    -0.005687277354951241
+     -0.00475142959603149
+       0.1172983243408198
+    0.0005155572378322615
+    -0.005737846872006832
+      -0.0168111130575938
+       0.1179021062040726
+ 1.56e+10    
+       0.1217782250867264
+     -0.01713132505749067
+       0.1208793052347187
+    -0.006462625105273474
+    -0.004545860629276638
+       0.1208284391848001
+    0.0006064343506798117
+    -0.006516096971160896
+     -0.01705911312166329
+       0.1215504876218735
+ 1.61e+10    
+       0.1254394358579163
+     -0.01738482324409377
+       0.1244158688901891
+     -0.00728754720634738
+    -0.004324880650226086
+       0.1243600895088623
+    0.0007079955684049539
+    -0.007342981816542161
+     -0.01730934100544912
+       0.1252021436095807
+ 1.66e+10    
+       0.1291017154040937
+     -0.01764117179603163
+        0.127953259513841
+    -0.008165611376382789
+    -0.004088662504121624
+       0.1278928210753963
+    0.0008215880643495026
+    -0.008221840305238828
+     -0.01756279755408124
+       0.1288560363970183
+ 1.71e+10    
+       0.1327643200381002
+     -0.01790128888112909
+       0.1314912422242682
+    -0.009100792065847338
+    -0.003837271665626015
+       0.1314264394447701
+    0.0009487019927797581
+    -0.009156376214825117
+     -0.01782041347502219
+       0.1325113610166072
+ 1.76e+10    
+       0.1364267154250944
+     -0.01816600476353702
+       0.1350297953451214
+     -0.01009752639770017
+     -0.00357063673390305
+       0.1349609640017856
+     0.001090985484119975
+     -0.01015070610830727
+     -0.01808303281813115
+       0.1361675111409898
+ 1.81e+10    
+       0.1400885444903355
+     -0.01843604566049183
+       0.1385690687375469
+      -0.0111607784087283
+    -0.003288518754088671
+        0.138496587133412
+     0.001250261908140548
+     -0.01120941387838523
+     -0.01835139808948111
+        0.139824048985978
+ 1.86e+10    
+       0.1437495997214993
+     -0.01871201889713616
+       0.1421093469706622
+     -0.01229611274170459
+    -0.002990479037550853
+       0.1420336384100762
+     0.001428549728252386
+     -0.01233761272939524
+     -0.01862613674171727
+       0.1434806791314452
+ 1.91e+10    
+       0.1474097996777815
+     -0.01899439905381174
+       0.1456510170924875
+     -0.01350977903075972
+    -0.002675845115603139
+       0.1455725535572006
+     0.001628085290085411
+     -0.01354101541776422
+     -0.01890774877146163
+       0.1471372260839228
+ 1.96e+10    
+       0.1510691694988423
+     -0.01928351479154042
+       0.1491945407150569
+      -0.0148088082792533
+    -0.002343674440857521
+       0.1491138479645698
+     0.001851348895818905
+     -0.01482601354772069
+      -0.0191965951530031
+       0.1507936153842712
+ 2.01e+10    
+       0.1547278251960874
+     -0.01957953604416471
+       0.1527404300959369
+     -0.01620112251528472
+    -0.001992715455193913
+       0.1526580944557032
+     0.002101094501249981
+     -0.01619976661693774
+     -0.01949288684736844
+       0.1544498580496071
+ 2.06e+10    
+       0.1583859615028672
+     -0.01988246128349609
+       0.1562892278802127
+     -0.01769565887290271
+    -0.001621365689545471
+       0.1562059050309643
+      0.00238038332098873
+     -0.01767030127811289
+     -0.01979667415106803
+       0.1581060381267243
+ 2.11e+10    
+       0.1620438430535562
+      -0.0201921046016085
+       0.1598414901554328
+     -0.01930250890281129
+    -0.001227626670322655
+       0.1597579162942822
+     0.002692621513190201
+     -0.01924662085525023
+     -0.02010783619310631
+       0.1617623031209748
+ 2.16e+10    
+       0.1657017986475856
+     -0.02050808242340431
+       0.1633977724672857
+     -0.02103307323513187
+   -0.0008090556193646138
+       0.1633147782742653
+     0.003041601903310025
+     -0.02093882441753079
+     -0.02042607046215355
+       0.1654188570443066
+ 2.21e+10    
+       0.1693602183242244
+     -0.02082979977763931
+       0.1669586184368503
+     -0.02290023050119607
+   -0.0003627143011976251
+         0.16687714634641
+     0.003431549339563978
+     -0.02275823350810225
+     -0.02075088236099246
+       0.1690759557920561
+ 2.26e+10    
+       0.1730195529142443
+     -0.02115643624160289
+       0.1705245506111055
+     -0.02491851736690127
+    0.0001148840187538093
+       0.1704456759463598
+     0.003867168668212783
+     -0.02471752270905905
+     -0.02108157496259216
+        0.172733904499949
+ 2.31e+10    
+       0.1766803156263045
+     -0.02148693197144081
+       0.1740960631604251
+     -0.02710431318197423
+    0.0006278275663671919
+       0.1740210197232924
+     0.004353693348409861
+     -0.02683084724768368
+     -0.02141723941298912
+       0.1763930564370498
+ 2.36e+10    
+       0.1803430850416164
+     -0.02181997469458298
+       0.1776736160056818
+     -0.02947601742349733
+     0.001180855532996376
+       0.1776038266998935
+     0.004896931209160114
+     -0.02911395630289207
+     -0.02175674683446316
+       0.1800538128372458
+ 2.41e+10    
+       0.1840085085880571
+     -0.02215398925815116
+       0.1812576299087411
+     -0.03205419980120894
+     0.001779398208374547
+       0.1811947428547947
+     0.005503301515388926
+     -0.03158427382976081
+     -0.02209874319376487
+       0.1837166228337725
+ 2.46e+10    
+       0.1876773050855291
+     -0.02248713242247127
+       0.1848484819876044
+     -0.03486169013348955
+     0.002429598377299806
+       0.1847944122886788
+     0.006179853967314186
+     -0.03426091856312845
+     -0.02244164950506232
+       0.1873819822994197
+ 2.51e+10    
+       0.1913502642114863
+     -0.02281729723720665
+        0.188446501016519
+     -0.03792355582667793
+     0.003138299251151343
+       0.1884034777193521
+     0.006934254967342493
+     -0.03716462000277237
+       -0.022783671062436
+       0.1910504298578177
+ 2.56e+10    
+       0.1950282396121095
+     -0.02314213378172071
+       0.1920519617405184
+     -0.04126688617235192
+     0.003912976373283476
+       0.1920225783983711
+     0.007774718721829077
+     -0.04031746581076359
+     -0.02312282130605218
+       0.1947225375493245
+ 2.61e+10    
+       0.1987121307259288
+      -0.0234590965999203
+       0.1956650772747786
+     -0.04492026109600188
+     0.004761579681050178
+       0.1956523425446594
+     0.008709849583858315
+     -0.04374238597554962
+     -0.02345696862343666
+       0.1983988925267895
+ 2.66e+10    
+       0.2024028460116695
+     -0.02376553417107867
+       0.1992859884845849
+     -0.04891272330004078
+     0.005692236188092729
+       0.1992933699224912
+     0.009748346460000659
+     -0.04746223802165628
+     -0.02378391808831883
+       0.2020800646326357
+ 2.71e+10    
+       0.2061012370103423
+     -0.02405884254833249
+       0.2029147490798225
+     -0.05327199332383716
+     0.006712742703927398
+       0.2029461981180609
+      0.01089849924404961
+     -0.05149830387194913
+     -0.02410154500490192
+       0.2057665527052765
+ 2.76e+10    
+       0.2098079884697189
+     -0.02433671391625282
+       0.2065513050591755
+     -0.05802156652380396
+     0.007829751647976597
+       0.2066112433249473
+      0.01216738112500923
+      -0.0558679436421191
+     -0.02440800309803165
+       0.2094587000029655
+ 2.81e+10    
+       0.2135234449190515
+     -0.02459752054849641
+        0.210195467168916
+     -0.06317621818922269
+     0.009047523741892976
+       0.2102887031907262
+      0.01355961163313325
+      -0.0605810818557446
+     -0.02470203665489776
+       0.2131565664603543
+ 2.86e+10    
+       0.2172473497280034
+     -0.02484088303857753
+       0.2138468752679046
+      -0.0687353474681591
+      0.01036609682155011
+       0.2139784062071172
+      0.01507554102988518
+     -0.06563514748303691
+     -0.02498343110321345
+       0.2168597433108581
+ 2.91e+10    
+       0.2209784715701751
+     -0.02506847290667004
+       0.2175049539042075
+     -0.07467358205856944
+      0.01177871782978454
+       0.2176795910764822
+      0.01670870461673648
+     -0.07100809470771358
+     -0.02525363646391256
+       0.2205670954608593
+ 2.96e+10    
+       0.2247141008639479
+     -0.02528508229613625
+       0.2211688588038983
+     -0.08092828002009288
+      0.01326843933607623
+         0.22139060424081
+      0.01844244956264695
+      -0.0766492780113374
+     -0.02551658543623674
+       0.2242764217826133
+ 3.01e+10    
+       0.2284494244967821
+     -0.02549993842398829
+       0.2248374138035858
+     -0.08738422779546838
+      0.01480394865045147
+       0.2251085208405151
+      0.02024580242799172
+     -0.08246837320636098
+     -0.02577969063178886
+       0.2279840378594967
+ 3.06e+10    
+       0.2321768433866954
+     -0.02572812274963061
+       0.2285090362100276
+      -0.0938572375782226
+      0.01633504989526522
+       0.2288287325514494
+        0.022068995163031
+     -0.08832339270334497
+     -0.02605492821270628
+       0.2316843157830876
+ 3.11e+10    
+       0.2358853938931378
+     -0.02599175569027744
+       0.2321816454783635
+      -0.1000807055720412
+      0.01778881341731356
+       0.2325446117035788
+      0.02383965649906008
+     -0.09401026940598024
+     -0.02635978566533016
+       0.2353692665603577
+ 3.16e+10    
+       0.2395605619454785
+     -0.02632034659847146
+       0.2358525484045465
+      -0.1057022546722165
+      0.01906819225282009
+       0.2362474474878911
+       0.0254614540416328
+     -0.09925838496362849
+     -0.02671767814841473
+       0.2390283204973075
+ 3.21e+10    
+       0.2431848847341198
+     -0.02674949530027799
+       0.2395183032776716
+      -0.1103000214104468
+      0.02005557818389721
+       0.2399269163298429
+      0.02681763836438807
+      -0.1037381611175362
+     -0.02715727929404249
+       0.2426485293574316
+ 3.26e+10    
+       0.2467397033849037
+     -0.02731720043098457
+       0.2431746010632674
+      -0.1134271584509173
+      0.02062366565163529
+       0.2435723091319281
+      0.02778183477331177
+      -0.1070869768219063
+     -0.02771020157872035
+       0.2462154321560039
+ 3.31e+10    
+       0.2502081221423767
+     -0.02805766208843519
+       0.2468162694415366
+      -0.1146854253734651
+      0.02065427647611716
+       0.2471744967752594
+      0.02823672477284974
+      -0.1089562482355635
+     -0.02840677869693344
+       0.2497147222917451
+ 3.36e+10    
+       0.2535786227450152
+     -0.02899370822463256
+       0.2504375688546071
+      -0.1138139454411482
+      0.02006222207370861
+       0.2507281763240897
+       0.0280977115302817
+      -0.1090744512764521
+     -0.02927043938515314
+       0.2531345778419364
+ 3.41e+10    
+       0.2568481441353834
+     -0.03013028949586268
+       0.2540329165487353
+      -0.1107638991463419
+      0.01881719141853519
+       0.2542335319604077
+      0.02733461152148185
+      -0.1073103486789653
+     -0.03031210839148768
+       0.2564681253543373
+ 3.46e+10    
+         0.26002328359911
+     -0.03145183231132306
+       0.2575979697645538
+      -0.1057265326902492
+      0.01695499186515233
+       0.2576964525069604
+      0.02598277356665267
+      -0.1037140173146884
+     -0.03152664298565251
+       0.2597152128643739
+ 3.51e+10    
+       0.2631189436306619
+     -0.03292491109418075
+       0.2611307030447462
+     -0.09909834776327431
+      0.01457261389331827
+       0.2611270536458995
+      0.02413815153312785
+     -0.09851737064916521
+     -0.03289290109770332
+       0.2628827410965834
+ 3.56e+10    
+       0.2661549291267948
+      -0.0345052882451242
+       0.2646319768882439
+     -0.09139608203235104
+       0.0118085037723137
+       0.2645371144717578
+      0.02193771550096314
+      -0.0920913600671526
+     -0.03437762420915593
+       0.2659833238305196
+ 3.61e+10    
+       0.2691518804763535
+     -0.03614650428822125
+       0.2681052970023773
+      -0.0831555024153144
+     0.008815705853154669
+       0.2679375143071503
+      0.01953280798568141
+      -0.0848752767028572
+     -0.03594171152305357
+       0.2690327493401918
+ 3.66e+10    
+       0.2721279480296348
+     -0.03780706593169406
+       0.2715558798594454
+     -0.07484855783746247
+     0.005737198854540947
+       0.2713365408323268
+      0.01706469287448953
+     -0.07730301305864562
+     -0.03754667840037904
+       0.2720471514305643
+ 3.71e+10    
+       0.2750969412119056
+     -0.03945460379561523
+       0.2749894490770637
+     -0.06683707851336643
+     0.002689652494194963
+       0.2747393239694356
+      0.01464846597911449
+     -0.06974727252361003
+     -0.03915948354297408
+       0.2750407363400137
+ 3.76e+10    
+       0.2780679148813737
+     -0.04106697288145083
+       0.2784112008907582
+     -0.05936229169357705
+   -0.0002430005896755169
+       0.2781481301026331
+      0.01236670283930539
+     -0.06249072266449397
+     -0.04075498173135823
+       0.2780244923540036
+ 3.81e+10    
+       0.2810457169731491
+     -0.04263123474897733
+       0.2818251751577808
+      -0.0525584922704753
+     -0.00300832962074799
+       0.2815630709020089
+      0.01027070376696809
+     -0.05572158788582302
+     -0.04231625517091933
+       0.2810058557096156
+ 3.86e+10    
+        0.284031962482485
+     -0.04414164169923761
+       0.2852340425051065
+     -0.04647757895650906
+    -0.005579889217814316
+       0.2849828661751714
+     0.008385979460718177
+     -0.04954522591264957
+     -0.04383357506426684
+       0.2839890421224324
+ 3.91e+10    
+        0.287026048524593
+     -0.04559746337078065
+       0.2886391884493796
+     -0.04111476762603319
+    -0.007950339744482069
+       0.2884054709551634
+     0.006719083202609402
+     -0.04400278749364604
+     -0.04530276762838783
+       0.2869757048262966
+ 3.96e+10    
+       0.2900260116834824
+     -0.04700111120584847
+        0.292040950009658
+     -0.03643040576757412
+     -0.01012502452317678
+       0.2918285146079694
+     0.005263985848781298
+     -0.03909053955181278
+     -0.04672353589077991
+       0.2899656592595617
+ 4.01e+10    
+       0.2930291666784549
+     -0.04835671754637558
+       0.2954388933965267
+     -0.03236627783351767
+     -0.01211681390146355
+       0.2952495728397481
+     0.004007191790935825
+     -0.03477642000957588
+         -0.0480980283546
+        0.292957526102704
+ 4.06e+10    
+       0.2960325403354489
+      -0.0496691557537954
+       0.2988320682837407
+     -0.02885670854459658
+     -0.01394236615621751
+       0.2986663172784025
+      0.00293144836011504
+     -0.03101265922698093
+     -0.04942975085342886
+       0.2959492346790712
+ 4.11e+10    
+       0.2990331436329244
+     -0.05094341711943923
+       0.3022192118745911
+      -0.0258355268868378
+     -0.01561962723454052
+        0.302076585591439
+     0.002018226027319903
+     -0.02774460545026862
+     -0.05072280715403198
+       0.2989383835419978
+ 4.16e+10    
+       0.3020281279033968
+     -0.05218424741845777
+       0.3055988989221418
+     -0.02324005654492054
+     -0.01716628366483561
+       0.3054784046715638
+     0.001249253188155366
+     -0.02491644701000781
+     -0.05198140728266446
+       0.3019224804025138
+ 4.21e+10    
+       0.3050148639080382
+     -0.05339595883653832
+       0.3089696447678428
+     -0.02101312134304028
+     -0.01859888997845778
+       0.3088699885598251
+    0.0006073821224541029
+     -0.02247463704074813
+      -0.0532095736110958
+       0.3048990905300419
+ 4.26e+10    
+       0.3079909725788028
+     -0.05458235326355373
+       0.3123299718872056
+     -0.01910380540067163
+     -0.01993244383881328
+        0.312249724347139
+    7.701114582853315e-05
+     -0.02036973307225927
+     -0.05441098319744907
+       0.3078659206402233
+ 4.31e+10    
+        0.310954327282318
+     -0.05574671210789286
+       0.3156784500810266
+     -0.01746748018375916
+     -0.02118024173852102
+       0.3156161535885008
+   -0.0003557712836727604
+     -0.01855720477311933
+     -0.05558889875196357
+       0.3108208598642052
+ 4.36e+10    
+       0.3139030405667907
+     -0.05689182295753126
+        0.319013718638776
+     -0.01606543373267219
+     -0.02235389992784991
+       0.3189679532137552
+   -0.0007032061514962318
+     -0.01699760699845018
+     -0.05674615409497145
+       0.3137619936378247
+ 4.41e+10    
+       0.3168354434752733
+     -0.05802002435364195
+        0.322334496727224
+     -0.01486431145354536
+     -0.02346346485124006
+       0.3223039178416237
+   -0.0009759721121346803
+      -0.0156563877582716
+     -0.05788517095675687
+       0.3166876014679002
+ 4.46e+10    
+       0.3197500622426898
+     -0.05913325737263447
+       0.3256395864342855
+     -0.01383549325603075
+     -0.02451756549559678
+       0.3256229442514943
+    -0.001183335195886073
+     -0.01450350608502748
+     -0.05900799210148878
+       0.3195961458208182
+ 4.51e+10    
+       0.3226455950958981
+     -0.06023311754499626
+       0.3289278714736712
+     -0.01295447732550968
+     -0.02552357904339562
+       0.3289240181646977
+    -0.001333311666493801
+     -0.01351296867961075
+     -0.06011632143002193
+       0.3224862567362264
+ 4.56e+10    
+       0.3255208905737688
+     -0.06132090367262816
+        0.332198313519356
+     -0.01220030695002319
+     -0.02648779356275009
+       0.3322062031978776
+    -0.001432827928988365
+     -0.01266235000769028
+      -0.0612115655093322
+       0.3253567149718063
+ 4.61e+10    
+       0.3283749280031382
+     -0.06239766194488031
+       0.3354499474148268
+     -0.01155505650623885
+      -0.0274155592193717
+       0.3354686317323934
+     -0.00148786906907486
+     -0.01193233196468237
+     -0.06229487342406954
+        0.328206435305011
+ 4.66e+10    
+       0.3312068003159185
+     -0.06346422482699415
+       0.3386818760163149
+     -0.01100338101111059
+      -0.0283114242074092
+       0.3387104974110997
+    -0.001503612273428308
+     -0.01130628136359487
+     -0.06336717337913045
+       0.3310344508665626
+ 4.71e+10    
+       0.3340156991474428
+       -0.064521244789898
+       0.3418932651099526
+     -0.01053212728622724
+      -0.0291792543501786
+       0.3419310489894645
+    -0.001484544105501591
+     -0.01076987269894114
+     -0.06442920540857153
+       0.3338398989162621
+ 4.76e+10    
+       0.3368009020332083
+     -0.06556922325335258
+       0.3450833386395378
+     -0.01013000163725482
+     -0.03002233684383945
+       0.3451295852940803
+    -0.001434562117988331
+     -0.01031075737819775
+     -0.06548155008415692
+       0.3366220081953006
+ 4.81e+10    
+       0.3395617614711355
+       -0.066608535246807
+       0.3482513743552779
+    -0.009787287684577244
+     -0.03084346938909297
+       0.3483054510810256
+    -0.001357062045023034
+    -0.009918277198788321
+     -0.06652465341067185
+       0.3393800878321342
+ 4.86e+10    
+       0.3422976956065351
+     -0.06763945032603733
+       0.3513966999174846
+    -0.009495607766411285
+     -0.03164503627769441
+       0.3514580336183147
+    -0.001255012135249327
+    -0.009583218177313666
+     -0.06755884823921915
+       0.3421135176960839
+ 4.91e+10    
+       0.3450081803083367
+     -0.06866215026483766
+       0.3545186894464215
+     -0.00924772167522997
+     -0.03242907307102567
+       0.3545867598496757
+    -0.001131016252336619
+     -0.00929760019798891
+     -0.06858437258548408
+       0.3448217400555698
+ 4.96e+10    
+       0.3476927424272216
+     -0.06967674399694969
+       0.3576167604854882
+    -0.009037357086229113
+     -0.03319732143357914
+       0.3576910940224071
+   -0.0009873672981630895
+    -0.009054497897519623
+     -0.06960138524482426
+       0.3475042523863463
+ 5.01e+10    
+       0.3503509540508147
+     -0.07068328022778819
+        0.360690371334764
+    -0.008859066723150476
+     -0.03395127555099803
+       0.3607705356855482
+   -0.0008260923769167377
+    -0.008847888463335294
+     -0.07060997907420841
+       0.3501606011789191
+ 5.06e+10    
+       0.3529824275975349
+     -0.07168175808090649
+       0.3637390187086675
+    -0.008708107993932878
+     -0.03469222139471526
+       0.3638246179810551
+   -0.0006489909542671071
+    -0.008672522433958944
+     -0.07161019227620954
+       0.3527903766055909
+ 5.11e+10    
+       0.3555868116134458
+     -0.07267213609000361
+       0.3667622356721815
+    -0.008580341464138891
+     -0.03542126993232319
+       0.3668529061682687
+   -0.0004576671018594672
+    -0.008523814049328046
+     -0.07260201798134108
+       0.3553932079221468
+ 5.16e+10    
+       0.3581637871581904
+     -0.07365433980016753
+       0.3697595898141315
+    -0.008472145105255825
+     -0.03613938522390712
+       0.3698549963311211
+   -0.0002535567599142973
+     -0.00839774815864648
+     -0.07358541238514507
+       0.3579687594943871
+ 5.21e+10    
+       0.3607130646843654
+     -0.07462826820012937
+       0.3727306816189948
+    -0.008380341748483016
+     -0.03684740820487188
+       0.3728305142298819
+   -3.795081194550706e-05
+    -0.008290801119128343
+     -0.07456030166115035
+       0.3605167273550943
+ 5.26e+10    
+       0.3632343813302755
+     -0.07559379917112322
+       0.3756751430049033
+    -0.008302137596267673
+     -0.03754607683095718
+       0.3757791142647394
+    0.0001879853593255414
+    -0.008199873504209275
+     -0.07552658783673125
+       0.3630368362101929
+ 5.31e+10    
+       0.3657274985599023
+     -0.07655079410813528
+       0.3785926359987261
+    -0.008235070001658084
+     -0.03823604315427138
+       0.3787004785269084
+    0.0004231952708892298
+    -0.008122232775002031
+     -0.07648415379103997
+       0.3655288368254297
+ 5.36e+10    
+       0.3681922000944063
+     -0.07749910184257319
+       0.3814828515242356
+    -0.008176963023980476
+     -0.03891788780833052
+        0.381594315916422
+    0.0006667172211996617
+    -0.008055464359738402
+     -0.07743286750887041
+       0.3679925037353065
+ 5.41e+10    
+       0.3706282900893632
+     -0.07843856197510808
+        0.384345508282227
+    -0.008125889519300437
+     -0.03959213230207171
+       0.3844603613103533
+    0.0009176722583567154
+    -0.007997429833035958
+     -0.07837258570311441
+       0.3704276332252617
+ 5.46e+10    
+       0.3730355915194691
+     -0.07936900770819484
+       0.3871803517050482
+    -0.008080138732087043
+     -0.04025924945886573
+       0.3872983747693938
+     0.001175253903790619
+     -0.00794623109665334
+      -0.0793031569008729
+       0.3728340415458606
+ 5.51e+10    
+       0.3754139447389058
+     -0.08029026825443618
+       0.3899871529722965
+    -0.008038188525754044
+     -0.04091967228251159
+       0.3901081407712065
+     0.001438719353638812
+    -0.007900179639576874
+     -0.08022442407246147
+       0.3752115633243731
+ 5.56e+10    
+       0.3777632061909595
+     -0.08120217088304593
+       0.3927657080738405
+    -0.007998681534094653
+     -0.04157380148528674
+       0.3928894674638989
+     0.001707381926190518
+    -0.007857770103858373
+     -0.08113622687056141
+        0.377560050144561
+ 5.61e+10    
+       0.3800832472446772
+     -0.08210454265741285
+       0.3955158369116866
+    -0.007960404632448289
+     -0.04222201187725217
+       0.3956421859320268
+     0.001980604560480149
+    -0.007817657506056497
+     -0.08203840353559416
+       0.3798793692703661
+ 5.66e+10    
+        0.382373953140492
+     -0.08299721190813131
+       0.3982373824318092
+    -0.007922271226452478
+     -0.04286465778331174
+       0.3983661494711475
+     0.002257794203163197
+    -0.007778637568100136
+      -0.0829307925148363
+       0.3821694024928721
+ 5.71e+10    
+       0.3846352220289894
+     -0.08388000947802604
+       0.4009302097793531
+    -0.007883305937533515
+     -0.04350207762804606
+       0.4010612328659972
+     0.002538396947245045
+     -0.00773962969834353
+     -0.08381323383489016
+       0.3844300450832749
+ 5.76e+10    
+       0.3868669640904147
+     -0.08475276977137007
+       0.4035942054727177
+    -0.007842631330988205
+      -0.0441345978082715
+       0.4037273316709218
+      0.00282189380702492
+    -0.007699662234886769
+     -0.08468557026179928
+       0.3866612048375807
+ 5.81e+10    
+       0.3890691007235455
+      -0.0856153316321871
+       0.4062292765900921
+    -0.007799456389876736
+     -0.04476253595169481
+       0.4063643614885249
+     0.003107797033845826
+    -0.007657859625272613
+     -0.08554764827638162
+       0.3888628012002018
+ 5.86e+10    
+       0.3912415637955146
+     -0.08646753907571426
+       0.4088353499678791
+    -0.007753066483732383
+     -0.04538620364836018
+       0.4089722572467448
+     0.003395646890419334
+    -0.007613431265794663
+     -0.08639931889011322
+         0.39103476445696
+ 5.91e+10    
+       0.3933842949442977
+     -0.08730924189029728
+       0.4114123714058369
+    -0.007702814620337574
+     -0.04600590872611912
+       0.4115509724721722
+     0.003685008816118709
+    -0.007565661767310463
+     -0.08724043832082554
+       0.3931770349878063
+ 5.96e+10    
+       0.3954972449278606
+     -0.08814029612675334
+       0.4139603048783508
+    -0.007648113801903878
+     -0.04662195713170736
+       0.4141004785596715
+     0.003975470925497206
+    -0.007513902448958013
+      -0.0880708685467112
+       0.3952895625727169
+ 6.01e+10    
+        0.397580373014072
+      -0.0889605644884022
+       0.4164791317497682
+    -0.007588430332849982
+     -0.04723465447026289
+       0.4166207640371792
+     0.004266641791143741
+    -0.007457563891579989
+     -0.08889047775269282
+       0.3973723057437071
+ 6.06e+10    
+       0.3996336464072376
+     -0.08976991663370193
+       0.4189688499923558
+    -0.007523277951236472
+     -0.04784430724739621
+       0.4191118338269427
+     0.004558148470894056
+    -0.007396109407800909
+     -0.08969914068269895
+       0.3994252311782589
+ 6.11e+10    
+       0.4016570397067643
+     -0.09056822940144889
+       0.4214294734072804
+    -0.007452212672788249
+     -0.04845122385331431
+       0.4215737085018081
+     0.004849634744201844
+    -0.007329049306409097
+     -0.09049673890794309
+       0.4014483131291314
+ 6.16e+10    
+       0.4036505343949824
+     -0.09135538696682756
+       0.4238610308467571
+    -0.007374828254907552
+     -0.04905571532109108
+        0.424006423538307
+     0.005140759529002538
+    -0.007255935846854194
+     -0.09128316102120893
+       0.4034415328868157
+ 6.21e+10    
+       0.4056141183510034
+     -0.09213128093631445
+       0.4262635654376602
+    -0.007290752199767308
+     -0.04965809588749884
+       0.4264100285658896
+     0.005431195454881564
+    -0.007176358794644368
+     -0.09205830276500175
+       0.4054048782713592
+ 6.26e+10    
+       0.4075477853883147
+     -0.09289581038740576
+        0.428637133807414
+    -0.007199642227987735
+     -0.05025868338261147
+       0.4287845866140043
+     0.005720627571861952
+    -0.007089941501044283
+     -0.09282206710057418
+       0.4073383431505145
+ 6.31e+10    
+       0.4094515348137235
+     -0.09364888185888418
+       0.4309818053107519
+    -0.007101183164345546
+     -0.05085779946744021
+        0.431130173356459
+      0.00600875217749427
+    -0.006996337441518289
+     -0.09357436422395177
+       0.4092419269819011
+ 6.36e+10    
+       0.4113253710061872
+     -0.09439040929657432
+       0.4332976612589057
+    -0.006995084184702981
+     -0.05145576973895373
+       0.4334468763547685
+     0.006295275748268686
+    -0.006895227156273661
+     -0.09431511153423372
+       0.4111156343769172
+ 6.41e+10    
+       0.4131693030134643
+     -0.09512031395847766
+       0.4355847941505302
+     -0.00688107638052312
+     -0.05205292371927452
+       0.4357347943009812
+     0.006579913963111078
+    -0.006786315544353364
+     -0.09504423355891717
+       0.4129594746845808
+ 6.46e+10    
+        0.414983344165712
+     -0.09583852428392256
+        0.437843306906472
+    -0.006758910603112392
+     -0.05264959474240377
+       0.4379940362604837
+     0.006862390808639286
+    -0.006669329468801748
+     -0.09576166184017271
+       0.4147734615938213
+ 6.51e+10    
+       0.4167675117043868
+     -0.09654497572855021
+       0.4400733121060253
+     -0.00662835555591528
+     -0.05324611975014275
+       0.4402247209160315
+     0.007142437758722664
+    -0.006544015637415308
+     -0.09646733478559757
+       0.4165576127525008
+ 6.56e+10    
+       0.4185218264257656
+     -0.09723961056974709
+       0.4422749312290991
+     -0.00648919610534969
+     -0.05384283901013855
+       0.4424269758135596
+     0.007419793020290952
+    -0.006410138726250835
+      -0.0971611974869839
+       0.4183119494024106
+ 6.61e+10    
+       0.4202463123378828
+     -0.09792237768373668
+       0.4444482939006667
+    -0.006341231787203924
+      -0.0544400957625086
+       0.4446009366106424
+     0.007694200840857373
+    -0.006267479719805229
+     -0.09784320150961751
+       0.4200364960288279
+ 6.66e+10    
+       0.4219409963302795
+     -0.09859323229752014
+       0.4465935371420967
+    -0.006184275486087889
+     -0.05503823580692634
+       0.4467467463286408
+     0.007965410872308277
+    -0.006115834443205214
+     -0.09851330465440458
+       0.4217312800236482
+ 6.71e+10    
+       0.4236059078558196
+     -0.09925213571732622
+        0.448710804626538
+    -0.006018152270143564
+     -0.05563760703417765
+       0.4488645546089898
+     0.008233177587283006
+    -0.005955012266010253
+     -0.09917147069581791
+       0.4233963313617595
+ 6.76e+10    
+       0.4252410786237824
+     -0.09989905503547342
+       0.4508002459414869
+    -0.005842698364520701
+     -0.05623855891152674
+        0.450954516974669
+     0.008497259745445244
+    -0.005784834959417676
+     -0.09981766909687384
+       0.4250316822892747
+ 6.81e+10    
+       0.4268465423041443
+      -0.1005339628179471
+       0.4528620158583442
+    -0.005657760249651679
+     -0.05684144192617661
+       0.4530167940979137
+     0.008757419906513242
+    -0.005605135690942256
+      -0.1004518747037016
+        0.426637367023637
+ 6.86e+10    
+       0.4284223342419371
+      -0.1011568367730693
+       0.4548962736080212
+    -0.005463193871954721
+     -0.05744660699173471
+       0.4550515510735672
+     0.009013423988459193
+     -0.00541575814320501
+      -0.1010740674206943
+       0.4282134214644288
+ 6.91e+10    
+        0.429968491181793
+      -0.1017676594041245
+       0.4569031821670286
+    -0.005258863955483754
+     -0.05805440482479592
+       0.4570589567013215
+     0.009265040868736602
+    -0.005216555743433918
+      -0.1016842318684981
+       0.4297598829150382
+ 6.96e+10    
+       0.4314850510021366
+      -0.1023664176461111
+       0.4588829075498088
+    -0.005044643406015356
+     -0.05866518529204001
+       0.4590391827746946
+     0.009512042027559162
+    -0.005007390994421938
+      -0.1022823570257058
+       0.4312767898141448
+ 7.01e+10    
+       0.4329720524584927
+        -0.10295310248852
+       0.4608356181121808
+    -0.004820412797858114
+     -0.05927929673542462
+       0.4609924033794282
+     0.009754201231926992
+    -0.004788134896107913
+      -0.1028684358556599
+       0.4327641814769936
+ 7.06e+10    
+       0.4344295349359587
+       -0.103527708584978
+       0.4627614838634544
+    -0.004586059936894642
+     -0.05989708527606837
+       0.4629187942012566
+       0.0099912942591863
+    -0.004558666450353169
+      -0.1034424649200552
+       0.4342220978461199
+ 7.11e+10    
+        0.435857538210316
+      -0.1040902338509156
+       0.4646606757892552
+    -0.004341479492503303
+     -0.06051889410113122
+       0.4648185318431621
+      0.01022309865957337
+    -0.004318872240809844
+        -0.10400444397957
+       0.4356505792509886
+ 7.16e+10    
+       0.4372561022177479
+      -0.1046406790505258
+       0.4665333651857371
+    -0.004086572692801077
+      -0.0611450627367188
+       0.4666917931541016
+      0.01044939355701125
+    -0.004068646081583232
+      -0.1045543755837855
+       0.4370496661765522
+ 7.21e+10    
+       0.4386252668327105
+      -0.1051790473733424
+        0.468379723004041
+    -0.003821247077541916
+     -0.06177592630841332
+       0.4685387545677359
+      0.01066995948678833
+    -0.003807888728539264
+      -0.1050922646501487
+       0.4384193990402993
+ 7.26e+10    
+       0.4399650716540712
+      -0.1057053440021673
+       0.4701999192072872
+    -0.003545416304435717
+     -0.06241181479255622
+       0.4703595914539327
+      0.01088457827047823
+    -0.003536507648073498
+      -0.1056181180339875
+       0.4397598179776601
+ 7.31e+10    
+       0.4412755557992322
+      -0.1062195756726731
+       0.4719941221401422
+    -0.003259000003994518
+     -0.06305305226016852
+       0.4721544774813501
+      0.01109303292657173
+     -0.00325441683871454
+       -0.106131944089883
+       0.4410709626356314
+ 7.36e+10    
+       0.4425567577058768
+      -0.1067217502256116
+        0.473762497910112
+    -0.002961923679254923
+     -0.06369995611533194
+       0.4739235839933892
+      0.01129510761599233
+    -0.002961536700622664
+      -0.1066337522255723
+       0.4423528719742865
+ 7.41e+10    
+       0.4438087149416722
+      -0.1072118761526578
+       0.4755052097821343
+    -0.002654118647191426
+      -0.0643528363300937
+       0.4756670793967089
+      0.01149058762276699
+    -0.002657793949817476
+      -0.1071235524489743
+       0.4436055840761413
+ 7.46e+10    
+       0.4450314640213039
+       -0.107689962136459
+       0.4772224175871383
+     -0.00233552201810988
+     -0.06501199467692335
+       0.4773851285629389
+      0.01167925936785925
+    -0.002343121573293953
+      -0.1076013549095815
+       0.4448291359634047
+ 7.51e+10    
+       0.4462250402312076
+      -0.1081560165859404
+        0.478914277143853
+    -0.002006076709990997
+     -0.06567772396197699
+       0.4790778922449861
+      0.01186091045554815
+    -0.002017458821398632
+      -0.1080671694345003
+        0.446023563422534
+ 7.56e+10    
+       0.4473894774615549
+      -0.1086100471672645
+       0.4805809396941755
+     -0.00166573149601935
+     -0.06635030725788653
+       0.4807455265063347
+      0.01203532975246406
+    -0.001680751235172539
+      -0.1085210050604755
+       0.4471889008365019
+ 7.61e+10    
+       0.4485248080456077
+      -0.1090520603316175
+       0.4822225513543625
+    -0.001314441081437339
+     -0.06703001714052491
+       0.4823881821658141
+      0.01220230749646344
+    -0.001332950705136665
+      -0.1089628695623147
+        0.448325181024409
+ 7.66e+10    
+       0.4496310626062429
+      -0.1094820608400813
+       0.4838392525785596
+   -0.0009521662085790836
+     -0.06771711492835161
+       0.4840060042560937
+      0.01236163543618037
+    -0.000974015559984226
+      -0.1093927689781855
+       0.4494324350881407
+ 7.71e+10    
+       0.4507082699097627
+      -0.1099000512869986
+       0.4854311776396577
+   -0.0005788737871461045
+     -0.06841184992782187
+       0.4855991314978135
+      0.01251310699837989
+   -0.0006039106813963686
+      -0.1098107071337426
+       0.4505106922667141
+ 7.76e+10    
+        0.451756456726652
+      -0.1103060316217472
+       0.4869984541232155
+   -0.0001945370482095701
+     -0.06911445868357065
+       0.4871676957888785
+      0.01265651748358883
+   -0.0002226076445430492
+      -0.1102166851642599
+       0.4515599797974041
+ 7.81e+10    
+       0.4527756476996256
+      -0.1106999986704304
+       0.4885412024374542
+    0.0002008642805925533
+     -0.06982516423760836
+       0.4887118217088355
+      0.01279166428700335
+    0.0001699151198678514
+      -0.1106107010366151
+        0.452580322784065
+ 7.86e+10    
+       0.4537658652184268
+      -0.1110819456577466
+       0.4900595353392815
+    0.0006073437794957323
+     -0.07054417539526557
+       0.4902316260392892
+      0.01291834714526504
+    0.0005736721416855928
+      -0.1109927490714764
+       0.4535717440725357
+ 7.91e+10    
+       0.4547271293018745
+      -0.1114518617298103
+       0.4915535574746043
+     0.001024908123352512
+       -0.071271686001217
+       0.4917272172998621
+      0.01303636840598877
+    0.0009886707094704543
+      -0.1113628194665092
+       0.4545342641330058
+ 7.96e+10    
+       0.4556594574866326
+      -0.1118097314790442
+       0.4930233649358922
+     0.001453556852013081
+     -0.07200787422585508
+        0.493198695300666
+      0.01314553331983414
+     0.001414910650954124
+      -0.1117208978214087
+       0.4554679009493443
+ 8.01e+10    
+       0.4565628647229207
+      -0.1121555344711571
+       0.4944690448347097
+     0.001893282125537794
+     -0.07275290186282402
+       0.4946461507100927
+      0.01324565035306046
+     0.001852384098470363
+       -0.112066964665134
+       0.4563726699152341
+ 8.06e+10    
+       0.4574373632773084
+      -0.1124892447759686
+       0.4958906748906899
+     0.002344068466061001
+     -0.07350691363845005
+       0.4960696646398708
+      0.01333653151963713
+     0.002301075240062326
+      -0.1124009949869413
+       0.4572485837374377
+ 8.11e+10    
+       0.4582829626420893
+      -0.1128108305017718
+       0.4972883230371963
+     0.002805892487941648
+     -0.07427003653519768
+       0.4974693082465673
+      0.01341799273060474
+     0.002760960058823673
+      -0.1127229577710013
+       0.4580956523455392
+ 8.16e+10    
+       0.4590996694517608
+      -0.1131202533349123
+       0.4986620470424246
+     0.003278722616900442
+     -0.07504237912770031
+       0.4988451423488368
+      0.01348985416041385
+     0.003232006060743987
+       -0.113032815536137
+       0.4589138828089084
+ 8.21e+10    
+       0.4598874874061783
+      -0.1134174680848073
+       0.5000118941481997
+     0.003762518800298325
+      -0.0758240309348989
+       0.5001972170620773
+      0.01355194062723235
+      0.00371417199343313
+      -0.1133305238808303
+       0.4597032792601888
+ 8.26e+10    
+       0.4606464172005243
+      -0.1137024222351177
+       0.5013379007239603
+     0.004257232209264332
+     -0.07661506178751727
+       0.5015255714502711
+      0.01360408198697282
+     0.004207407556947896
+      -0.1136160310351892
+       0.4604638428257418
+ 8.31e+10    
+       0.4613764564623692
+      -0.1139750555028178
+       0.5026400919393132
+     0.004762804934098881
+     -0.07741552121163238
+       0.5028302331942093
+      0.01364611353884946
+     0.004711653107079942
+      -0.1138892774195506
+       0.4611955715629185
+ 8.36e+10    
+       0.4620775996952061
+       -0.114235299404436
+       0.5039184814516067
+     0.005279169674428929
+     -0.07822543783060391
+        0.504111218277089
+      0.01367787644114602
+     0.005226839354062238
+      -0.1141501952114744
+       0.4618984604039137
+ 8.41e+10    
+        0.462749838229198
+      -0.1144830768319716
+        0.505173071112238
+     0.005806249424663503
+     -0.07904481878426808
+       0.5053685306875683
+      0.01369921813584758
+     0.005752887056218036
+      -0.1143987079216395
+       0.4625725011068627
+ 8.46e+10    
+       0.4633931601785204
+      -0.1147183016377608
+       0.5064038506882017
+     0.006343957156746684
+     -0.07987364916778721
+       0.5066021621398864
+      0.01370999278018831
+     0.006289706710851771
+      -0.1146347299792422
+       0.4632176822133044
+ 8.51e+10    
+       0.4640075504057516
+      -0.1149408782305093
+         0.50761079760273
+     0.006892195500701589
+     -0.08071189149029617
+        0.507812091811599
+      0.01371006168425297
+     0.006837198243309339
+       -0.114858166328183
+       0.4638339890128301
+ 8.56e+10    
+       0.4645929904932493
+      -0.1151507011825589
+       0.5087938766922224
+     0.007450856424382127
+     -0.08155948515431691
+       0.5089982860990354
+      0.01369929375272826
+     0.007395250695130366
+      -0.1150689120346308
+       0.4644214035144444
+ 8.61e+10    
+       0.4651494587213565
+      -0.1153476548494289
+       0.5099530399809649
+     0.008019820913387495
+     -0.08241634595682766
+       0.5101606983907128
+      0.01367756592986736
+     0.007963741912535294
+      -0.1152668519071771
+       0.4649799044250366
+ 8.66e+10    
+       0.4656769300537429
+       -0.115531613002656
+       0.5110882264733854
+     0.008598958652373279
+     -0.08328236561229491
+       0.5112992688576956
+      0.01364476364559122
+     0.008542538236450476
+      -0.1154518601298309
+       0.4655094671346649
+ 8.71e+10    
+       0.4661753761297931
+      -0.1157024384769199
+       0.5121993619645225
+     0.009188127708471374
+     -0.08415741129975782
+       0.5124139242638335
+       0.0136007812622355
+     0.009131494195092443
+      -0.1156237999099499
+       0.4660100637089959
+ 8.76e+10    
+       0.4666447652642701
+      -0.1158599828323025
+       0.5132863588683311
+      0.00978717421859162
+     -0.08504132523368087
+       0.5135045777923295
+      0.01354552251991226
+     0.009730452200066356
+      -0.1157825231404858
+       0.4664816628887192
+ 8.81e+10    
+        0.467085062454057
+      -0.1160040860326056
+       0.5143491160639742
+      0.01039593208069562
+     -0.08593392425964454
+       0.5145711288923465
+       0.0134789009799211
+       0.0103392422470809
+      -0.1159278700792533
+       0.4669242300964525
+ 8.86e+10    
+       0.4674962293922475
+      -0.1161345761404859
+       0.5153875187603773
+      0.01101422265040507
+     -0.08683499947589304
+       0.5156134631427157
+      0.01340084046402923
+      0.01095768162213626
+      -0.1160596690443426
+        0.467337727450448
+ 8.91e+10    
+       0.4678782244898194
+      -0.1162512690312505
+       0.5164014383802822
+      0.01164185444461402
+     -0.08774431588244275
+       0.5166314521362434
+      0.01331127548948678
+      0.01158557461504839
+      -0.1161777361287655
+       0.4677221137861776
+ 8.96e+10    
+       0.4682310029046868
+       -0.116353968125236
+        0.517390732462008
+      0.01227862285197162
+     -0.08866161205667832
+       0.5176249533815288
+       0.0132101516979767
+      0.01222271223940785
+      -0.1162818749332034
+       0.4680773446849964
+ 9.01e+10    
+       0.4685545165784315
+      -0.1164424641406034
+       0.5183552445813054
+      0.01292430985204992
+     -0.08958659985862984
+        0.518593810224766
+      0.01309742627728659
+      0.01286887196233596
+      -0.1163718763195249
+       0.4684033725107459
+ 9.06e+10    
+       0.4688487142809504
+      -0.1165165348671449
+       0.5192948042913728
+       0.0135786837435148
+     -0.09051896416474867
+       0.5195378517914743
+      0.01297306837538945
+      0.01352381744315844
+      -0.1164475181853822
+       0.4687001464537962
+ 9.11e+10    
+       0.4691135416628254
+      -0.1165759449624584
+       0.5202092270839379
+      0.01424149888326685
+     -0.09145836263327206
+       0.5204568929472159
+      0.01283705950471474
+       0.0141872982826056
+      -0.1165085652608697
+       0.4689676125831821
+ 9.16e+10    
+       0.4693489413159908
+      -0.1166204457712463
+       0.5210983143688594
+      0.01491249543608644
+     -0.09240442550008605
+       0.5213507342796693
+      0.01268939393667204
+      0.01485904978401772
+      -0.1165547689290087
+       0.4692057139067836
+ 9.21e+10    
+       0.4695548528425239
+      -0.1166497751694444
+       0.5219618534755035
+      0.01559139913701673
+      -0.0933567554071167
+       0.5222191620994144
+      0.01253007908491437
+       0.0155387927262185
+      -0.1165858670700117
+        0.469414390439482
+ 9.26e+10    
+        0.469731212931891
+      -0.1166636574331346
+        0.522799617672541
+      0.01627792106675278
+     -0.09431492726448416
+       0.5230619484638329
+      0.01235913587653153
+      0.01622623315019021
+      -0.1166015839317816
+       0.4695935792800513
+ 9.31e+10    
+       0.4698779554469358
+       -0.116661803135143
+        0.523611366211719
+      0.01697175744114594
+     -0.09527848814700575
+       0.5238788512201493
+       0.0121765991097634
+      0.01692106216034592
+      -0.1166016300265294
+       0.4697432146963021
+ 9.36e+10    
+        0.469995011518499
+      -0.1166439090683595
+       0.5243968443899271
+      0.01767258941582034
+     -0.09624695722544868
+        0.524669614071172
+       0.0119825177986164
+      0.01762295574000233
+      -0.1165857020555465
+       0.4698632282192812
+ 9.41e+10    
+       0.4700823096492918
+      -0.1166096581988133
+       0.5251557836352849
+      0.01838008290655508
+     -0.09721982573479708
+        0.525433966662642
+      0.01177695550169154
+      0.01833157458415467
+      -0.1165534828627375
+       0.4699535487463252
+ 9.46e+10    
+       0.4701397758268962
+      -0.1165587196482019
+       0.5258879016140043
+      0.01909388842688736
+     -0.09819655698002436
+       0.5261716246930898
+      0.01155999063619604
+      0.01904656394840935
+      -0.1165046414183514
+       0.4700141026532995
+ 9.51e+10    
+       0.4701673336462908
+      -0.1164907487081475
+       0.5265929023608701
+      0.01981364094349443
+     -0.09917658638002703
+       0.5268822900467499
+       0.0113317167746658
+      0.01976755351634808
+      -0.1164388328340082
+       0.4700448139165608
+ 9.56e+10    
+       0.4701649044422934
+      -0.1164053868865763
+       0.5272704764319169
+      0.02053895975010571
+       -0.100159321551256
+       0.5275656509494705
+      0.01109224292518662
+       0.0204941572856449
+      -0.1163556984100603
+        0.470045604244396
+ 9.61e+10    
+       0.4701324074317247
+      -0.1163022619878356
+       0.5279203010817984
+      0.02126944836158362
+      -0.1011441424322512
+       0.5282213821476858
+      0.01084169379251301
+      0.02122597347389483
+      -0.1162548657161947
+       0.4700163932183483
+ 9.66e+10    
+       0.4700697598661661
+        -0.11618098822742
+       0.5285420404639412
+       0.0220046944283834
+      -0.1021304014497661
+       0.5288491451145527
+      0.01058021002131053
+      0.02196258444522967
+       -0.116135948707991
+       0.4699570984453798
+ 9.71e+10    
+       0.4699768771951871
+      -0.1160411663829637
+       0.5291353458568699
+      0.02274426967271349
+      -0.1031174237280769
+       0.5294485882770203
+       0.0103079484190532
+      0.02270355665859084
+      -0.1159985478779228
+       0.4698676357197888
+ 9.76e+10    
+       0.4698536732401793
+      -0.1158823839817973
+       0.5296998559138012
+      0.02348772984710604
+      -0.1041045073414893
+       0.5300193472712109
+      0.01002508215833555
+      0.02344844063842467
+      -0.1158422504445236
+        0.469747919196531
+ 9.81e+10    
+       0.4697000603797436
+      -0.1157042155275021
+       0.5302351969401184
+      0.02423461471697907
+      -0.1050909236133772
+       0.5305610452226275
+     0.009731800958711409
+      0.02419677096899111
+      -0.1156666305794422
+       0.4695978615753305
+ 9.86e+10    
+       0.4695159497462241
+      -0.1155062227653506
+       0.5307409831954915
+      0.02498444806682466
+      -0.1060759174601032
+       0.5310732930531249
+     0.009428311245709113
+      0.02494806631290276
+      -0.1154712496739939
+       0.4694173742963948
+ 9.91e+10    
+       0.4693012514341121
+      -0.1152879549887553
+        0.531216817223548
+       0.0257367377327276
+      -0.1070587077834262
+       0.5315556898149564
+     0.009114836287972319
+      0.02570182945496371
+       -0.115255656646684
+       0.4692063677479201
+ 9.96e+10    
+       0.4690558747204144
+       -0.115048949387141
+       0.5316622902092617
+       0.0264909756604046
+      -0.1080384879106064
+       0.5320078230525699
+     0.008791616310076768
+      0.02645754737239138
+      -0.1150193882917584
+        0.468964751485247
+ 1.001e+11   
+       0.4687797282975171
+      -0.1147887314370486
+       0.5320769823636424
+         0.02724663799096
+      -0.1090144260847363
+       0.5324292691924924
+     0.008458908582029159
+      0.02721469133176647
+      -0.1147619696713243
+       0.4686924344628531
+ 1.006e+11   
+       0.4684727205186097
+      -0.1145068153370218
+       0.5324604633381262
+      0.02800318517478125
+      -0.1099856660058135
+        0.532819593962907
+     0.008116987483169016
+      0.02797271701452386
+      -0.1144829145511411
+       0.4683893252786178
+ 1.011e+11   
+       0.4681347596560738
+      -0.1142027044876253
+       0.5328122926675346
+      0.02876006211458045
+      -0.1109513274233334
+       0.5331783528419457
+     0.007766144540657724
+      0.02873106467106751
+      -0.1141817258815856
+       0.4680553324313405
+ 1.016e+11   
+       0.4677657541734179
+       -0.113875892017629
+       0.5331320202431622
+      0.02951669833828209
+      -0.1119105067823121
+        0.533505091536817
+     0.007406688442085124
+       0.0294891593047056
+      -0.1138578963247287
+       0.4676903645914141
+ 1.021e+11   
+       0.4673656130103775
+       -0.113525861357483
+       0.5334191868166487
+      0.03027250820363573
+      -0.1128622779234301
+       0.5337993464928806
+     0.007038945019764482
+      0.03024641088652331
+      -0.1135109088283607
+       0.4672943308850774
+ 1.026e+11   
+       0.4669342458824036
+      -0.1131520868607121
+       0.5336733245350042
+      0.03102689113379142
+      -0.1138056928381479
+        0.534060645435635
+     0.006663257208682626
+      0.03100221460178634
+      -0.1131402372484726
+       0.4668671411925249
+ 1.031e+11   
+       0.4664715635938448
+      -0.1127540344744308
+       0.5338939575063135
+      0.03177923188646663
+      -0.1147397824796626
+       0.5342885079433306
+     0.006279984974657911
+      0.03175595112886745
+      -0.1127453470207458
+       0.4664087064604175
+ 1.036e+11   
+       0.4659774783659162
+      -0.1123311624600708
+       0.5340806023999118
+      0.03252890085653812
+      -0.1156635576320923
+       0.5344824460524776
+     0.005889505214226572
+      0.03250698695157977
+      -0.1123256958816451
+       0.4659189390285772
+ 1.041e+11   
+       0.4654519041793387
+      -0.1118829221647121
+       0.5342327690765643
+      0.03327525441313198
+      -0.1165760098363464
+       0.5346419648967308
+     0.005492211623688487
+       0.0332546747056764
+      -0.1118807346406995
+       0.4653977529714178
+ 1.046e+11   
+       0.4648947571318102
+      -0.1114087588440196
+       0.5343499612546766
+      0.03401763527274913
+      -0.1174761123767282
+       0.5347665633801467
+      0.00508851453826252
+        0.033998353560691
+      -0.1114099080044362
+       0.4648450644546701
+ 1.051e+11   
+       0.4643059558106352
+      -0.1109081125376075
+       0.5344316772085873
+       0.0347553729077316
+      -0.1183628213257588
+       0.5348557348828719
+     0.004678840739374026
+      0.03473734963714782
+      -0.1109126554519965
+       0.4642607921068641
+ 1.056e+11   
+       0.4636854216809476
+      -0.1103804189972478
+       0.5344774105022342
+      0.03548778399276886
+      -0.1192350766511928
+       0.5349089680030734
+     0.004263633230343591
+      0.03547097646092003
+       -0.110388412164211
+       0.4636448574063243
+ 1.061e+11   
+       0.4630330794893324
+       -0.109825110668754
+       0.5344866507567272
+      0.03621417288871675
+      -0.1200918033834231
+       0.5349257473334962
+     0.003843350979080806
+      0.03619853545480151
+      -0.1098366100061095
+       0.4629971850839376
+ 1.066e+11   
+       0.4623488576830223
+      -0.1092416177274936
+        0.534458884453851
+      0.03693383216513936
+      -0.1209319128453079
+       0.5349055542729058
+     0.003418468627599692
+       0.0369193164680244
+       -0.109256678563132
+       0.4623177035414401
+ 1.071e+11   
+       0.4616326888450282
+      -0.1086293691683834
+        0.534393595774122
+       0.0376460431623114
+       -0.121754303945391
+       0.5348478678742944
+     0.002989476167864103
+      0.03763259834495142
+      -0.1086480462316946
+       0.4616063452853801
+ 1.076e+11   
+       0.4608845101451947
+      -0.1079877939506206
+       0.5342902674711207
+      0.03835007659278683
+      -0.1225578645324902
+       0.5347521657279714
+     0.002556878582597569
+      0.03833764953282249
+       -0.108010141364283
+       0.4608630473772039
+ 1.081e+11   
+        0.460104263806886
+      -0.1073163221969608
+       0.5341483817816529
+      0.03904519318392149
+      -0.1233414728158778
+       0.5346179248820034
+     0.002121195451661973
+        0.039033728729594
+       -0.107342393469444
+       0.4600877518991933
+ 1.086e+11   
+       0.4592918975897617
+      -0.1066143864477008
+       0.5339674213708503
+      0.03973064436113378
+      -0.1241039988475426
+       0.5344446227982489
+     0.001682960522572479
+       0.0397200855724078
+      -0.1066442344662434
+       0.4592804064360369
+ 1.091e+11   
+       0.4584473652880424
+       -0.105881422969311
+       0.5337468703149792
+      0.04040567297274424
+      -0.1248443060693027
+       0.5342317383442952
+     0.001242721244751461
+       0.0403959613668021
+      -0.1059150999931445
+       0.4584409645724373
+ 1.096e+11   
+       0.4575706272448131
+      -0.1051168731175399
+        0.533486215118014
+      0.04106951405677006
+      -0.1255612529231741
+       0.5339787528233721
+    0.0008010382678413971
+      0.04106058985737512
+      -0.1051544307720292
+       0.4575693864064405
+ 1.101e+11   
+        0.456661650881169
+      -0.1043201847540265
+       0.5331849457653989
+      0.04172139564965428
+      -0.1262536945254496
+       0.5336851510374273
+    0.0003584849029050303
+      0.04171319803977323
+      -0.1043616740247672
+       0.4566656390778327
+ 1.106e+11   
+       0.4557204112412593
+      -0.1034908137169383
+       0.5328425568120481
+      0.04236053963788747
+      -0.1269204844046421
+       0.5333504223891171
+   -8.435345397855409e-05
+      0.04235300701508286
+      -0.1035362849442668
+       0.4557296973121221
+ 1.111e+11   
+       0.4547468915513039
+      -0.1026282253432511
+       0.5324585485057918
+      0.04298616265155712
+      -0.1275604763012391
+       0.5329740620160995
+   -0.0005268799344769716
+      0.04297923288520173
+      -0.1026777282174722
+       0.4547615439792477
+ 1.116e+11   
+       0.4537410837937537
+      -0.1017318960433316
+       0.5320324279449601
+      0.04359747700062768
+      -0.1281725260305775
+        0.532555571962312
+   -0.0009684868495853471
+      0.04359108769102568
+       -0.101785479599931
+       0.4537611706665323
+ 1.121e+11   
+       0.4527029892948541
+      -0.1008013149256318
+       0.5315637102689655
+       0.0441936916536841
+      -0.1287554934056806
+        0.532094462381852
+    -0.001408556377750684
+      0.04418778039164188
+      -0.1008590275409962
+        0.452728578265944
+ 1.126e+11   
+       0.4516326193256257
+     -0.09983598547016415
+       0.5310519198821307
+       0.0447740132587254
+      -0.1293082442211664
+       0.5315902527761275
+    -0.001846461292022066
+      0.04476851788547245
+     -0.09989787485755498
+       0.4516637775741585
+ 1.131e+11   
+       0.4505299957154923
+     -0.09883542724982916
+       0.5304965917086746
+      0.04533764720568192
+      -0.1298296522953164
+       0.5310424732631305
+     -0.00228156572345418
+      0.04533250607252924
+     -0.09890154045563676
+       0.4505667899057401
+ 1.136e+11   
+       0.4493951514775429
+     -0.09779917769664595
+       0.5298972724778188
+      0.04588379872993239
+      -0.1303186015680198
+       0.5304506658772903
+    -0.002713225963173953
+      0.04587895095669012
+     -0.09786956109689521
+       0.4494376477178593
+ 1.141e+11   
+        0.448228131444729
+     -0.09672679391184184
+       0.5292535220382197
+      0.04641167405682099
+      -0.1307739882561779
+       0.5298143858988696
+    -0.003140791301077913
+      0.04640705978884611
+     -0.09680149320897194
+       0.4482763952459333
+ 1.146e+11   
+       0.4470289929158691
+      -0.0956178545165389
+        0.528564914698762
+      0.04692048158531546
+      -0.1311947230588312
+       0.5291332032101945
+    -0.003563604901436534
+      0.04691604224794434
+     -0.09569691473661023
+       0.4470830891492094
+ 1.151e+11   
+       0.4457978063102525
+     -0.09447196154063435
+       0.5278310405950279
+        0.047409433110121
+      -0.1315797334146158
+       0.5284067036781631
+    -0.003981004714528148
+      0.04740511166074633
+     -0.09455542703053646
+       0.4458577991650511
+ 1.156e+11   
+       0.4445346558296979
+     -0.09328874234728428
+       0.5270515070790572
+      0.04787774508208816
+       -0.131927965806259
+       0.5276344905600151
+    -0.004392324424454233
+      0.04787348625796053
+     -0.09337665677215079
+       0.4446006087704397
+ 1.161e+11   
+       0.4432396401263251
+     -0.09206785158844495
+       0.5262259401290431
+      0.04832463990303289
+      -0.1322383881079524
+       0.5268161859299093
+    -0.004796894431575476
+      0.04832039046570077
+      -0.0921602579297576
+       0.4433116158499126
+ 1.166e+11   
+       0.4419128729750005
+     -0.09080897318974245
+       0.5253539857780917
+      0.04874934725602636
+      -0.1325099919750342
+       0.5259514321245964
+    -0.005194042868485387
+      0.04874505623070263
+     -0.09090591374291931
+       0.4419909333672763
+ 1.171e+11   
+       0.4405544839479659
+     -0.08951182235800084
+       0.5244353115566648
+      0.04915110546710487
+      -0.1327417952686905
+       0.5250398932040712
+    -0.005583096648897726
+       0.0491467243766167
+      -0.0896133387311694
+       0.4406386900406384
+ 1.176e+11   
+       0.4391646190905003
+     -0.08817614760977877
+       0.5234696079482082
+      0.04952916289755535
+      -0.1329328445133733
+       0.5240812564237323
+    -0.005963382548366888
+      0.04952464599038613
+     -0.08828228072189644
+       0.4392550310175732
+ 1.181e+11   
+       0.4377434415950666
+     -0.08680173281410336
+       0.5224565898522581
+      0.04988277936346532
+      -0.1330822173818171
+       0.5230752337169267
+    -0.006334228314484385
+      0.04987808383545311
+     -0.08691252289392372
+       0.4378401185495012
+ 1.186e+11   
+       0.4362911324717884
+     -0.08538839924495305
+       0.5213959980522217
+      0.05021122758066679
+      -0.1331890252013981
+        0.522021563180232
+    -0.006694963805823385
+      0.05020631378944422
+     -0.08550388583012251
+         0.43639413266234
+ 1.191e+11   
+       0.4348078912130598
+     -0.08393600763801838
+       0.5202876006832178
+      0.05051379463149098
+      -0.1332524154774872
+       0.5209200105604117
+    -0.007044922157009311
+      0.05050862630308026
+     -0.08405622957408024
+       0.4349172718208943
+ 1.196e+11   
+       0.4332939364491641
+     -0.08244446024509361
+       0.5191311946954533
+      0.05078978345010458
+      -0.1332715744260383
+       0.5197703707366954
+    -0.007383440968449101
+      0.05078432787745334
+     -0.08256945568536819
+       0.4334097535853799
+ 1.201e+11   
+        0.431749506592869
+     -0.08091370288008091
+       0.5179266073082178
+      0.05103851432317385
+      -0.1332457295097845
+       0.5185724691941306
+    -0.007709863518199892
+      0.05103274255571049
+     -0.08104350928546966
+       0.4318718152557217
+ 1.206e+11   
+       0.4301748604690585
+     -0.07934372694938786
+       0.5166736974491046
+      0.05125932640144759
+      -0.1331741519700156
+       0.5173261634816103
+    -0.008023539993445445
+      0.05125321342523376
+     -0.07947838108839994
+       0.4303037145019731
+ 1.211e+11   
+       0.4285702779269177
+      -0.0777345714590439
+       0.5153723571732695
+      0.05145157921869865
+      -0.1330561593473628
+       0.5160313446505985
+    -0.008323828738629991
+      0.05144510412670592
+     -0.07787410940833854
+       0.4287057299769942
+ 1.216e+11   
+       0.4269360604308662
+     -0.07608632499073978
+       0.5140225130544406
+      0.05161465421228585
+      -0.1328911179799508
+       0.5146879386663269
+    -0.008610097517928824
+      0.05160780036401742
+     -0.07623078213600587
+       0.4270781619079198
+ 1.221e+11   
+       0.4252725316265843
+     -0.07439912763821696
+       0.5126241275447512
+      0.05174795624181679
+      -0.1326784454744617
+       0.5132959077859305
+    -0.008881724788133372
+      0.05174071141206105
+     -0.07454853867518861
+       0.4254213326630458
+ 1.226e+11   
+       0.4235800378783425
+     -0.07267317289468797
+       0.5111772002920798
+      0.05185091509923323
+      -0.1324176131360859
+       0.5118552518962327
+    -0.009138100978709256
+      0.05184327161493094
+     -0.07282757183062658
+       0.4237355872897917
+ 1.231e+11   
+       0.4218589487734942
+     -0.07090870948205868
+       0.5096817694110104
+      0.05192298700496814
+      -0.1321081483494544
+       0.5103660098030796
+    -0.009378629775121539
+      0.05191494187041935
+     -0.07106812963760192
+       0.4220212940204113
+ 1.236e+11   
+       0.4201096575897293
+     -0.06910604311132552
+       0.5081379126970799
+        0.051963656084945
+      -0.1317496368992034
+       0.5088282604651381
+    -0.009602729402548704
+      0.05195521109406116
+     -0.06927051712248641
+       0.4202788447399856
+ 1.241e+11   
+       0.4183325817203995
+     -0.06726553816333615
+       0.5065457487763024
+      0.05197243582004653
+      -0.1313417252173862
+       0.5072421241621895
+    -0.009809833902881397
+      0.05196359765560511
+     -0.06743509798426693
+       0.4185086554132537
+ 1.246e+11   
+       0.4165281630533277
+      -0.0653876192791368
+       0.5049054381819484
+      0.05194887046289758
+      -0.1308841225467586
+       0.5056077635896348
+    -0.009999394403868956
+      0.05193965078223648
+     -0.06556229618476762
+       0.4167111664644262
+ 1.251e+11   
+       0.4146968682978258
+     -0.06347277284696234
+       0.5032171843473251
+      0.05189253641326377
+      -0.1303766030055813
+       0.5039253848703197
+     -0.01017088037306567
+      0.05188295191990529
+     -0.06365259743631918
+       0.4148868431057352
+ 1.256e+11   
+       0.4128391892546101
+     -0.06152154837423381
+       0.5014812345065034
+      0.05180304354515933
+      -0.1298190075405713
+       0.5021952384712444
+     -0.01032378085265597
+       0.0517931160456637
+     -0.06170655057394372
+       0.4130361756089376
+ 1.261e+11   
+       0.4109556430230495
+     -0.05953455973026661
+       0.4996978804896758
+      0.05168003647650746
+      -0.1292112457536762
+       0.5004176200169855
+     -0.01045760566872558
+      0.05166979292248548
+      -0.0597247687985494
+       0.4111596795141126
+ 1.266e+11   
+       0.4090467721401046
+     -0.05751248624686883
+       0.4978674594050112
+      0.05152319577304205
+      -0.1285532975858254
+        0.498592870986462
+     -0.01057188660980127
+      0.05151266828774037
+     -0.05770793077764236
+       0.4092578957704642
+ 1.271e+11   
+       0.4071131446445105
+     -0.05545607366140566
+       0.4959903541925754
+      0.05133223907782124
+      -0.1278452148437817
+       0.4967213792825728
+     -0.01066617856933777
+      0.05132146496656165
+     -0.05565678158898112
+       0.4073313908024612
+ 1.276e+11   
+       0.4051553540605055
+     -0.05336613488808949
+       0.4940669940401236
+      0.05110692215537081
+      -0.1270871225499944
+       0.4948035796610487
+      -0.0107400606436439
+      0.05109594389986288
+     -0.05357213349167283
+       0.4053807564954937
+ 1.281e+11   
+       0.4031740192939086
+     -0.05124355060063476
+       0.4920978546457866
+        0.050847039841961
+      -0.1262792201014438
+       0.4928399540073535
+     -0.01079313718105489
+      0.05083590507753286
+     -0.05145486650964467
+        0.403406610094342
+ 1.286e+11   
+       0.4011697844342907
+     -0.04908926961073797
+       0.4900834583157573
+      0.05055242688976529
+      -0.1254217822142039
+       0.4908310314450376
+     -0.01082503877368034
+      0.05054118836594913
+     -0.04930592881004908
+        0.401409594007635
+ 1.291e+11   
+       0.3991433184561508
+     -0.04690430902502252
+       0.4880243738820116
+      0.05022295869540431
+       -0.124515159637866
+        0.488777388264087
+     -0.01083542318451331
+      0.05021167421844075
+     -0.04712633686044923
+       0.3993903755115045
+ 1.296e+11   
+       0.3970953148117097
+     -0.04468975416260234
+       0.4859212164255219
+      0.04985855190059921
+      -0.1235597796186463
+       0.4866796476526715
+     -0.01082397620411299
+      0.04984728425849836
+     -0.04491717534644062
+       0.3973496463450371
+ 1.301e+11   
+       0.3950264909083235
+     -0.04244675821522639
+       0.4837746467901892
+      0.04945916485326512
+      -0.1225561460885638
+       0.4845384792176312
+     -0.01079041242649356
+      0.04944798172221017
+     -0.04267959683189083
+       0.3952881221904488
+ 1.306e+11   
+       0.3929375874625082
+     -0.04017654163077258
+       0.4815853708696016
+      0.04902479791624094
+      -0.1215048395599287
+       0.4823545982768531
+     -0.01073447593781771
+      0.04901377174898525
+     -0.04041482114272221
+       0.3932065420302399
+ 1.311e+11   
+       0.3908293677231779
+     -0.03788039120100314
+        0.479354138652613
+      0.04855549361183422
+      -0.1204065167023657
+       0.4801287649079061
+     -0.01065594090923668
+      0.04854470150698179
+     -0.03812413445446761
+        0.391105667373393
+ 1.316e+11   
+       0.3887026165562631
+     -0.03555965883337116
+       0.4770817430092487
+       0.0480513365880584
+      -0.1192619095776798
+       0.4778617827338624
+     -0.01055461208420382
+      0.04804086014035542
+     -0.03580888806383126
+       0.3889862813432282
+ 1.321e+11   
+       0.3865581393821263
+      -0.0332157599860706
+       0.4747690181982093
+      0.04751245339368961
+      -0.1180718245093621
+       0.4755544974299533
+     -0.01043032515349902
+      0.04750237852541411
+     -0.03347049682403595
+       0.3868491876184583
+ 1.326e+11   
+       0.3843967609583993
+     -0.03085017174574067
+       0.4724168380797232
+      0.04693901204733041
+      -0.1168371405597566
+        0.473207794931816
+     -0.01028294700570323
+      0.04692942882002631
+     -0.03111043722187082
+       0.3846952092194329
+ 1.331e+11   
+       0.3822193239994584
+     -0.02846443052588998
+       0.4700261140132776
+      0.04633122138736114
+      -0.1155588075910888
+       0.4708225993262158
+     -0.01011237584716375
+      0.04632222379431918
+      -0.0287302450761409
+       0.3825251871315072
+ 1.336e+11   
+       0.3800266876245127
+     -0.02606012936423834
+       0.4675977924200981
+      0.04568933018667426
+      -0.1142378438805158
+       0.4683998704038426
+    -0.009918541178875973
+      0.04568101592624145
+     -0.02633151283481716
+       0.3803399787570048
+ 1.341e+11   
+        0.377819725625913
+      -0.0236389147969534
+       0.4651328519927371
+      0.04501362601904264
+      -0.1128753332649485
+        0.465940600854873
+    -0.009701403623375357
+      0.04500609624802836
+     -0.02391588644836539
+       0.3781404561876235
+ 1.346e+11   
+       0.3755993245492398
+     -0.02120248328663509
+       0.4626323005279328
+      0.04430443385957834
+       -0.111472421784167
+        0.463445813086217
+    -0.009460954588406846
+      0.04429779292798529
+     -0.02148506179789006
+       0.3759275042889279
+ 1.351e+11   
+       0.3733663815774236
+     -0.01875257718191568
+       0.4600971713646169
+      0.04356211440636606
+      -0.1100303137962112
+       0.4609165556382076
+    -0.009197215761309014
+      0.04355646957292249
+     -0.01904078065368062
+       0.3737020185886633
+ 1.356e+11   
+       0.3711218022098167
+     -0.01629098018486725
+        0.457528519401758
+      0.04278706210538676
+      -0.1085502675326822
+       0.4583538991793702
+    -0.008910238419412521
+      0.04278252323409693
+     -0.01658482614242948
+       0.3714649029606419
+ 1.361e+11   
+       0.3688664977290819
+     -0.01381951230405812
+       0.4549274166784137
+       0.0419797028643349
+      -0.1070335900666451
+       0.4557589320575421
+    -0.008600102550729285
+       0.0419763821033113
+     -0.01411901769963106
+       0.3692170670964154
+ 1.366e+11   
+       0.3666013824474095
+      -0.0113400242695889
+       0.4522949474887666
+      0.04114049143911136
+      -0.1054816316603065
+       0.4531327553833823
+    -0.008266915771408697
+      0.04113850288099756
+      -0.0116452054838352
+       0.3669594237563711
+ 1.371e+11   
+       0.3643273707248211
+    -0.008854391387539367
+       0.4496322030130991
+      0.04026990847626891
+      -0.1038957794629553
+       0.4504764776234491
+    -0.007910812030654491
+      0.04026936780225762
+    -0.009165264230563044
+       0.3646928857931379
+ 1.376e+11   
+       0.3620453737517291
+    -0.006364506811085731
+       0.4469402754387074
+      0.03936845719688337
+      -0.1022774505277425
+       0.4477912086804284
+     -0.00753195009312679
+      0.03936948130371881
+    -0.006681086522711151
+       0.3624183629395636
+ 1.381e+11   
+       0.3597562960894775
+     -0.00387227420615733
+       0.4442202515486758
+      0.03843665970487107
+      -0.1006280841151202
+       0.4450780534349288
+    -0.007130511789020741
+      0.03843936631701143
+    -0.004194575455601614
+       0.3601367583546256
+ 1.386e+11   
+       0.3574610319616052
+    -0.001379599789916493
+       0.4414732057546953
+      0.03747505290442722
+     -0.09894913325234338
+       0.4423381047269339
+    -0.006706700019902622
+      0.03747956017165409
+    -0.001707636674875682
+       0.3578489649203558
+ 1.391e+11   
+       0.3551604612905375
+     0.001111616278638315
+       0.4387001925500286
+         0.03648418401159
+     -0.09724205551769187
+       0.4395724357516316
+    -0.006260736512004365
+      0.03649061009349379
+    0.0007778302336935231
+       0.3555558612841436
+ 1.396e+11   
+        0.352855445473464
+     0.003599489176553119
+       0.4359022383588703
+       0.0354646056442685
+     -0.09550830301736535
+       0.4367820918462338
+    -0.005792859307747888
+      0.03547306828354121
+     0.003259941022237317
+       0.3532583076409305
+ 1.401e+11   
+       0.3505468228936554
+     0.006082159381536618
+       0.4330803327583993
+      0.03441687047698323
+      -0.0937493115252535
+        0.433968081644445
+    -0.005303319983526758
+      0.03442748656192842
+     0.005736836746017684
+       0.3509571412501515
+ 1.406e+11   
+       0.3482354041626946
+     0.008557803341067401
+       0.4302354190523894
+      0.03334152544538222
+     -0.09196648875566876
+       0.4311313675746139
+    -0.004792380587814033
+      0.03335441056501431
+     0.008206694432661256
+       0.3486531716845391
+ 1.411e+11   
+       0.3459219670908785
+       0.0110246448619614
+       0.4273683841697835
+      0.03223910548852769
+     -0.09016120173893391
+       0.4282728556793733
+     -0.00426031028915209
+      0.03225437348068702
+      0.01066773847202622
+       0.3463471758066746
+ 1.416e+11   
+       0.3436072513841933
+      0.01348096723472735
+       0.4244800478703623
+      0.03111012681530191
+     -0.08833476327251526
+       0.4253933847341828
+    -0.003707381725932806
+      0.03112788931132426
+      0.01311825274001415
+       0.3440398924724193
+ 1.421e+11   
+       0.3412919530667996
+      0.01592512610339918
+       0.4215711512344401
+      0.02995507968520323
+     -0.08648841742174143
+       0.4224937146441635
+     -0.00313386705197595
+      0.02997544565247888
+      0.01555659346860301
+        0.341732016959985
+ 1.426e+11   
+       0.3389767186301975
+      0.01835556309155431
+       0.4186423444168844
+      0.02877442069227466
+     -0.08462332404420569
+       0.4195745140989125
+    -0.002540033670531852
+      0.02879749597781243
+      0.01798120287072744
+       0.3394241951257493
+ 1.431e+11   
+       0.3366621389112184
+      0.02077082018935346
+       0.4156941736482547
+       0.0275685645444569
+     -0.08274054231694244
+       0.4166363474675617
+    -0.001926139650134315
+      0.02759445142224132
+      0.02039062352675922
+       0.3371170172888428
+ 1.436e+11   
+       0.3343487427028097
+      0.02316955490537345
+       0.4127270674654165
+      0.02633787533161659
+     -0.08084101324574622
+       0.4136796609166535
+     -0.00129242881981507
+      0.02636667205657327
+      0.02278351353469858
+       0.3348110118486893
+ 1.441e+11   
+       0.3320369901039611
+      0.02555055618141818
+       0.4097413221587404
+       0.0250826572771508
+     -0.07892554114039302
+       0.4107047677383208
+   -0.0006391255385214179
+      0.02511445764879529
+      0.02515866242368918
+       0.3325066386415289
+ 1.446e+11   
+       0.3297272656166683
+      0.02791276106560268
+       0.4067370864242215
+      0.02380314497139603
+      -0.0769947740443694
+       0.4077118328760207
+     3.35708622484492e-05
+      0.02383803791086363
+      0.02751500782460339
+       0.3302042820441861
+ 1.451e+11   
+        0.327419871000927
+      0.03025527213241629
+       0.4037143452130275
+      0.02249949308691634
+     -0.07504918311005888
+       0.4047008566415776
+    0.0007254919629891357
+      0.02253756223062203
+      0.02985165288766198
+       0.3279042438355145
+ 1.456e+11   
+       0.3251150179011032
+      0.03257737563420853
+       0.4006729027736295
+      0.02117176557917091
+     -0.07308904091700487
+       0.4016716576180642
+     0.001436506466881666
+      0.02121308889237537
+      0.03216788443097501
+       0.3256067358291423
+ 1.461e+11   
+       0.3228128202601531
+      0.03487856036156731
+       0.3976123648888069
+       0.0198199243796094
+      -0.0711143987370183
+       0.3986238547507942
+     0.002166526731355093
+       0.0198645737946666
+      0.03446319179695945
+       0.3233118722941138
+ 1.466e+11   
+       0.3205132865417465
+      0.03715853718293308
+       0.3945321203125517
+      0.01844381759277526
+     -0.06912506275741166
+       0.3955568486325347
+     0.002915515615776416
+      0.01849185867458391
+      0.03673728638791469
+       0.3210196621829045
+ 1.471e+11   
+       0.3182163117840929
+      0.03941725922585862
+       0.3914313214209065
+      0.01704316721260234
+     -0.06712056928069775
+        0.392469801996027
+     0.003683493635094749
+      0.01709465885606447
+      0.03899012184257233
+        0.318730001190758
+ 1.476e+11   
+       0.3159216695129555
+      0.04165494265440049
+       0.3883088640941934
+       0.0156175563791115
+     -0.06510015892828895
+        0.389361619432696
+     0.004470546406931914
+      0.01567255054226986
+      0.04122191480761341
+       0.3164426636742951
+ 1.481e+11   
+        0.313629003546993
+      0.04387208798523633
+       0.3851633668637985
+      0.01416641620317749
+     -0.06306274988983203
+       0.3862309263702029
+     0.005276832376623011
+       0.0142249576797915
+      0.04343316624810808
+       0.3141572944613486
+ 1.486e+11   
+       0.3113378197325982
+      0.04606950187673425
+       0.3819931493573366
+      0.01268901219240441
+     -0.06100691026680438
+       0.3830760473434088
+      0.00610259079940512
+      0.01275113842755575
+      0.04562468322952326
+       0.3118734005901548
+ 1.491e+11   
+       0.3090474776518228
+      0.04824831931081545
+       0.3787962100960141
+      0.01118443032056426
+     -0.05893082957874558
+        0.379894983613571
+     0.006948149954435004
+      0.01125017127341675
+      0.04779760109234612
+       0.3095903430207924
+ 1.496e+11   
+       0.3067571823528243
+      0.05041002607595627
+       0.3755702037043558
+     0.009651562789918997
+     -0.05683228951038818
+       0.3766853901961445
+     0.007813935560427013
+     0.009720940846715855
+      0.04995340592684298
+       0.3073073283681811
+ 1.501e+11   
+       0.3044659761589897
+      0.05255648144339077
+       0.3723124176120521
+     0.008089093547378468
+     -0.05470863400122647
+       0.3734445523770378
+     0.008700479356515706
+     0.008162123488179079
+      0.05209395724066302
+       0.3050234007132204
+ 1.506e+11   
+       0.3021727306208114
+      0.05468994091392203
+       0.3690197483404303
+     0.006495483624383676
+     -0.05255673879495786
+       0.3701693618121948
+     0.009608427804906439
+     0.006572172646335214
+      0.05422151069620493
+       0.3027374335551866
+ 1.511e+11   
+       0.2998761386820811
+      0.05681307889360072
+       0.3656886774887771
+     0.004868956384793583
+     -0.05037298059166246
+       0.3668562923253096
+      0.01053855086416863
+     0.004949304184365805
+      0.05633874077640666
+       0.3004481219774809
+ 1.516e+11   
+       0.2975747071412625
+      0.05892901113860273
+       0.3623152475526418
+     0.003207482776109245
+     -0.04815320596758538
+       0.3635013755372873
+      0.01149175077466638
+     0.003291481692864279
+         0.05844876321924
+       0.2981539751072541
+ 1.521e+11   
+       0.2952667494983888
+      0.06104131678764035
+       0.3588950377342361
+     0.001508766697140529
+     -0.04589270025876269
+       0.3601001764897548
+      0.01246907078602295
+     0.001596401920477237
+      0.06055515703896826
+       0.2958533089587373
+ 1.526e+11   
+       0.2929503792879468
+      0.06315405977781986
+       0.3554231399292971
+   -0.0002297693901593177
+     -0.04358615663257269
+       0.3566477694452876
+      0.01347170374931436
+   -0.0001385195504143861
+      0.06266198593097985
+       0.2935442397612773
+ 1.531e+11   
+       0.2906235040098065
+      0.06527180941547447
+       0.3518941351026845
+    -0.002010998457765741
+     -0.04122764560599058
+       0.3531387140829479
+      0.01450100048191244
+    -0.001916162235816135
+      0.06477381883062026
+       0.2912246778832345
+ 1.536e+11   
+       0.2882838197815381
+      0.06739965984670737
+       0.3483020703022622
+    -0.003838102350063848
+     -0.03881058530916747
+       0.3495670323353051
+      0.01555847780337434
+    -0.003739714124447436
+      0.06689574937217949
+        0.288892322475313
+ 1.541e+11   
+       0.2859288068486937
+      0.06954324814444615
+       0.3446404365902424
+     -0.00571458447516836
+     -0.03632771282911479
+       0.3459261861515633
+       0.0166458261243752
+    -0.005612684305173201
+      0.06903341396371444
+       0.2865446569698093
+ 1.546e+11   
+        0.283555726102866
+      0.07170877069810271
+       0.3409021482167625
+    -0.007644281535644793
+     -0.03377105701820282
+       0.3422090565112439
+      0.01776491645807754
+    -0.007538914635872512
+      0.07119300816481584
+       0.2841789455850667
+ 1.551e+11   
+       0.2811616167712501
+      0.07390299756074108
+       0.3370795233966928
+    -0.009631374060033508
+     -0.03113191319525286
+       0.3384079240523818
+      0.01891780670624009
+    -0.009522590215378945
+       0.0733813010221899
+       0.2817922309987781
+ 1.556e+11   
+       0.2787432954561315
+      0.07613328437510425
+       0.3331642671018615
+      -0.0116803954691217
+     -0.02840082022256708
+       0.3345144517294444
+      0.02010674705644362
+     -0.01156824839349899
+      0.07560564698382764
+       0.2793813333688731
+ 1.561e+11   
+       0.2762973567183633
+      0.07840758146421475
+       0.3291474563267017
+      -0.0137962393804148
+     -0.02556754049492895
+       0.3305196699597757
+      0.02133418430621251
+     -0.01368078602331681
+      0.07787399497887154
+       0.2769428508949994
+ 1.566e+11   
+       0.2738201754135204
+      0.08073443963721694
+        0.325019528339995
+     -0.01598416482492501
+     -0.02262104343653862
+       0.3264139647752117
+       0.0226027649148398
+     -0.01586546463080568
+      0.08019489421304889
+       0.2744731621299563
+ 1.571e+11   
+       0.2713079110055435
+      0.08312301222349854
+       0.3207702724903101
+     -0.01824979901652298
+     -0.01954949316294929
+       0.3221870695482226
+      0.02391533656031559
+     -0.01812791314301071
+      0.08257749619323802
+       0.2719684302652991
+ 1.576e+11   
+        0.268756514097741
+      0.08558305281181047
+       0.3163888261893473
+     -0.02059913728196043
+     -0.01634024102899562
+       0.3178280609209045
+      0.02527494796111898
+     -0.02047412778363665
+      0.08503155245832943
+       0.2694246096310113
+ 1.581e+11   
+       0.2661617354359382
+      0.08812490813332789
+       0.3118636757599608
+     -0.02303853972502116
+     -0.01297982384863253
+       0.3133253596253006
+      0.02668484670083638
+      -0.0229104687103709
+      0.08756740745497073
+       0.2668374546638202
+ 1.586e+11   
+       0.2635191376521627
+      0.09075950549267071
+       0.3071826628936847
+     -0.02557472416464033
+    -0.009453968641463988
+       0.3086667369445609
+      0.02814847477485367
+     -0.02544365293472121
+      0.09019598596312384
+       0.2642025316126735
+ 1.591e+11   
+       0.2608241100298934
+      0.09349833411656042
+       0.3023329975260356
+     -0.02821475485401327
+    -0.005747604823985045
+       0.3038393276250896
+      0.02966946155747835
+     -0.02808074303211286
+      0.09292877444086634
+       0.2615152332619974
+ 1.596e+11   
+       0.2580718865818435
+      0.09635341975939776
+       0.2973012779956541
+     -0.03096602645567546
+    -0.001844884830570075
+       0.2988296501105708
+      0.03125161387090191
+     -0.03082913111796012
+      0.09577779562809176
+       0.2587707969641633
+ 1.601e+11   
+       0.2552575677394257
+      0.09933729187795622
+       0.2920735194111059
+     -0.03383624271954975
+     0.002270785790477592
+        0.293623635023976
+      0.03289890282190431
+     -0.03369651753724281
+      0.09875557572194102
+       0.2559643262796937
+ 1.606e+11   
+       0.2523761459559606
+       0.1024629426678807
+       0.2866351912010349
+     -0.03683338928540433
+      0.00661670770535127
+        0.288206662878545
+      0.03461544705720283
+     -0.03669088369014706
+       0.1018751034161489
+       0.2530908165279595
+ 1.611e+11   
+       0.2494225355265175
+       0.1057437772401998
+       0.2809712648680947
+     -0.03996570001376851
+       0.0112108353997441
+       0.2825636120395882
+      0.03640549208193031
+     -0.03982045839733692
+       0.1051497800838111
+       0.2501451845505758
+ 1.616e+11   
+       0.2463916069197447
+       0.1091935542141568
+       0.2750662730015022
+     -0.04324161623539377
+      0.01607171187551069
+       0.2766789179974807
+      0.03827338527916457
+     -0.04309367719653186
+       0.1085933603791906
+       0.2471223029838555
+ 1.621e+11   
+       0.2432782259056105
+       0.1128263160093648
+       0.2689043806244398
+     -0.04666973830967425
+      0.02121838923351908
+        0.270536645030551
+      0.04022354627256206
+     -0.04651913395974241
+       0.1122198825430421
+       0.2440170393232296
+ 1.626e+11   
+       0.2400772977410305
+       0.1166563081445213
+       0.2624694699592501
+      -0.0502587688896831
+      0.02667033393266975
+       0.2641205713449789
+      0.04226043228260404
+     -0.05010552422993384
+       0.1160435877175416
+       0.2408243000428801
+ 1.631e+11   
+        0.236783816645916
+       0.1206978868878595
+       0.2557452396747651
+     -0.05401744731625322
+      0.03244731553545173
+       0.2574142887577266
+      0.04438849814847471
+     -0.05386157969912927
+       0.1200788276179336
+       0.2375390800025347
+ 1.636e+11   
+       0.2333929207609424
+       0.1249654146649843
+       0.2487153196416459
+     -0.05795447460391154
+      0.03856927779514865
+       0.2504013179536532
+      0.04661215071462643
+     -0.05779599328983109
+       0.1243399599655464
+       0.2341565173331672
+ 1.641e+11   
+       0.2298999527246877
+       0.1294731427113819
+       0.2413634021485848
+     -0.06207842854090166
+      0.04505619102117762
+       0.2430652402700418
+      0.04893569732772481
+     -0.06191733436280077
+       0.1288412311707535
+       0.2306719539397414
+ 1.646e+11   
+       0.2263005259410106
+       0.1342350805654396
+       0.2336733904268043
+     -0.06639766850921601
+      0.05192788477432739
+       0.2353898468591817
+      0.05136328824424635
+     -0.06623395365503758
+       0.1335966458615136
+       0.2270810016917451
+ 1.651e+11   
+       0.2225905965245112
+       0.1392648521351869
+       0.2256295651834992
+     -0.07092022973926143
+      0.05920386010412496
+       0.2273593059311228
+      0.05389885282411385
+     -0.07075387766205972
+       0.1386198229910617
+       0.2233796142900907
+ 1.656e+11   
+       0.2187665408127104
+       0.1445755382415619
+       0.2172167696516095
+     -0.07565370685096766
+      0.06690308075160156
+       0.2189583485849575
+      0.05654602947718286
+     -0.07548469231516437
+       0.1439238384283526
+       0.2195641646990382
+ 1.661e+11   
+       0.2148252382160709
+       0.1501795057465369
+       0.2084206134197708
+     -0.08060512670263548
+      0.07504374300358181
+       0.2101724734920101
+      0.05930808943987962
+     -0.08043341597267031
+       0.1495210541389345
+       0.2156315279151738
+ 1.666e+11   
+       0.2107641590411862
+       0.1560882236153827
+       0.1992276950067447
+       -0.085780810772418
+      0.08364302420995978
+       0.2009881703957077
+      0.06218785459171447
+     -0.08560636194820967
+       0.1554229343065749
+       0.2115791687089687
+ 1.671e+11   
+        0.206581456766843
+       0.1623120665452378
+       0.1896258427848068
+     -0.09118622753623168
+      0.09271681036281389
+        0.191393162029329
+      0.06518760967381572
+      -0.0910089910368295
+       0.1616398490275769
+       0.2074052338192321
+ 1.676e+11   
+       0.2022760640779012
+       0.1688601071127712
+       0.1796043734333161
+     -0.09682583558235783
+       0.1022794035925753
+       0.1813766636313695
+      0.06830900944609718
+     -0.09664575477632034
+       0.1681808665304862
+       0.2031086479065238
+ 1.681e+11   
+        0.197847791769299
+       0.1757398977560125
+       0.1691543666177779
+      -0.1027029185172569
+       0.1123432109614241
+       0.1709296587485412
+      0.07155298151655079
+      -0.1025199304940977
+       0.1750535352364376
+       0.1986892123782925
+ 1.686e+11   
+       0.1932974294224067
+       0.1829572443047033
+       0.1582689540358663
+      -0.1088194130661598
+       0.1229184165268319
+        0.160045189463175
+      0.07491962579117438
+      -0.1086334495386265
+       0.1822636573740972
+       0.1941477059891895
+ 1.691e+11   
+       0.1886268465320212
+       0.1905159732088796
+       0.1469436203616134
+      -0.1151757321557058
+       0.1340126393091131
+        0.148718658568668
+        0.078408111726541
+      -0.1149867204773377
+        0.189815056298502
+       0.1894859858961429
+ 1.696e+11   
+       0.1838390925281517
+       0.1984176950797587
+       0.1351765129481165
+      -0.1217705851776125
+       0.1456305805159595
+       0.1369481405442989
+      0.08201657481481614
+      -0.1215784494535495
+       0.1977093401276543
+        0.184707087613386
+ 1.701e+11   
+       0.1789384938972162
+       0.2066615676435977
+       0.1229687564352445
+       -0.128600798066021
+       0.1577736641485586
+       0.1247346974663184
+      0.08574201398694332
+      -0.1284054603273858
+       0.2059456647961095
+       0.1798153220740229
+ 1.706e+11   
+       0.1739307463694423
+        0.215244061707426
+       0.1103247676608383
+      -0.1356611362682707
+       0.1704396759208433
+       0.1120826952407423
+      0.08958019188013831
+      -0.1354625176717736
+       0.2145205001241239
+       0.1748163677662308
+ 1.711e+11   
+       0.1688229999103677
+       0.2241587342329468
+      0.09725256550879458
+      -0.1429441341357626
+        0.183622406251621
+       0.0990001147779636
+      0.09352554016829845
+      -0.1427421561399443
+       0.2234274029966485
+       0.1697173556843971
+ 1.716e+11   
+       0.1636239340454976
+       0.2333960130947862
+      0.08376406957204227
+      -0.1504399346970825
+       0.1973113039126295
+      0.08549885197077992
+      0.09757107239418138
+      -0.1502345201537824
+       0.2326568022272213
+       0.1645269446257165
+ 1.721e+11   
+       0.1583438208674555
+       0.2429429985439074
+      0.06987538078304679
+      -0.1581361441793318
+       0.2114911477077444
+      0.07159499961162222
+       0.1017083069571203
+      -0.1579272182655858
+       0.2421958001255307
+       0.1592553841839133
+ 1.726e+11   
+       0.1529945729382559
+        0.252783286784314
+      0.05560703650719667
+      -0.1660177059986202
+       0.2261417442869928
+      0.05730910372466741
+       0.1059272030825991
+      -0.1658051968960484
+       0.2520279961740421
+       0.1539145626545425
+ 1.731e+11   
+       0.1475897732184752
+       0.2628968213784618
+       0.0409842320351758
+      -0.1740667992253054
+       0.2412376608264082
+       0.0426663862294258
+       0.1102161127272271
+      -0.1738506384339708
+        0.262133338526727
+       0.1485180369853782
+ 1.736e+11   
+       0.1421446841434641
+       0.2732597783972692
+      0.02603699999455648
+      -0.1822627667210597
+       0.2567480017909686
+      0.02769692543363535
+       0.1145617514297654
+      -0.1820428888695333
+       0.2724880092424439
+       0.1430810418930087
+ 1.741e+11   
+       0.1366762330393517
+       0.2838444913002163
+      0.01080033896258193
+      -0.1905820782193309
+       0.2726362392984867
+      0.01243578561678274
+       0.1189491910975909
+      -0.1903584202018021
+       0.2830643492343429
+       0.1376204753389116
+ 1.746e+11   
+       0.1312029712404999
+       0.2946194214420479
+        0.384708695324211
+      -0.1989983335601047
+       0.2888601066769676
+       0.3836926019447007
+       0.1233618776044091
+      -0.1987708327924603
+       0.2938308288276035
+       0.1321548577256741
+ 1.751e+11   
+       0.1257450045485716
+       0.3055491798315202
+        0.403669841834463
+      -0.2074823110683096
+       0.3053715646085612
+       0.4026413230857376
+       0.1277816758545225
+      -0.2072509026062311
+       0.3047520695455452
+       0.1267042624507329
+ 1.756e+11   
+       0.1203238930696348
+       0.3165946052935094
+        0.422944776170639
+      -0.2160020656756673
+       0.3221168487464653
+       0.4219037053390645
+       0.1321889446345371
+      -0.2157666778731903
+       0.3157889222686312
+       0.1212902158491397
+ 1.761e+11   
+       0.1149625189876696
+       0.3277129034916225
+       0.4424658812257394
+      -0.2245230808115177
+       0.3390366068416347
+        0.441412132245275
+       0.1365626431161768
+      -0.2242836291149367
+       0.3268986062158394
+        0.115935565074635
+ 1.766e+11   
+       0.1096849214815646
+       0.3388578503440858
+       0.4621591268584033
+      -0.2330084773374134
+       0.3560661321989571
+       0.4610925671317997
+       0.1408804702953056
+      -0.2327648556959921
+       0.3380349122712653
+        0.110664313112703
+ 1.771e+11   
+       0.1045160987664043
+       0.3499800622112885
+       0.4819444098190936
+      -0.2414192818796928
+       0.3731356986927598
+       0.4808648898326462
+        0.145119037950568
+      -0.2411713511006673
+        0.349148473020927
+        0.105501420886135
+ 1.776e+11   
+      0.09948177813092482
+       0.3610273338536386
+       0.5017360064623833
+      -0.2497147558569176
+       0.3901710006078259
+       0.5006433452314353
+       0.1492540768970516
+      -0.2494623280196498
+       0.3601871004822241
+       0.1004725772951482
+ 1.781e+11   
+        0.094608155837939
+       0.3719450435764389
+       0.5214431387695488
+      -0.2578527853500697
+       0.4070936982618331
+       0.5203371038294995
+       0.1532606754059079
+      -0.2575956030947303
+        0.371096190919792
+      0.09560393901566268
+ 1.786e+11   
+      0.08992160983509472
+       0.3826766232214485
+       0.5409706511242107
+      -0.2657903307975186
+       0.4238220677497738
+       0.5398509313259416
+        0.157113547690028
+      -0.2655280398791495
+       0.3818191943761107
+      0.09092184294114894
+ 1.791e+11   
+      0.08544838936937343
+       0.3931640887756733
+       0.5602197918045616
+      -0.2734839344175084
+       0.4402717502936822
+       0.5590859605177154
+       0.1607873293457633
+      -0.2732160473038889
+       0.3922981446443415
+       0.0864524952710784
+ 1.796e+11   
+      0.08121428678578239
+       0.4033486253987736
+       0.5790890892984126
+       -0.280890282417284
+       0.4563565936697073
+       0.5779405546728872
+       0.1642568956344198
+      -0.2806161298171191
+       0.4024742434236444
+       0.0822216423944192
+ 1.801e+11   
+      0.07724429800168936
+       0.4131712186793915
+       0.5974753093210879
+      -0.2879668186425284
+        0.471989575119504
+        0.596311246852159
+       0.1674976975257669
+      -0.2876854845340327
+        0.412288490378747
+      0.07825422986481496
+ 1.806e+11   
+      0.07356227937317124
+       0.4225733219800786
+       0.6152744737981648
+      -0.2946724066416468
+       0.4870837921595417
+        0.614093734350322
+       0.1704861095619515
+      -0.2943826404083555
+        0.421682348836371
+      0.07457405689066632
+ 1.811e+11   
+      0.07019060992027804
+       0.4314975478789048
+       0.6323829179766943
+      -0.3009680385712108
+       0.5015535049078395
+       0.6311839012719749
+       0.1731997828853212
+      -0.3006681348894932
+       0.4305984349396596
+      0.07120343486161271
+ 1.816e+11   
+      0.06714986920295346
+       0.4398883700081062
+       0.6486983560493695
+       -0.306817592536579
+       0.5153152110928354
+       0.6474788348368519
+       0.1756179962591574
+      -0.3065052251459107
+       0.4389812162852568
+      0.06816285951369409
+ 1.821e+11   
+      0.06445854264449692
+       0.4476928200437156
+       0.6641209188346053
+      -0.3121886456894871
+       0.5282887329212708
+       0.6628777916169742
+       0.1777219976434219
+      -0.3118606342426106
+       0.4467777043901607
+      0.06547070744932847
+ 1.826e+11   
+      0.06213276798816583
+        0.454861163181142
+       0.6785541184927912
+       -0.317053359903115
+       0.5403982935690405
+       0.6772830573833561
+       0.1794953288974033
+      -0.3167053383913743
+        0.453938123722644
+      0.06314296898280221
+ 1.831e+11   
+      0.06018613918003719
+       0.4613475340220977
+       0.6919056839385798
+      -0.3213894717515167
+       0.5515735602733334
+       0.6906006268700323
+       0.1809241264554627
+       -0.321015410517632
+       0.4604165383535642
+      0.06119303086333776
+ 1.836e+11   
+      0.05862958780257405
+       0.4671105131395281
+       0.7040881950709523
+      -0.3251814406787524
+        0.561750630778234
+       0.7027406053838521
+       0.1819973912475159
+      -0.3247729490410623
+       0.4661714152896828
+      0.05963152462514823
+ 1.841e+11   
+      0.05747136783202347
+       0.4721136221998703
+       0.7150194226183494
+      -0.3284218393783794
+       0.5708729398805926
+       0.7136172013803057
+       0.1827072213443538
+      -0.3279671396987835
+       0.4711661008830941
+      0.05846625948307386
+ 1.846e+11   
+      0.05671717711656379
+        0.476325711619362
+       0.7246222532248566
+      -0.3311131029527965
+       0.5788920620432227
+       0.7231481421591418
+       0.1830489997664942
+      -0.3305955207289503
+       0.4753691830729717
+      0.05770226303227776
+ 1.851e+11   
+      0.05637045610188408
+        0.479721208250193
+       0.7328240538213726
+      -0.3332697589189496
+       0.5857683818925815
+       0.7312533311911198
+       0.1830215248657782
+      -0.3326655366837881
+       0.4787547082203057
+      0.05734195764343029
+ 1.856e+11   
+        0.056432897997235
+       0.4822801809896351
+       0.7395553402005555
+      -0.3349211282657854
+        0.591471590283317
+       0.7378526836865082
+       0.1826270544529374
+      -0.3341964315287409
+       0.4813022216692611
+      0.05738550024596474
+ 1.861e+11   
+      0.05690513486585435
+       0.4839881736228863
+       0.7447477875363302
+      -0.3361138512463424
+       0.5959809230840161
+       0.7428636976885338
+       0.1818711888292492
+      -0.3352213097517768
+       0.4829966258469078
+      0.05783128856327385
+ 1.866e+11   
+       0.0577872618948985
+       0.4848357730662702
+       0.7483323632694734
+      -0.3369113214001632
+       0.5992849549743928
+       0.7462016025006308
+       0.1807623971000121
+      -0.3357883655172695
+       0.4838279689156942
+      0.05867652258873515
+ 1.871e+11   
+      0.05907782377875963
+       0.4848180419338083
+       0.7502408998000258
+       -0.337380157254947
+       0.6013805224945244
+       0.7477920696926017
+       0.1793107065289495
+      -0.3359576655844387
+       0.4837917044323328
+      0.05991730985923129
+ 1.876e+11   
+      0.06076700470215951
+       0.4839346517962158
+        0.750421937759951
+      -0.3375366019451029
+       0.6022699707659075
+       0.7476245498250809
+       0.1775245744284384
+      -0.3357826859981478
+       0.4828911809710763
+      0.06154661640632943
+ 1.881e+11   
+      0.06281499724551955
+       0.4821937981734526
+       0.7488992631330399
+       -0.337204065406535
+       0.6019561335644007
+       0.7458983070327119
+       0.1754049797070677
+      -0.3352506699929524
+       0.4811462388320125
+      0.06354563853982004
+ 1.886e+11   
+      0.06511367602343349
+       0.4796265690988477
+       0.7459181667539834
+      -0.3358041353309642
+       0.6004387575688723
+       0.7432440765575281
+       0.1729403039048874
+      -0.3341471612479545
+       0.4786094542824076
+      0.06586166976334792
+ 1.891e+11   
+      0.06749029397668856
+       0.4763102114457934
+       0.7421287714036928
+      -0.3324868393634531
+       0.5977270883767836
+       0.7406085559974753
+       0.1701188510304887
+      -0.3319085291959828
+       0.4753683069756685
+       0.0683791955846059
+ 1.896e+11   
+      0.06984765840209803
+       0.4723556837934141
+        0.738379945710989
+      -0.3270579746273002
+       0.5938733780414773
+       0.7383110743409713
+       0.1669679835797603
+      -0.3278491159320272
+       0.4714956709551976
+        0.070945028783111
+ 1.901e+11   
+      0.07227261626540873
+       0.4678260925940658
+       0.7348381587573669
+      -0.3204456954859298
+       0.5889775699645683
+       0.7355350137781762
+       0.1635654582784477
+       -0.321965502858236
+       0.4670031393515964
+       0.0734976368074348
+ 1.906e+11   
+      0.07489727870169476
+       0.4627040117860521
+        0.730711481554597
+      -0.3136659989009719
+       0.5831397232379799
+       0.7313495351112858
+       0.1599887125437078
+      -0.3151322523636866
+       0.4618758108314206
+      0.07612566007399102
+ 1.911e+11   
+      0.07776685899375911
+       0.4569649142388027
+       0.7252025550541055
+      -0.3071081622000255
+       0.5764303088597427
+       0.7254415775527914
+       0.1562781787932495
+      -0.3081926671355447
+       0.4561194309433879
+      0.07893625773646208
+ 1.916e+11   
+      0.08085722181449277
+       0.4506254195904073
+        0.718071136173675
+      -0.3007564613914362
+       0.5689034582133604
+       0.7179146083050102
+        0.152449679659682
+      -0.3014577409848668
+       0.4497676115227818
+      0.08195959647918541
+ 1.921e+11   
+      0.08412270049392906
+       0.4437322913572803
+       0.7094344313811892
+      -0.2944994673576071
+       0.5606145650717407
+       0.7089854105965538
+       0.1485148936167422
+      -0.2949124246152969
+       0.4428703129121678
+      0.08516973077693057
+ 1.926e+11   
+      0.08751820322268605
+         0.43634319575539
+       0.6995046388814626
+      -0.2882481611053435
+       0.5516255916328879
+       0.6988611301474179
+       0.1444889485172417
+      -0.2884641482217009
+       0.4354836996416984
+      0.08852366970973539
+ 1.931e+11   
+      0.09100447033157665
+       0.4285175716422744
+       0.6884827685554962
+      -0.2819533817916418
+       0.5420039084485215
+       0.6877157728661791
+       0.1403904309645101
+      -0.2820387113472165
+       0.4276652462252082
+      0.09197934032201874
+ 1.936e+11   
+      0.09454795648705507
+       0.4203138614737934
+       0.6765384337516676
+      -0.2755966733571791
+       0.5318199851080585
+       0.6756952642473462
+       0.1362397442983283
+      -0.2755954127051713
+       0.4194719525080629
+       0.0955000639912859
+ 1.941e+11   
+      0.09811976985154286
+       0.4117889144564678
+       0.6638146083539223
+      -0.2691791632459189
+       0.5211454781266923
+       0.6629260559534914
+       0.1320577222890791
+      -0.2691197841453786
+       0.4109597410811887
+      0.09905455210136782
+ 1.946e+11   
+       0.1016947820374094
+       0.4029978826740787
+       0.6504354819915728
+      -0.2627134237524558
+       0.5100518295967054
+       0.6495215904529801
+       0.1278647207843907
+      -0.2626142302224886
+       0.4021831846149307
+       0.1026160257310941
+ 1.951e+11   
+       0.1052510379343503
+       0.3939941420485721
+       0.6365123754704144
+      -0.2562181930946597
+       0.4986092312342542
+        0.635586326792109
+       0.1236800570833823
+      -0.2560909977738086
+       0.3931952886570556
+       0.1061614300726326
+ 1.956e+11   
+       0.1087693864592734
+       0.3848291575726855
+       0.6221474489345759
+      -0.2497150664832242
+       0.4868858319215758
+       0.6212180339315787
+       0.1195216673390707
+      -0.2495675405333319
+        0.384047268496547
+       0.1096708847847616
+ 1.961e+11   
+       0.1122332439356582
+       0.3755523076730006
+       0.6074358372325658
+      -0.2432264338958721
+       0.4749471164563376
+         0.60650900372209
+       0.1154058999298163
+      -0.2430635868787941
+       0.3747883211640395
+       0.1131273183438894
+ 1.966e+11   
+       0.1156284279388016
+       0.3662106950704602
+       0.5924668021822895
+      -0.2367741938490698
+       0.4628554157524516
+       0.5915466279776328
+       0.1113473978872814
+      -0.2365993086284249
+       0.3654654060759916
+       0.1165162165874443
+ 1.971e+11   
+       0.1189430233582889
+       0.3568489653480766
+       0.5773243056207423
+      -0.2303789557015808
+       0.4506695260186476
+       0.5764136166534617
+        0.107359043661416
+      -0.2301941857378045
+       0.3561230463376308
+       0.1198254338396019
+ 1.976e+11   
+       0.1221672587925286
+       0.3475091465851509
+       0.5620872557386798
+      -0.2240595570529959
+       0.4384444228278701
+       0.5611880243709504
+       0.1034519502508258
+      -0.2238663136689749
+        0.346803158596932
+       0.1230450341096758
+ 1.981e+11   
+       0.1252933816565871
+       0.3382305173818803
+        0.546829579332222
+      -0.2178327903805561
+       0.4262310597987429
+       0.5459431850507359
+      0.09963548832437823
+      -0.2176319978450055
+       0.3375449156331196
+       0.1261671435648449
+ 1.986e+11   
+       0.1283155266159481
+       0.3290495065100102
+       0.5316202109333621
+      -0.2117132726457524
+       0.4140762432126849
+       0.5307476136877309
+      0.09591734189464389
+      -0.2115055387873188
+        0.328384643121154
+       0.1291858043002233
+ 1.991e+11   
+       0.1312295756732706
+       0.3199996247918129
+       0.5165230524610668
+      -0.2057134149256301
+       0.4020225745017968
+       0.5156649097165189
+      0.09230358669538129
+      -0.2054991468314934
+       0.3193557501405462
+       0.1320968248516607
+ 1.996e+11   
+       0.1340330104004671
+       0.3111114281639772
+        0.501596934485903
+      -0.1998434630898353
+       0.3901084527676456
+       0.5007536814573745
+      0.08879878634370904
+      -0.1996229464453394
+       0.3104886917796377
+       0.1348976261373092
+ 2.001e+11   
+       0.1367247580155264
+       0.3024125098938587
+       0.4868955964994907
+      -0.1941115891156419
+       0.3783681296202555
+       0.4860675019449713
+      0.08540610197706483
+      -0.1938850430147005
+        0.301810961440342
+       0.1375870833874911
+ 2.006e+11   
+       0.1393050336106126
+       0.2939275193601564
+       0.4724676951928142
+      -0.1885240180697419
+       0.3668318087920545
+       0.4716549007555264
+      0.08212741151855228
+      -0.1882916329597795
+       0.2933471100331326
+       0.1401653656423342
+ 2.011e+11   
+       0.1417751810653841
+       0.2856782045440288
+       0.4583568445889867
+        -0.18308517937963
+       0.3555257832344152
+       0.4575593929229078
+       0.0789634351255257
+      -0.1828471431900374
+        0.285118789067995
+       0.1426337748812398
+ 2.016e+11   
+       0.1441375151658625
+       0.2776834753032726
+        0.444601688708045
+      -0.1777978735118004
+       0.3444726027551882
+       0.4438195438661447
+      0.07591386375401625
+      -0.1775543893511156
+       0.2771448146225967
+       0.1449945869964347
+ 2.021e+11   
+       0.1463951672840138
+       0.2699594845547307
+       0.4312360055177892
+      -0.1726634469985117
+       0.3336912656946277
+       0.4304690679483944
+      0.07297748814067735
+      -0.1724147447323327
+       0.2694412492520965
+       0.1472508967609061
+ 2.026e+11   
+         0.14855193671653
+       0.2625197246248521
+       0.4182888397922468
+      -0.1676819701588891
+       0.3231974286455291
+       0.4175369575451344
+      0.07015232586764839
+       -0.167428313478923
+        0.262021499058299
+       0.1494064687508241
+ 2.031e+11   
+       0.1506121494738253
+       0.2553751362101416
+       0.4057846618719911
+       -0.162852412989739
+       0.3130036287803045
+       0.4050476391218228
+      0.06743574453217586
+      -0.1625941031192412
+       0.2548964233310552
+        0.151465595918777
+ 2.036e+11   
+       0.1525805259807546
+       0.2485342275977923
+       0.3937435490207415
+      -0.1581728156409123
+        0.303119513931399
+       0.3930211526820535
+      0.06482457938729759
+      -0.1579101925092145
+       0.2480744543913626
+       0.1534329672134727
+ 2.041e+11   
+       0.1544620588188021
+       0.2420032020134248
+       0.3821813859822552
+      -0.1536404506897758
+       0.2935520761633365
+       0.3814733509627228
+      0.06231524414787252
+      -0.1533738921952373
+       0.2415617254889596
+       0.1553135453294105
+ 2.046e+11   
+       0.1562619013196769
+       0.2357860911777734
+       0.3711100813857562
+      -0.1492519751182418
+       0.2843058851582402
+       0.3704161148669866
+      0.05990383396321378
+      -0.1489818949509477
+       0.2353622048267897
+       0.1571124553635562
+ 2.051e+11   
+       0.1579852675218041
+       0.2298848933589509
+       0.3605377967759201
+      -0.1450035704919223
+       0.2753833182991182
+       0.3598575818003041
+      0.05758621984030825
+      -0.1447304148827939
+       0.2294778339929165
+       0.1588348848668249
+ 2.056e+11   
+       0.1596373437303247
+       0.2242997143975336
+       0.3504691852216938
+      -0.1408910703553178
+       0.2667847848662796
+        0.349802383785609
+      0.05535813405733679
+      -0.1406153140427162
+       0.2239086692744625
+       0.1604859955139926
+ 2.061e+11   
+       0.1612232116815771
+        0.219028910355551
+       0.3409056366646479
+      -0.1369100742976393
+       0.2585089422550722
+       0.3402518924616591
+      0.05321524633472181
+      -0.1366322159465242
+       0.2186530245040503
+       0.1620708463805697
+ 2.066e+11   
+       0.1627477831061821
+       0.2140692305966978
+       0.3318455273873496
+      -0.1330560485167316
+       0.2505529025730249
+       0.3312044683042379
+       0.0511532307297447
+      -0.1327766057828751
+       0.2137076142477781
+       0.1635943286119371
+ 2.071e+11   
+       0.1642157453111028
+       0.2094159602445108
+     0.002915372897803001
+      -0.1293244130191617
+        0.242912428378907
+     0.004731837879202654
+       0.0491678233908765
+      -0.1290439174175414
+       0.2090676962845943
+       0.1650611110987049
+ 2.076e+11   
+       0.1656315172593607
+       0.2050630610887929
+     0.009609486448374468
+      -0.1257106158478176
+       0.2355821166845755
+      0.01142693702998166
+      0.04725487145040307
+      -0.1254296075574454
+       0.2047272124520275
+       0.1664755966326054
+ 2.081e+11   
+       0.1669992155147163
+       0.2010033101199486
+      0.01611358410411182
+      -0.1222101949295074
+       0.2285555706534584
+      0.01793002488230529
+      0.04541037345020949
+       -0.121929217644669
+       0.2006789270435757
+       0.1678418879072986
+ 2.086e+11   
+       0.1683226293353822
+       0.1972284349681859
+      0.02243092672798748
+      -0.1188188282890565
+       0.2218255586988014
+      0.02424446414345681
+      0.04363051178720599
+      -0.1185384242080847
+       0.1969145620411245
+       0.1691637626463853
+ 2.091e+11   
+       0.1696052041429433
+       0.1937292456114255
+      0.02856489460085312
+      -0.1155323734884418
+       0.2153841609129489
+      0.03037374415177588
+      0.04191167773403868
+      -0.1152530785147871
+       0.1934249285535082
+       0.1704446570840192
+ 2.096e+11   
+       0.1708500325574632
+       0.1904957617944815
+      0.03451892848080322
+      -0.1123468972246244
+       0.2092229029489602
+      0.03632142062083937
+      0.04025048963951155
+      -0.1120692364406893
+       0.1902000539110707
+       0.1716876569889056
+ 2.101e+11   
+       0.1720598521742008
+       0.1875173356737176
+      0.04029648230047429
+      -0.1092586960628527
+       0.2033328776311355
+       0.0420910670680857
+      0.03864380494395343
+      -0.1089831795243664
+       0.1872293039382465
+       0.1728954954076588
+ 2.106e+11   
+       0.1732370492587948
+       0.1847827692680424
+      0.04590098627519047
+      -0.1062643092980984
+        0.197704854694938
+      0.04768623671007721
+      0.03708872665945993
+      -0.1059914281855309
+       0.1845014999927544
+       0.1740705563052723
+ 2.111e+11   
+       0.1743836675533306
+        0.182280426359238
+      0.05133581920474563
+      -0.1033605249304374
+       0.1923293791529852
+      0.05311043361474403
+      0.03558260496633182
+      -0.1030907480838584
+       0.1820050304220482
+       0.1752148832964455
+ 2.116e+11   
+       0.1755014214129277
+       0.1799983385437531
+      0.05660428878522972
+      -0.1005443797146631
+       0.1871968588554825
+      0.05836709193289256
+      0.03412303456653119
+      -0.1002781505695218
+       0.1797279561466085
+       0.1763301926889834
+ 2.121e+11   
+       0.1765917125289157
+       0.1779243051942511
+      0.06170961879917542
+     -0.09781315420420017
+       0.1822976418640807
+      0.06345956208165503
+       0.0327078484152083
+     -0.09755088813755793
+       0.1776581101354903
+       0.1774178900971822
+ 2.126e+11   
+        0.177655649538345
+       0.1760459871432735
+      0.06665494211808269
+     -0.09516436365775985
+       0.1776220842905953
+      0.06839110281701755
+      0.03133510842369612
+     -0.09490644574751965
+       0.1757831905932672
+       0.1784790899268855
+ 2.131e+11   
+       0.1786940698683274
+       0.1743509939532673
+      0.07144329852685348
+     -0.09259574561731609
+       0.1731606092691263
+       0.0731648782067927
+       0.0300030936938076
+     -0.09234252881090796
+       0.1740908477288604
+       0.1795146370828028
+ 2.136e+11   
+       0.1797075632160735
+       0.1728269646870631
+      0.07607763646156736
+     -0.09010524490045323
+       0.1689037577345797
+       0.0777839585962475
+      0.02871028680515493
+      -0.0898570485842077
+       0.1725687640261364
+        0.180525130301078
+ 2.141e+11   
+       0.1806964961199332
+       0.1714616421406434
+      0.08056081783718602
+     -0.08769099668136494
+       0.1648422316743983
+       0.0822513247428415
+      0.02745535863606451
+     -0.08744810563734309
+        0.171204727983389
+       0.1815109465645842
+ 2.146e+11   
+       0.1816610371319513
+       0.1702429405455475
+       0.0848956252279687
+      -0.0853513082646335
+       0.1609669305058255
+      0.08656987438184915
+      0.02623715215547499
+     -0.08511397199797394
+       0.1699867013336638
+        0.182472266113528
+ 2.151e+11   
+       0.1826011821574034
+       0.1691590067911362
+      0.08908477074848702
+     -0.08308464008603626
+       0.1572689812098219
+      0.09074243056909913
+      0.02505466557928701
+     -0.08285307250288407
+       0.1689028798003631
+       0.1834090976189875
+ 2.156e+11   
+       0.1835167795807255
+       0.1681982752573573
+      0.09313090606571554
+     -0.08088958640635775
+       0.1537397628264764
+       0.0947717512290288
+      0.02390703524057528
+     -0.08066396582001914
+         0.16794174748227
+       0.1843213031406919
+ 2.161e+11   
+        0.184407554849183
+       0.1673495163858487
+      0.09703663305137364
+      -0.0787648560985406
+       0.1503709258867334
+      0.09866053941446866
+      0.02279351847988673
+     -0.07854532553974407
+       0.1670921249988735
+       0.1852086225423576
+ 2.166e+11   
+       0.1852731342353796
+        0.166601879151506
+       0.1008045146578889
+     -0.07670925386629038
+       0.1471544073226475
+       0.1024114538583599
+      0.02171347681992632
+     -0.07649592167214292
+        0.166343211560611
+       0.1860706970873956
+ 2.171e+11   
+       0.1861130675464733
+       0.1659449276274044
+       0.1044370856701163
+     -0.07472166217407815
+       0.1440824413641307
+       0.1060271194660702
+      0.02066635964894218
+     -0.07451460282950118
+       0.1656846211588975
+       0.1869070919845122
+ 2.176e+11   
+       0.1869268495917632
+       0.1653686718634422
+       0.1079368630482739
+     -0.07280102411466864
+       0.1411475668951022
+       0.1095101374600468
+      0.01965168859925272
+     -0.07260027931974618
+       0.1651064130978251
+       0.1877173176963404
+ 2.181e+11   
+       0.1877139402606613
+       0.1648635933228254
+       0.1113063556348691
+     -0.07094632739120361
+       0.1383426317067423
+       0.1128630949456919
+      0.01866904277210353
+      -0.0707519073278479
+       0.1645991171127196
+       0.1885008498644451
+ 2.186e+11   
+       0.1884737831000836
+       0.1644206651408575
+       0.1145480730500295
+     -0.06915658954644967
+       0.1356607940507002
+       0.1160885737188922
+      0.01771804492737834
+     -0.06896847431811172
+       0.1641537533406738
+       0.1892571477408828
+ 2.191e+11   
+        0.189205822313736
+       0.1640313674871168
+       0.1176645336454902
+     -0.06743084453216924
+       0.1330955218611523
+        0.119189158181374
+      0.01679834872688293
+     -0.06724898575094086
+       0.1637618474244475
+       0.1899856710498366
+ 2.196e+11   
+       0.1899095181358483
+       0.1636876983253525
+       0.1206582714277139
+     -0.06576813067658503
+       0.1306405899816713
+       0.1221674422703506
+      0.01590962709295786
+     -0.06559245317280796
+       0.1634154410440053
+       0.1906858952326487
+ 2.201e+11   
+        0.190584360558455
+       0.1633821798751776
+       0.1235318418956984
+     -0.06416748007729632
+       0.1282900757014813
+       0.1250260353439372
+      0.01505156172004361
+     -0.06399788370787983
+       0.1631070981794497
+       0.1913573250561202
+ 2.206e+11   
+       0.1912298814147812
+       0.1631078610862438
+       0.1262878267690361
+     -0.06262790942075878
+       0.1260383528757656
+       0.1277675669939713
+      0.01422383375549716
+     -0.06246427095352944
+       0.1628299074154088
+       0.1919995065870848
+ 2.211e+11   
+        0.191845664841412
+       0.1628583164390171
+       0.1289288376071838
+     -0.06114841220708039
+       0.1238800848765287
+       0.1303946907833277
+      0.01342611564732044
+     -0.06099058725980577
+        0.162577480600199
+       0.1926120375563788
+ 2.216e+11   
+       0.1924313561592432
+       0.1626276413869369
+       0.1314575183421399
+     -0.05972795234027714
+       0.1218102165941834
+       0.1329100869261815
+        0.012658064140439
+     -0.05957577735436315
+       0.1623439481734998
+       0.1931945761523958
+ 2.221e+11   
+       0.1929866692276505
+        0.162410444752748
+       0.1338765467640002
+     -0.05836545902887898
+       0.1198239656854033
+       0.1353164639470875
+      0.01191931438952319
+     -0.05821875325921815
+       0.1621239514741733
+       0.1937468482988401
+ 2.226e+11   
+       0.1935113923382567
+       0.1622018383874026
+       0.1361886350127354
+     -0.05705982292965814
+        0.117916813240142
+       0.1376165593687769
+      0.01120947514507582
+     -0.05691839043355575
+       0.1619126323352842
+       0.1942686534830002
+ 2.231e+11   
+       0.1940053927241853
+       0.1619974243934142
+       0.1383965291402207
+     -0.05580989345787163
+       0.1160844940196885
+       0.1398131394894317
+      0.01052812496024835
+     -0.05567352506747848
+       0.1617056202668197
+       0.1947598692103459
+ 2.236e+11   
+       0.1944686197680988
+       0.1617932802061805
+       0.1405030078145769
+     -0.05461447718051236
+       0.1143229863985089
+        0.141908998318382
+     0.009874809358625858
+      -0.0544829524447059
+       0.1614990175180958
+       0.1952204541685433
+ 2.241e+11   
+       0.1949011069977409
+        0.161585941816743
+       0.1425108802443895
+     -0.05347233720438641
+       0.1126285021250823
+       0.1439069557449005
+     0.009249038897669161
+     -0.05334542628748871
+       0.1612893823018053
+       0.1956504501892967
+ 2.246e+11   
+       0.1953029729614205
+       0.1613723854080901
+       0.1444229834038968
+     -0.05238219346801226
+       0.1109974760010767
+       0.1458098550184246
+     0.008650288058646288
+     -0.05225965899419151
+       0.1610737104501896
+       0.1960499831000847
+ 2.251e+11   
+        0.195674421077995
+       0.1611500076645652
+       0.1462421786418753
+     -0.05134272384522551
+       0.1094265555638362
+        0.147620559620422
+     0.008077994891296698
+     -0.05122432267882845
+       0.1608494157613345
+       0.1964192625599335
+ 2.256e+11   
+        0.196015738556755
+        0.160916605000516
+       0.1479713477571241
+     -0.05035256596862907
+       0.1079125908442415
+       0.1493419496084386
+      0.00753156134029639
+     -0.05023805092201241
+       0.1606143092800903
+        0.196758580974088
+ 2.261e+11   
+       0.1963272944821624
+       0.1606703519401671
+        0.149613388622353
+     -0.04941031968249173
+       0.1064526242604562
+       0.1509769175119429
+     0.007010354180362643
+     -0.04929944114424507
+       0.1603665777440552
+        0.197068311582081
+ 2.266e+11   
+       0.1966095371570937
+       0.1604097788661188
+       0.1511712104360748
+     -0.04851455003712928
+       0.1050438806977316
+       0.1525283638576078
+     0.006513706487647479
+     -0.04840705751476342
+       0.1601047614104279
+       0.1973489058121793
+ 2.271e+11   
+       0.1968629907959204
+       0.1601337493388747
+       0.1526477286791331
+     -0.04766379074009251
+       0.1036837578153274
+        0.153999192398842
+     0.006040919576602223
+     -0.04755943431243222
+       0.1598277314646516
+       0.1976008899930223
+ 2.276e+11   
+       0.1970882516558497
+       0.1598414371747779
+       0.1540458598488378
+      -0.0468565479832893
+       0.1023698166135307
+       0.1553923051208607
+     0.005591265333766926
+     -0.04675507965890608
+       0.1595346671967318
+       0.1978248615102238
+ 2.281e+11   
+       0.1972859836914203
+       0.1595323034545978
+       0.1553685160394439
+     -0.04609130456963891
+       0.1010997722866582
+        0.156710597088637
+     0.005163988882703764
+     -0.04599247954860611
+       0.1592250331160925
+       0.1980214844921951
+ 2.286e+11   
+       0.1974569138130333
+       0.1592060736201001
+       0.1566185994332671
+     -0.04536652426750432
+      0.09987148538174304
+        0.157956951200603
+     0.004758311517528269
+     -0.04527010210475903
+       0.1588985561609139
+       0.1981914851054709
+ 2.291e+11   
+       0.1976018268260897
+        0.158862714801227
+       0.1577989967618471
+     -0.04468065632618784
+       0.0986829532772437
+       0.1591342329064252
+     0.004373433846047251
+     -0.04458640199557212
+       0.1585552031433297
+       0.1983356465354396
+ 2.296e+11   
+       0.1977215601226743
+       0.1585024135021396
+       0.1589125737917096
+     -0.04403214009088383
+      0.09753230199147124
+       0.1602452849423341
+     0.004008539087355733
+     -0.04393982494975767
+       0.1581951585575135
+       0.1984548037238404
+ 2.301e+11   
+       0.1978169981929911
+       0.1581255537605097
+       0.1599621698842703
+     -0.04341940966068036
+      0.09641777832647073
+       0.1612929221326578
+     0.003662796472716172
+     -0.04332881231568365
+       0.1578188028638885
+       0.1985498379295628
+ 2.306e+11   
+       0.1978890670188598
+       0.1577326958809867
+       0.1609505926744474
+     -0.04284089853841141
+      0.09533774234970081
+       0.1622799263013711
+     0.003335364702656613
+     -0.04275180561360965
+       0.1574266913493468
+       0.1986216711745293
+ 2.311e+11   
+       0.1979387284066579
+       0.1573245558309504
+         0.16188061290768
+     -0.04229504422625686
+       0.0942906602130572
+       0.1632090413326988
+     0.003025395417352497
+     -0.04220725103544931
+       0.1570195336505859
+       0.1986712606314177
+ 2.316e+11   
+       0.1979669743122731
+       0.1569019853743984
+       0.1627549594703062
+     -0.04178029272603798
+      0.09327509730639187
+       0.1640829684151867
+     0.002732036641515207
+     -0.04169360385154146
+       0.1565981740155032
+       0.1986995930052698
+ 2.321e+11   
+       0.1979748212057183
+       0.1564659530082291
+       0.1635763146436155
+     -0.04129510290796383
+       0.0922897117407364
+       0.1649043614991243
+     0.002454436169054954
+     -0.04120933268859953
+       0.1561635723660722
+       0.1987076789560908
+ 2.326e+11   
+       0.1979633045184247
+       0.1560175257542283
+       0.1643473096075559
+     -0.04083795071628384
+      0.09133324815487615
+       0.1656758229929517
+     0.002191744856807442
+     -0.04075292364770348
+       0.1557167862152472
+        0.198696547604975
+ 2.331e+11   
+       0.1979334732115823
+       0.1555578518497946
+       0.1650705202158786
+     -0.04040733318474164
+      0.09040453183766832
+       0.1663998997201853
+     0.001943119800450826
+     -0.04032288423554198
+       0.1552589534802468
+       0.1986672411616541
+ 2.336e+11   
+       0.1978863844995496
+       0.1550881443709027
+       0.1657484630605646
+     -0.04000177223893443
+       0.0895024631574983
+       0.1670790791545397
+      0.00170772736947551
+     -0.03991774708628514
+       0.1547912762250855
+       0.1986208097070288
+ 2.341e+11   
+       0.1978230987580389
+       0.1546096658118624
+       0.1663835918397309
+      -0.0396198182666479
+      0.08862601228958793
+       0.1677157859473316
+     0.001484746081600152
+     -0.03953607345539958
+       0.1543150053563753
+       0.1985583061600251
+ 2.346e+11   
+       0.1977446746428227
+       0.1541237136382553
+       0.1669782940397384
+     -0.03926005344097771
+      0.08777421423128627
+       0.1683123787578685
+     0.001273369300389644
+      -0.0391764564703932
+       0.1538314262882758
+       0.1984807814541016
+ 2.351e+11   
+       0.1976521644408304
+       0.1536316068218646
+       0.1675348879390954
+     -0.03892109478447466
+      0.08694616409519355
+       0.1688711473944665
+     0.001072807743000091
+     -0.03883752412684553
+       0.1533418455850201
+       0.1983892799449662
+ 2.356e+11   
+       0.1975466096719304
+       0.1531346733595512
+       0.1680556199388147
+     -0.03860159696575693
+      0.08614101266971172
+       0.1693943102707941
+    0.0008822917879177388
+     -0.03851794202131081
+       0.1528475785825607
+       0.1982848350674599
+ 2.361e+11   
+       0.1974290369562718
+        0.152634238771728
+       0.1685426622212045
+     -0.03830025482296672
+      0.08535796223660136
+       0.1698840121797268
+    0.0007010735753211711
+     -0.03821641581549417
+       0.1523499379847482
+       0.1981684652562312
+ 2.366e+11   
+       0.1973004541589387
+       0.1521316155705066
+       0.1689981107366921
+     -0.03801580561112703
+      0.08459626263512227
+       0.1703423223844331
+    0.0005284288952083832
+     -0.03793169342881871
+       0.1518502234237983
+        0.198041170141668
+ 2.371e+11   
+       0.1971618468207075
+       0.1516280936824642
+       0.1694239835160416
+     -0.03774703097289659
+      0.08385520756245467
+       0.1707712330243229
+    0.0003636588607695025
+     -0.03766256695886844
+       0.1513497119698585
+       0.1979039270296912
+ 2.376e+11   
+       0.1970141748809716
+       0.1511249318065458
+       0.1698222193034059
+     -0.03749275863438185
+      0.08313413110030757
+       0.1711726578315386
+     0.000206091366590197
+     -0.03740787433134356
+       0.1508496495700053
+       0.1977576876712644
+ 2.381e+11   
+       0.1968583696964279
+       0.1506233496836315
+       0.1701946765038956
+     -0.03725186382966183
+      0.08243240445781994
+       0.1715484311519608
+    5.508233316411622e-05
+     -0.03716650068314663
+       0.1503512433931079
+       0.1976033753250624
+ 2.386e+11   
+       0.1966953313567905
+       0.1501245212508531
+       0.1705431324378138
+     -0.03702327045938746
+      0.08174943292117105
+       0.1719003072631973
+   -8.998325908533833e-05
+     -0.03693737948387908
+       0.1498556550535759
+       0.1974418821144276
+ 2.391e+11   
+       0.1965259262967441
+       0.1496295686507731
+        0.170869282892336
+      -0.0368059519903642
+      0.08108465300058425
+       0.1722299599806913
+   -0.0002296905415689273
+     -0.03671949340256415
+        0.149363994684102
+       0.1972740666777214
+ 2.396e+11   
+        0.196350985201453
+       0.1491395570630482
+       0.1711747419602992
+     -0.03659893210433712
+      0.08043752976576407
+       0.1725389825419435
+   -0.0003645941290560156
+      -0.0365118749277237
+       0.1488773158249876
+       0.1971007521092858
+ 2.401e+11   
+       0.1961713012011942
+       0.1486554903240348
+       0.1714610421547131
+     -0.03640128510534005
+      0.07980755436111348
+       0.1728288877578628
+   -0.0004952176837813083
+      -0.0363136067500421
+       0.1483966110956125
+       0.1969227241865718
+ 2.406e+11   
+       0.1959876283492557
+       0.1481783072981651
+       0.1717296347868019
+      -0.0362121360959397
+      0.07919424169242709
+       0.1731011084194386
+   -0.0006220536639560785
+     -0.03612382191780619
+       0.1479228086119054
+       0.1967407298774846
+ 2.411e+11   
+       0.1958006803758153
+       0.1477088789635264
+       0.1719818905947007
+     -0.03603066093350757
+      0.07859712827708677
+       0.1733569979472497
+    -0.000745563247735058
+     -0.03594170377610767
+       0.1474567691123725
+       0.1965554761206618
+ 2.416e+11   
+       0.1956111297093427
+       0.1472480061730952
+       0.1722191006093284
+     -0.03585608597825519
+      0.07801577025011572
+       0.1735978312707555
+   -0.0008661764229420104
+      -0.0357664857014128
+       0.1469992837542545
+       0.1963676288702685
+ 2.421e+11   
+       0.1954196067560719
+       0.1467964180523633
+       0.1724424772436135
+     -0.03568768764533372
+      0.07744974151878593
+       0.1738248059239413
+   -0.0009842922323828778
+     -0.03559745064360571
+       0.1465510725407072
+       0.1961778123958235
+ 2.426e+11   
+       0.1952266994271773
+       0.1463547709937143
+       0.1726531555908129
+     -0.03552479177362988
+      0.07689863205873805
+       0.1740390433434985
+      -0.0011002791641429
+       -0.035433930487982
+       0.1461127833395182
+       0.1959866088267586
+ 2.431e+11   
+       0.1950329529025364
+        0.145923648207723
+        0.172852194917581
+     -0.03536677282414852
+      0.07636204634492101
+       0.1742415903555913
+    -0.001214475675962655
+      -0.0352753052499177
+       0.1456849914537272
+       0.1957945579306484
+ 2.436e+11   
+       0.1948388696193379
+        0.145503559791661
+       0.1730405803372288
+     -0.03521305292101992
+      0.07583960191090378
+       0.1744334208370772
+    -0.001327190842642025
+     -0.03512100211506613
+       0.1452681997046329
+       0.1956021571134373
+ 2.441e+11   
+       0.1946449094733312
+       0.1450949432757694
+       0.1732192246486297
+     -0.03506310074824779
+      0.07533092803038428
+       0.1746154375370659
+    -0.001438705115303359
+     -0.03497049433800475
+       0.1448628389879546
+       0.1954098616295193
+ 2.446e+11   
+         0.19445149022005
+       0.1446981646083709
+       0.1733889703262675
+     -0.03491643031519785
+      0.07483566451496713
+       0.1747884740446885
+    -0.001549271181381469
+     -0.03482330001218858
+       0.1444692692644417
+       0.1952180849891241
+ 2.451e+11   
+       0.1942589880631116
+       0.1443135195415217
+       0.1735505916470481
+     -0.03477259960379287
+      0.07435346062253334
+       0.1749532968891466
+    -0.001659114914286895
+     -0.03467898072395286
+       0.1440877809468803
+       0.1950271995502043
+ 2.456e+11   
+       0.1940677384164709
+       0.1439412353797418
+       0.1737047969396406
+     -0.03463120911011765
+      0.07388397407068875
+       0.1751106077581706
+    -0.001768436401849928
+     -0.03453714010312198
+       0.1437185966462512
+       0.1948375372818042
+ 2.461e+11   
+       0.1938780368274153
+       0.1435814730552981
+       0.1738522309424019
+     -0.03449190029292337
+      0.07342687015003833
+       0.1752610458213533
+    -0.001877411042896003
+      -0.0343974222825114
+       0.1433618732407758
+       0.1946493906858243
+ 2.466e+11   
+       0.1936901400470453
+        0.143234329494543
+       0.1739934772561911
+     -0.03435435394120601
+      0.07298182093217205
+       0.1754051901450272
+    -0.001986190701557332
+     -0.03425951027833887
+       0.1430177042325833
+       0.1944630138640469
+ 2.471e+11   
+       0.1935042672350188
+       0.1428998402410154
+       0.1741290608787052
+     -0.03421828847264216
+      0.07254850456744903
+       0.1755435621857233
+    -0.002094904909292282
+     -0.03412312430313852
+       0.1426861223579834
+       0.1942786237173437
+ 2.476e+11   
+       0.1933206012855039
+       0.1425779823022123
+       0.1742594508073625
+     -0.03408345817433323
+      0.07212660466778752
+        0.175676628349549
+     -0.00220366210493725
+     -0.03398802002247551
+       0.1423671024184631
+       0.1940964012641215
+ 2.481e+11   
+       0.1931392902613834
+       0.1422686771882566
+       0.1743850626981388
+     -0.03394965139681979
+      0.07171580976985685
+       0.1758048026052925
+    -0.002312550903529943
+     -0.03385398676623835
+       0.1420605643009254
+       0.1939164930652104
+ 2.486e+11   
+       0.1929604489240362
+       0.1419717941120695
+       0.1745062615681939
+      -0.0338166887118871
+      0.07131581287416518
+       0.1759284491393789
+    -0.002421641385079623
+     -0.03372084570489228
+       0.1417663761569835
+       0.1937390127426416
+ 2.491e+11   
+       0.1927841603462644
+       0.1416871533220272
+       0.1746233645305833
+     -0.03368442104423093
+       0.0709263110556813
+       0.1760478850413539
+    -0.002530986394939488
+     -0.03358844800057418
+       0.1414843577125877
+       0.1935640425800485
+ 2.496e+11   
+       0.1926104775962666
+       0.1414145295395654
+       0.1747366435498195
+     -0.03355272778650201
+      0.07054700514173498
+        0.176163383008912
+    -0.002640622847886905
+     -0.03345667294242933
+       0.1412142836806337
+       0.1933916351927065
+ 2.501e+11   
+       0.1924394254809168
+       0.1411536554756303
+       0.1748463282075247
+     -0.03342151490678705
+      0.07017759945304117
+       0.1762751740620625
+    -0.002750573028547365
+      -0.0333254260750754
+       0.1409558872507296
+       0.1932218152556297
+ 2.506e+11   
+       0.1922710023369691
+       0.1409042254013531
+       0.1749526084679498
+     -0.03329071305701835
+      0.06981780160382856
+       0.1763834502564552
+    -0.002860845881256895
+     -0.03319463732856397
+       0.1407088636317111
+       0.1930545812784874
+ 2.511e+11   
+       0.1921051818592771
+        0.140665898749835
+       0.1750556374335988
+     -0.03316027569032734
+      0.06946732235708913
+       0.1764883673863999
+    -0.002971438283027168
+      -0.0330642591577085
+       0.1404728736240153
+       0.1928899074165538
+ 2.516e+11   
+       0.1919419149554795
+       0.1404383037273384
+        0.175155534081737
+     -0.03303017719478556
+      0.06912587553112441
+       0.1765900476686147
+    -0.003082336293705529
+     -0.03293426469810085
+       0.1402475472004475
+       0.1927277453073077
+ 2.521e+11   
+       0.1917811316171648
+       0.1402210409137399
+       0.1752523859730933
+     -0.03290041105049391
+      0.06879317795358526
+       0.1766885823982423
+    -0.003193516378008058
+     -0.03280464594564166
+       0.1400324870753814
+       0.1925680259227836
+ 2.526e+11   
+       0.1916227427978942
+       0.1400136868334775
+       0.1753462519245712
+     -0.03277098801641157
+      0.06846894945934927
+       0.1767840345691816
+    -0.003304946594551774
+     -0.03267541196590004
+       0.1398272722438345
+       0.1924106614282473
+ 2.531e+11   
+       0.1914666422890513
+        0.139815797479656
+       0.1754371646382834
+     -0.03264193435287917
+      0.06815291292860676
+       0.1768764414512925
+     -0.00341658774751775
+     -0.03254658713908283
+        0.139631461473298
+       0.1922555470382245
+ 2.536e+11   
+       0.1913127085849032
+       0.1396269117754232
+       0.1755251332797888
+     -0.03251329008520078
+      0.06784479436164742
+       0.1769658171175145
+    -0.003528394497083054
+     -0.03241820944594042
+       0.1394445967325939
+        0.192102562861452
+ 2.541e+11   
+        0.191160806728835
+       0.1394465549580306
+       0.1756101459988806
+     -0.03238510731323603
+      0.06754432298689901
+       0.1770521549144615
+    -0.003640316425181139
+     -0.03229032879941787
+       0.1392662065433573
+       0.1919515757267734
+ 2.546e+11   
+       0.1910107901331528
+       0.1392742418723686
+       0.1756921723867922
+     -0.03225744857141091
+      0.06725123139885299
+       0.1771354298705291
+    -0.003752299053654054
+      -0.0321630054263982
+        0.139095809241114
+       0.1918024409825486
+ 2.551e+11   
+       0.1908625023654278
+       0.1391094801620195
+       0.1757711658641906
+      -0.0321303852431546
+      0.06696525572259872
+       0.1772156010360361
+    -0.003864284812270667
+     -0.03203630830344569
+       0.1389329161341352
+       0.1916550042626048
+ 2.556e+11   
+        0.190715778894817
+       0.1389517733471498
+       0.1758470659948013
+     -0.03200399603327236
+      0.06668613580176568
+       0.1772926137504127
+    -0.003976213954518245
+     -0.03191031364997478
+       0.1387770345495633
+       0.1915091032122974
+ 2.561e+11   
+       0.1905704487923021
+        0.138800623779743
+       0.1759198007199952
+     -0.03187836550134105
+      0.06641361540673918
+       0.1773664018318613
+    -0.004088025419469007
+     -0.03178510348190511
+       0.1386276707574163
+       0.1913645691687257
+ 2.566e+11   
+       0.1904263363793137
+       0.1386555354678198
+       0.1759892885101131
+     -0.03175358265885152
+      0.06614744246013349
+       0.1774368896854451
+    -0.004199657638424668
+     -0.03166076422837908
+        0.138484332764296
+       0.1912212287896325
+ 2.571e+11   
+       0.1902832628196568
+       0.1385160167614438
+        0.176055440428793
+     -0.03162973963233646
+      0.06588736927654809
+       0.1775039943259135
+    -0.004311049285400984
+     -0.03153738541381811
+       0.1383465329696564
+       0.1910789056260194
+ 2.576e+11   
+       0.1901410476501635
+       0.1383815828942897
+       0.1761181621069477
+     -0.03150693039443992
+      0.06563315281375832
+       0.1775676273120734
+    -0.004422139970834128
+     -0.03141505840712944
+       0.1382137906785876
+       0.1909374216339696
+ 2.581e+11   
+       0.1899995102459485
+       0.1382517583756408
+       0.1761773556235112
+      -0.0313852495644529
+      0.06538455493253424
+       0.1776276965898532
+    -0.004532870878275033
+     -0.03129387523961297
+       0.1380856344660253
+        0.190796598621634
+ 2.586e+11   
+       0.1898584712166046
+        0.138126079228566
+       0.1762329212904543
+     -0.03126479127955231
+      0.06514134266242144
+       0.1776841082416863
+    -0.004643185344077097
+     -0.03117392749270852
+       0.1379616043882723
+       0.1906562596277855
+ 2.591e+11   
+       0.1897177537301157
+       0.1380040950709714
+        0.176284759339978
+      -0.0311456481376141
+      0.06490328847087537
+       0.1777367681401404
+    -0.004753029380399239
+     -0.03105530525645857
+       0.1378412540385785
+       0.1905162302287848
+ 2.596e+11   
+       0.1895771847617104
+       0.1378853710370568
+       0.1763327715121419
+     -0.03102791021223573
+      0.06467017053321972
+       0.1777855835041451
+    -0.004862352142124246
+      -0.0309380961592478
+       0.1377241524444073
+       0.1903763397712202
+ 2.601e+11   
+       0.1894365962652396
+        0.137769489537499
+       0.1763768625415892
+     -0.03091166414025032
+      0.06444177300103546
+       0.1778304643564894
+     -0.00497110633850483
+     -0.03082238446911184
+       0.1376098858047708
+       0.1902364225278972
+ 2.606e+11   
+       0.1892958262651321
+       0.1376560518574621
+       0.1764169415423335
+     -0.03079699228178381
+      0.06421788626665913
+       0.1778713248816087
+    -0.005079248590565199
+     -0.03070825026662594
+       0.1374980590667735
+       0.1900963187752265
+ 2.611e+11   
+       0.1891547198672948
+        0.137544679592194
+        0.176452923289917
+     -0.03068397195270015
+      0.06399830722153223
+       0.1779080846829876
+     -0.00518673973555713
+     -0.03059576868919347
+       0.1373882973412139
+       0.1899558757904709
+ 2.616e+11   
+       0.1890131301877294
+       0.1374350159206486
+       0.1764847294005773
+     -0.03057267472897393
+      0.06378283950632867
+       0.1779406699398381
+      -0.0052935450798502
+     -0.03048500924627221
+       0.1372802471576823
+       0.1898149487676064
+ 2.621e+11   
+       0.1888709191979633
+       0.1373267267181772
+       0.1765122894073069
+     -0.03046316582239433
+      0.06357129375076195
+       0.1779690144629374
+    -0.005399634601908219
+     -0.03037603520492476
+       0.1371735775602587
+       0.1896734016509626
+ 2.626e+11   
+       0.1887279584867181
+       0.1372195015098538
+       0.1765355417330323
+     -0.03035550352676972
+      0.06336348780120134
+       0.1779930606498649
+    -0.005504983107061464
+     -0.03026890304485939
+       0.1370679810454058
+       0.1895311078860895
+ 2.631e+11   
+       0.1885841299375673
+       0.1371130542665584
+       0.1765544345613465
+     -0.03024973873364164
+      0.06315924693422278
+       0.1780127603400454
+    -0.005609570335975449
+     -0.03016366198196485
+        0.136963174344178
+       0.1893879510875911
+ 2.636e+11   
+       0.1884393263226109
+       0.1370071240463656
+       0.1765689266054962
+     -0.03014591451636452
+      0.06295840405437092
+       0.1780280755703128
+    -0.005713381028794831
+     -0.03006035355919832
+       0.1368588990513399
+       0.1892438256240155
+ 2.641e+11   
+       0.1882934518124627
+       0.1369014754842426
+       0.1765789877765704
+      -0.0300440657812538
+      0.06276079987450761
+       0.1780389792318982
+    -0.005816404947082288
+     -0.02995901130352664
+       0.1367549221043829
+       0.1890986371200727
+ 2.646e+11   
+        0.188146422403138
+       0.1367958991334101
+       0.1765845997520121
+     -0.02994421898438297
+      0.06256628307719375
+       0.1780454556299543
+    -0.005918636855677964
+     -0.02985966044751812
+       0.1366510361158031
+       0.1889523028767838
+ 2.651e+11   
+       0.1879981662606068
+       0.1366902116620899
+       0.1765857564458174
+     -0.02984639191248628
+      0.06237471045568332
+       0.1780475009469355
+    -0.006020076466759207
+      -0.0297623177140433
+       0.1365470595623728
+       0.1888047522103568
+ 2.656e+11   
+       0.1878486239840842
+       0.1365842559096692
+       0.1765824643819313
+     -0.02975059352634422
+      0.06218594703317491
+       0.1780451236113208
+    -0.006120728348382773
+     -0.02966699116247016
+       0.1364428368354035
+       0.1886559267108058
+ 2.661e+11   
+       0.1876977487892473
+        0.136477900806556
+       0.1765747429725589
+     -0.02965682386490523
+      0.06199986615909724
+        0.178038344573339
+    -0.006220601799835771
+     -0.02957368009464969
+       0.1363382381562833
+       0.1885057804215708
+ 2.666e+11   
+       0.1875455066128215
+       0.1363710411622359
+       0.1765626247032104
+     -0.02956507400838286
+      0.06181634958126245
+       0.1780271974894952
+    -0.006319710696172668
+     -0.02948237501888924
+       0.1362331593617851
+       0.1883542799415036
+ 2.671e+11   
+       0.1873918761401239
+        0.136263597326301
+       0.1765461552265025
+     -0.02947532609841503
+      0.06163528749285376
+       0.1780117288178492
+    -0.006418073304318544
+     -0.02939305767009478
+       0.1361275215638625
+       0.1882014044508502
+ 2.676e+11   
+       0.1872368487573124
+       0.1361555147272965
+       0.1765253933668265
+     -0.02938755341340286
+       0.0614565785532887
+       0.1779919978260978
+     -0.00651571207310364
+     -0.02930570108416026
+       0.1360212706887892
+       0.1880471456629377
+ 2.681e+11   
+       0.1870804284302292
+       0.1360467632944451
+       0.1765004110381037
+     -0.02930172049706867
+      0.06128012988208568
+       0.1779680765146722
+    -0.006612653399655745
+     -0.02922026972468207
+       0.1359143769006725
+       0.1878915077034549
+ 2.686e+11   
+       0.1869226315118808
+       0.1359373367674175
+       0.1764712930769907
+     -0.02921778333821549
+      0.06110585702496994
+       0.1779400494570828
+    -0.006708927374479335
+     -0.02913671966003411
+       0.1358068339144285
+       0.1877345069193253
+ 2.691e+11   
+       0.1867634864806596
+       0.1358272518993464
+       0.1764381369939354
+      -0.0291356895997021
+      0.06093368389153069
+       0.1779080135599258
+    -0.006804567507592698
+     -0.02905499878878539
+        0.135698658203461
+        0.187576171619295
+ 2.696e+11   
+       0.1866030336115565
+       0.1357165475584308
+       0.1764010526446147
+     -0.02905537889456514
+       0.0607635426638351
+       0.1778720777449479
+    -0.006899610438042336
+     -0.02897504711149004
+        0.135589888107275
+       0.1874165417484387
+ 2.701e+11   
+       0.1864413245827098
+       0.1356052837334435
+       0.1763601618243125
+     -0.02897678310729727
+      0.06059537367547826
+        0.177832362555733
+    -0.006994095629074742
+     -0.02889679704680682
+       0.1354805828443584
+       0.1872556684988964
+ 2.706e+11   
+        0.186278422019631
+       0.1354935404485223
+       0.1763155977878772
+     -0.02889982675816937
+      0.06042912526065063
+       0.1777889996915144
+    -0.007088065051200322
+      -0.0288201737899477
+       0.1353708214356241
+       0.1870936138591948
+ 2.711e+11   
+       0.1861143989796486
+       0.1353814165926032
+        0.176267504697936
+     -0.02882442740863779
+      0.06026475357286377
+        0.177742131470794
+    -0.007181562855353646
+     -0.02874509571143754
+        0.135260701543772
+       0.1869304501046107
+ 2.716e+11   
+       0.1859493383790019
+       0.1352690286688454
+       0.1762160370040909
+      -0.0287504961057371
+      0.06010222237306359
+       0.1776919102273468
+    -0.007274635038278028
+     -0.02867147479420727
+       0.1351503382338262
+       0.1867662592310439
+ 2.721e+11   
+       0.1857833323652125
+       0.1351565094693464
+       0.1761613587558399
+      -0.0286779378635195
+      0.05994150278693345
+        0.177638497641364
+    -0.007367329102212019
+     -0.02859921710702528
+       0.1350398626601516
+       0.1866011323349424
+ 2.726e+11   
+       0.1856164816372716
+       0.1350440066804378
+       0.1761036428519951
+     -0.02860665217949246
+       0.0597825730312625
+        0.177582064008362
+    -0.007459693710900907
+     -0.02852822331232243
+       0.1349294206851361
+       0.1864351689418207
+ 2.731e+11   
+       0.1854488947162874
+       0.1349316814237355
+       0.1760430702293876
+     -0.02853653358413591
+      0.05962541810932762
+       0.1775227874486343
+    -0.007551778343866641
+     -0.02845838920646935
+       0.1348191714347134
+       0.1862684762859669
+ 2.736e+11   
+       0.1852806871691816
+       0.1348197067380524
+       0.1759798289936221
+     -0.02846747222157306
+      0.05947002947528551
+       0.1774608530599211
+     -0.00764363295083449
+     -0.02838960629063428
+       0.1347092857957742
+        0.186101168543926
+ 2.741e+11   
+       0.1851119807881181
+       0.1347082660072768
+       0.1759141134947214
+     -0.02839935445945183
+      0.05931640466767839
+       0.1773964520160411
+    -0.007735307608098094
+     -0.02832176237032954
+       0.1345999448604694
+       0.1859333660243569
+ 2.746e+11   
+       0.1849429027282287
+       0.1345975513390433
+       0.1758461233503732
+     -0.02833206352626363
+      0.05916454691214523
+       0.1773297806141706
+    -0.007826852178574505
+     -0.02825474218184944
+       0.1344913383222726
+       0.1857651943168525
+ 2.751e+11   
+       0.1847735846063127
+       0.1344877618991463
+       0.1757760624196095
+     -0.02826548017419284
+      0.05901446469359561
+       0.1772610392735015
+    -0.007918315977192473
+     -0.02818842804378582
+       0.1343836628286096
+       0.1855967834023225
+ 2.756e+11   
+       0.1846041615630723
+        0.134379102206305
+        0.175704137729626
+     -0.02819948336580114
+      0.05886617129803799
+       0.1771904314879227
+    -0.008009747443188222
+     -0.02812270053191599
+       0.1342771202946769
+       0.1854282667274963
+ 2.761e+11   
+        0.184434771291488
+        0.134271780391946
+       0.1756305583584742
+     -0.02813395098277042
+      0.05871968432440475
+        0.177118162735408
+    -0.008101193820815328
+     -0.02805743917572715
+       0.1341719161830422
+       0.1852597802461056
+ 2.766e+11   
+       0.1842655530338736
+       0.1341660064294287
+       0.1755555342763334
+     -0.02806876055504696
+      0.05857502516671747
+       0.1770444393467149
+    -0.008192700849882604
+     -0.02799252317496993
+        0.134068257753383
+       0.1850914614292468
+ 2.771e+11   
+       0.1840966465501336
+       0.1340619903370432
+       0.1754792751480043
+     -0.02800379000875466
+      0.05843221846699509
+       0.1769694673360111
+    -0.008284312467451552
+     -0.02792783213460222
+       0.1339663522866955
+       0.1849234482474424
+ 2.776e+11   
+       0.1839281910597224
+       0.1339599403590092
+       0.1754019890992584
+     -0.02793891843128456
+      0.05829129153934803
+       0.1768934511959669
+    -0.008376070521970544
+     -0.02786324681659513
+       0.1338664052880837
+       0.1847558781268106
+ 2.781e+11   
+       0.1837603241597151
+       0.1338600611284823
+       0.1753238814496218
+     -0.02787402685203676
+       0.0581522737657602
+       0.1768165926598413
+    -0.008468014501003353
+      -0.0277986499070858
+       0.1337686186721481
+       0.1845888868817873
+ 2.786e+11   
+       0.1835931807214092
+        0.133762551816492
+       0.1752451534141274
+     -0.02780899903734391
+      0.05801519596407539
+       0.1767390894330466
+    -0.008560181273669119
+      -0.0277339267974407
+       0.1336731889348181
+       0.1844226076267443
+ 2.791e+11   
+       0.1834268917677877
+       0.1336676042705882
+       0.1751660007765286
+     -0.02774372229812998
+      0.05788008972874998
+       0.1766611338965916
+    -0.008652604848821133
+     -0.02766896637781706
+       0.1335803053153622
+       0.1842571696688212
+ 2.796e+11   
+       0.1832615833341492
+       0.1335754011467919
+       0.1750866125364213
+     -0.02767808830893525
+      0.05774698674500448
+       0.1765829117848255
+     -0.00874531614989338
+     -0.02760366184186809
+       0.1334901479521269
+       0.1840926973842251
+ 2.801e+11   
+       0.1830973753141332
+       0.1334861140383153
+       0.1750071695326402
+     -0.02761199393699879
+      0.05761591807694545
+       0.1765046008397622
+    -0.008838342807308794
+     -0.02753791150132931
+       0.1334028860354219
+       0.1839293090802271
+ 2.806e+11   
+       0.1829343802933069
+       0.1333999016043635
+       0.1749278430452785
+     -0.02754534208010393
+      0.05748691343038277
+       0.1764263694443089
+    -0.008931708969231896
+      -0.0274716196091911
+        0.133318675960834
+       0.1837671158449679
+ 2.811e+11   
+       0.1827727023724674
+       0.1333169077022043
+       0.1748487933786109
+     -0.02747804251197992
+      0.05736000039099222
+       0.1763483752366011
+    -0.009025435131398843
+     -0.02740469719029923
+       0.1332376594860903
+       0.1836062203872011
+ 2.816e+11   
+       0.1826124359826787
+       0.1332372595255076
+       0.1747701684271203
+     -0.02741001273408985
+      0.05723520363852258
+       0.1762707637075839
+    -0.009119537986695198
+     -0.02733706287823972
+       0.1331599618944398
+       0.1834467158679792
+ 2.821e+11   
+       0.1824536646940653
+       0.1331610657518277
+       0.1746921022268161
+     -0.02734117883268628
+      0.05711254413784531
+       0.1761936667840184
+    -0.009214030295041692
+     -0.02726864375738266
+       0.1330856901673874
+       0.1832886847262462
+ 2.826e+11   
+       0.1822964600202674
+       0.1330884147019561
+       0.1746147134938962
+     -0.02727147634006553
+      0.05699203830750473
+       0.1761172013988689
+    -0.009308920774140984
+     -0.02719937620908042
+       0.1330149311694729
+       0.1831321975002582
+ 2.831e+11   
+       0.1821408802204428
+       0.1330193725137366
+       0.1745381041528526
+     -0.02720085109899916
+      0.05687369716663335
+        0.176041468051151
+    -0.009404214011521897
+     -0.02712920676099444
+       0.1329477498476247
+       0.1829773116466413
+ 2.836e+11   
+       0.1819869691005817
+        0.132953981332762
+        0.174462357855953
+     -0.02712926012938695
+      0.05675752546096273
+       0.1759665493571224
+    -0.009499910398307734
+     -0.02705809293862252
+       0.1328841874475087
+       0.1828240703588818
+ 2.841e+11   
+       0.1818347548159076
+       0.1328922575222786
+       0.1743875384960247
+     -0.02705667249618785
+      0.05664352076874668
+       0.1758925085946936
+     -0.00959600608500495
+      -0.0269860041181098
+       0.1328242597491162
+       0.1826725013869362
+ 2.846e+11   
+       0.1816842486759624
+       0.1328341898944413
+       0.1743136887144047
+     -0.02698307017777376
+      0.05653167258741212
+       0.1758193882428863
+    -0.009692492959653789
+      -0.0269129223795052
+       0.1327679553237419
+       0.1825226158595991
+ 2.851e+11   
+       0.1815354439540312
+       0.1327797379649684
+       0.1742408284058417
+     -0.02690844893386311
+       0.0564219614017652
+       0.1757472085180743
+    -0.009789358648520078
+     -0.02683884335963682
+        0.132715233814323
+       0.1823744071111952
+ 2.856e+11   
+       0.1813883147023714
+       0.1327288302330681
+       0.1741689532220713
+     -0.02683281917225563
+      0.05631435773457546
+       0.1756759659087225
+    -0.009886586539530976
+     -0.02676377710384494
+       0.1326660242410417
+       0.1822278495141138
+ 2.861e+11   
+       0.1812428145747502
+       0.1326813624884601
+       0.1740980330757485
+     -0.02675620681361698
+      0.05620882118036898
+       0.1756056317101964
+    -0.009984155828598362
+     -0.02668774891586589
+       0.1326202233338827
+       0.1820828973185811
+ 2.866e+11   
+       0.1810988756576221
+       0.1326371961470581
+       0.1740280106463251
+     -0.02667865415363105
+       0.0561052994233102
+       0.1755361505613137
+     -0.01008204158888117
+      -0.0266108002051433
+       0.1325776938938192
+       0.1819394835010745
+ 2.871e+11   
+       0.1809564073113164
+       0.1325961566169332
+       0.1739587998894417
+      -0.0266002207218404
+      0.05600372723996514
+       0.1754674389840379
+     -0.01018021486307128
+     -0.02653298933098077
+       0.1325382631840678
+       0.1817975186226464
+ 2.876e+11   
+       0.1808152950224399
+       0.1325580316958942
+       0.1738902845512914
+     -0.02652098413656846
+      0.05590402548784578
+       0.1753993839278541
+      -0.0102786427786755
+     -0.02645439244287168
+       0.1325017213528492
+       0.1816568896983994
+ 2.881e+11   
+       0.1806753992687038
+       0.1325225700020167
+       0.1738223166894116
+     -0.02644104095534783
+      0.05580610008055086
+       0.1753318413201788
+     -0.01037728868628052
+     -0.02637510431649931
+       0.1324678198888726
+       0.1815174590792748
+ 2.886e+11   
+       0.1805365543972541
+       0.1324894794382933
+       0.1737547152012403
+     -0.02636050752028542
+      0.05570984095036972
+       0.1752646346241504
+     -0.01047611232071977
+     -0.02629523918483245
+       0.1324362701107426
+       0.1813790633472485
+ 2.891e+11   
+       0.1803985675176026
+       0.1324584256924933
+       0.1736872643617744
+      -0.0262795207978989
+      0.05561512099919741
+       0.1751975534050973
+     -0.01057506998505846
+     -0.02621493156384674
+         0.13240674169132
+       0.1812415122249514
+ 2.896e+11   
+       0.1802612174100753
+       0.1324290307731846
+       0.1736197123715672
+     -0.02619823921292341
+      0.05552179503858923
+        0.175130351906899
+     -0.01067411475726302
+     -0.02613433707242135
+       0.1323788612180042
+       0.1811045875007188
+ 2.901e+11   
+       0.1801242534507486
+       0.1324008715828355
+       0.1735517699162629
+     -0.02611684347564263
+      0.05542969871981499
+       0.1750627476393911
+       -0.010773196719391
+     -0.02605363324596157
+       0.1323522107897671
+       0.1809680419699066
+ 2.906e+11   
+       0.1799873945536897
+       0.1323734785287277
+        0.173483108738815
+     -0.02603553740238549
+      0.05533864745474483
+       0.1749944199780055
+     -0.01087226320915248
+     -0.02597302034336465
+       0.1323263266517498
+       0.1808315983933735
+ 2.911e+11   
+       0.1798503281312976
+        0.132346334172415
+       0.1734133602254835
+     -0.02595454872875155
+      0.05524843532838607
+       0.1749250087766167
+     -0.01097125909361009
+     -0.02589272214698179
+       0.1323006978680252
+       0.1806949484738625
+ 2.916e+11   
+       0.1797127090734678
+       0.1323188719182883
+       0.1733421140066256
+     -0.02587412991528353
+      0.05515883400390784
+       0.1748541129946959
+     -0.01107012706483264
+     -0.02581298675522129
+       0.1322747650331657
+       0.1805577518510089
+ 2.921e+11   
+       0.1795741587462527
+       0.1322904747418035
+       0.1732689165732918
+     -0.02579455894522167
+      0.05506959162096373
+       0.1747812893396854
+     -0.01116880795723684
+     -0.02573408736749772
+       0.1322479190230823
+       0.1804196351156252
+ 2.926e+11   
+       0.1794342640106034
+       0.1322604739577742
+       0.1731932699105442
+     -0.02571614011408323
+      0.05498043168812041
+       0.1747060509255317
+     -0.01126724108638944
+      -0.0256563230612518
+       0.1322194997855702
+       0.1802801908438533
+ 2.931e+11   
+       0.1792925762617437
+       0.1322281480290899
+       0.1731146301483894
+     -0.02563920481080036
+      0.05489105197020271
+       0.1746278659482617
+     -0.01136536460898104
+     -0.02558001956078426
+       0.1321887951708953
+       0.1801389766517296
+ 2.936e+11   
+       0.1791486104896828
+       0.1321927214161698
+       0.1730324062311648
+     -0.02556411229016974
+      0.05480112337133605
+       0.1745461563793913
+     -0.01146311590370382
+     -0.02550552999767925
+       0.1321550398026837
+       0.1799955142706139
+ 2.941e+11   
+       0.1790018443612456
+       0.1321533634673081
+         0.17294595860616
+     -0.02549125043640447
+      0.05471028881447523
+       0.1744602966779645
+     -0.01156043197271135
+      -0.0254332356626047
+       0.1321174139893188
+        0.179849288643939
+ 2.946e+11   
+       0.1788517173240734
+       0.1321091873501002
+       0.1728545979322385
+     -0.02542103651760752
+       0.0546181621182003
+       0.1743696125219757
+     -0.01165724986336127
+     -0.02536354674831257
+       0.1320750426759731
+       0.1796997470456392
+ 2.951e+11   
+       0.1786976297328554
+       0.1320592490239942
+       0.1727575838091314
+     -0.02535391793096833
+      0.05452432687152626
+       0.1742733795597982
+     -0.01175350710989138
+     -0.02529690308367403
+        0.132026994437311
+       0.1795462982205599
+ 2.956e+11   
+       0.1785389419981036
+       0.1320025462539537
+       0.1726541235280812
+     -0.02529037293854882
+      0.05442833530752415
+       0.1741708221823549
+     -0.01184914219464332
+     -0.02523377485857007
+        0.131972280510891
+       0.1793883115471542
+ 2.961e+11   
+       0.1783749737577037
+       0.1319380176652171
+       0.1725433708444276
+     -0.02523091139349288
+      0.05432970717646148
+       0.1740611123165495
+     -0.01194409502846388
+     -0.02517466333954149
+       0.1319098538711723
+       0.1792251162226782
+ 2.966e+11   
+       0.1782050030714213
+       0.1318645418389866
+       0.1724244247727207
+     -0.02517607545653825
+      0.05422792861923637
+       0.1739433682405564
+     -0.01203830744982318
+     -0.02512010157604141
+       0.1318386083439924
+       0.1790560004710703
+ 2.971e+11   
+       0.1780282656385208
+       0.1317809364488681
+       0.1722963284048456
+     -0.02512644030269375
+      0.05412245104184406
+       0.1738166534214843
+     -0.01213172374215302
+     -0.02507065509715455
+       0.1317573777613418
+       0.1788802107736705
+ 2.976e+11   
+       0.1778439540386452
+        0.131685957437835
+       0.1721580677516826
+     -0.02508261481795288
+       0.0540126899916064
+       0.1736799753758603
+     -0.01222429116885393
+     -0.02502692259869588
+       0.1316649351561431
+       0.1786969511229027
+ 2.981e+11   
+       0.1776512169959925
+        0.131578298235349
+       0.1720085706086844
+     -0.02504524228591879
+       0.0538980240359006
+        0.173532284553376
+     -0.01231596052533503
+     -0.02498953662053417
+       0.1315599919967469
+       0.1785053822990138
+ 2.986e+11   
+       0.1774491586669423
+       0.1314565890143165
+       0.1718467054457867
+     -0.02501500106418466
+      0.05377779364415961
+        0.173372473244267
+     -0.01240668670732403
+     -0.02495916421400251
+        0.131441197460722
+        0.178304621169921
+ 2.991e+11   
+       0.1772368379511153
+       0.1313193959873581
+       0.1716712803219403
+      -0.0249926052503248
+      0.05365130007383612
+        0.173199374510648
+     -0.01249642929458667
+     -0.02493650759924297
+       0.1313071377475247
+       0.1780937400142778
+ 2.996e+11   
+       0.1770132678259788
+       0.1311652207419341
+       0.1714810418245921
+     -0.02497880533727745
+      0.05351780426115117
+       0.1730117611420673
+     -0.01258515314901785
+     -0.02492230481230144
+        0.131156335429458
+       0.1778717658677401
* NOTE: Solution at 1e+08 Hz used as DC point.
* NOTE: Repaired negative diagonal entries at these frequencies:
* 1.7e+11 Hz, 1.8e+11 Hz, 1.8e+11 Hz, 1.8e+11 Hz, 1.8e+11 Hz, 1.8e+11 Hz,
* 1.8e+11 Hz, 1.8e+11 Hz, 1.8e+11 Hz, 1.8e+11 Hz, 1.8e+11 Hz, 1.8e+11 Hz,
* 1.8e+11 Hz, 1.8e+11 Hz, 1.8e+11 Hz, 1.8e+11 Hz, 1.8e+11 Hz, 1.8e+11 Hz,
* 1.8e+11 Hz, 1.8e+11 Hz, 1.8e+11 Hz, 1.9e+11 Hz, 1.9e+11 Hz, 1.9e+11 Hz,
* 1.9e+11 Hz, 1.9e+11 Hz, 1.9e+11 Hz, 1.9e+11 Hz, 1.9e+11 Hz, 1.9e+11 Hz,
* 1.9e+11 Hz, 1.9e+11 Hz, 1.9e+11 Hz, 1.9e+11 Hz, 1.9e+11 Hz, 1.9e+11 Hz,
* 1.9e+11 Hz, 1.9e+11 Hz, 1.9e+11 Hz, 1.9e+11 Hz, 1.9e+11 Hz,  2e+11 Hz,  2e+11
* Hz,  2e+11 Hz,  2e+11 Hz,  2e+11 Hz,  2e+11 Hz,  2e+11 Hz,  2e+11 Hz,  2e+11
* Hz,  2e+11 Hz,  2e+11 Hz,  2e+11 Hz,  2e+11 Hz,  2e+11 Hz,  2e+11 Hz,  2e+11
* Hz,  2e+11 Hz,  2e+11 Hz,  2e+11 Hz,  2e+11 Hz, 2.1e+11 Hz, 2.1e+11 Hz,
* 2.1e+11 Hz, 2.1e+11 Hz

.model c_m4lines_veryHighFreq_W_1 sp N=4 SPACING=nonuniform VALTYPE=real
+ INTERPOLATION=spline
+ INFINITY =
+    2.556655466176534e-11
+    9.268425817011095e-12
+    2.156998960948431e-11
+   -6.859396432269608e-12
+     9.34619274581565e-12
+    2.161768467603702e-11
+    2.632801425425317e-12
+   -6.852347032335529e-12
+    9.255230899294873e-12
+    2.558850389628505e-11
+ DATA = 600
+ 0           
+    8.534587023821072e-11
+   -2.095537631618298e-11
+    8.700278160855642e-11
+   -8.333425087446117e-13
+    -1.00146231354576e-11
+    8.700833294804957e-11
+   -3.001520909585882e-13
+   -8.340223463885308e-13
+   -2.095267790319996e-11
+    8.533136511217923e-11
+ 6e+08       
+    8.382832960109412e-11
+   -2.067707140972717e-11
+    8.547535367610619e-11
+   -8.294020486188888e-13
+   -9.894210167572235e-12
+    8.548076777391741e-11
+   -2.987086909803617e-13
+   -8.300937867507662e-13
+   -2.067467792287946e-11
+    8.381465318278806e-11
+ 1.1e+09     
+    8.334810868479389e-11
+   -2.059121934820341e-11
+    8.499214140494965e-11
+    -8.18881935820887e-13
+   -9.853726734990029e-12
+    8.499750421513857e-11
+     -2.9435584249241e-13
+   -8.195798034256017e-13
+   -2.058893794930097e-11
+     8.33347521669252e-11
+ 1.6e+09     
+    8.308595056965689e-11
+   -2.054921651409513e-11
+    8.472919813150369e-11
+   -7.961551364103809e-13
+   -9.825204700011652e-12
+    8.473449090041724e-11
+   -2.851862193011009e-13
+   -7.968995291213799e-13
+   -2.054702749682081e-11
+    8.307294963589833e-11
+ 2.1e+09     
+     8.28512439568956e-11
+   -2.048994652363002e-11
+    8.449054545466936e-11
+   -7.834588666982741e-13
+   -9.791677048883485e-12
+    8.449581031284603e-11
+   -2.743821175161544e-13
+   -7.842476286218247e-13
+   -2.048779979641761e-11
+    8.283840651774569e-11
+ 2.6e+09     
+    8.266210617938783e-11
+   -2.043290074231705e-11
+    8.429640740127586e-11
+   -7.752127415642067e-13
+   -9.761858411496454e-12
+    8.430168081181285e-11
+   -2.640525590744896e-13
+   -7.760247250275329e-13
+   -2.043077314128556e-11
+    8.264930841709244e-11
+ 3.1e+09     
+    8.251435251111614e-11
+   -2.038301173796945e-11
+    8.414352987488794e-11
+   -7.689887653279709e-13
+   -9.736916161674159e-12
+    8.414883214137587e-11
+   -2.548391596061061e-13
+   -7.698090128740904e-13
+   -2.038089537381567e-11
+    8.250153916162057e-11
+ 3.6e+09     
+    8.239836258992773e-11
+   -2.034019481181515e-11
+    8.402261604313476e-11
+   -7.636870209622401e-13
+   -9.715783785898967e-12
+     8.40279553488723e-11
+   -2.468158155898402e-13
+   -7.645071112212154e-13
+    -2.03380886623147e-11
+    8.238551874874267e-11
+ 4.1e+09     
+    8.230525062018109e-11
+   -2.030315733766645e-11
+    8.392479654115126e-11
+   -7.588347837571892e-13
+   -9.696822689428766e-12
+    8.393017422701204e-11
+   -2.398999869772967e-13
+   -7.596510042865255e-13
+   -2.030106225184734e-11
+    8.229237948068277e-11
+ 4.6e+09     
+    8.222824425203734e-11
+   -2.027059584009324e-11
+    8.384319797628771e-11
+   -7.542719236393658e-13
+   -9.678478163571562e-12
+    8.384861203386318e-11
+   -2.340159966100852e-13
+   -7.550840041476279e-13
+   -2.026851198270185e-11
+    8.221535465604496e-11
+ 5.1e+09     
+    8.216253313558021e-11
+   -2.024148446949355e-11
+    8.377296767753378e-11
+   -7.499302562585699e-13
+    -9.65999364047249e-12
+    8.377841469507962e-11
+   -2.291589252611353e-13
+   -7.507405959319253e-13
+   -2.023941035768888e-11
+     8.21496337880002e-11
+ 5.6e+09     
+    8.210480230053793e-11
+   -2.021509977603933e-11
+    8.371093188004562e-11
+   -7.456899074862549e-13
+   -9.641967941573058e-12
+    8.371640815959047e-11
+   -2.254147783107254e-13
+   -7.465029873726773e-13
+   -2.021303250072621e-11
+    8.209189967140609e-11
+ 6.1e+09     
+    8.205281209092483e-11
+   -2.019099558754913e-11
+    8.365510150467174e-11
+   -7.414360003144429e-13
+   -9.625786257666624e-12
+    8.366060388732448e-11
+   -2.229401256111643e-13
+   -7.422577508242103e-13
+   -2.018893209355883e-11
+    8.203991021182806e-11
+ 6.6e+09     
+    8.200508985593444e-11
+   -2.016897970659024e-11
+    8.360417111382243e-11
+   -7.372365690601159e-13
+   -9.612371117997702e-12
+    8.360969776233471e-11
+   -2.219220562585463e-13
+   -7.380735119150832e-13
+   -2.016691888690244e-11
+    8.199219101130244e-11
+ 7.1e+09     
+    8.196070957691166e-11
+   -2.014908044040713e-11
+    8.355723159841698e-11
+   -7.334130760365638e-13
+   -9.601735251547769e-12
+    8.356278262388271e-11
+   -2.225572989336987e-13
+   -7.342710983694121e-13
+   -2.014702510752682e-11
+    8.194781515903818e-11
+ 7.6e+09     
+    8.191912435475591e-11
+   -2.013147095894043e-11
+    8.351366620036273e-11
+   -7.304981484817801e-13
+   -9.593356044004992e-12
+    8.351924362616666e-11
+   -2.250531047053712e-13
+   -7.313808954098013e-13
+   -2.012942775923138e-11
+    8.190623510090621e-11
+ 8.1e+09     
+    8.188002516537551e-11
+   -2.011632544215767e-11
+    8.347307557917038e-11
+   -7.291952063255376e-13
+   -9.586578914158917e-12
+    8.347868209629577e-11
+   -2.296333692598832e-13
+   -7.301022694473272e-13
+    -2.01143008302214e-11
+    8.186714013902343e-11
+ 8.6e+09     
+    8.184321664948838e-11
+   -2.010362656898619e-11
+    8.343517971227247e-11
+     -7.3036690358339e-13
+   -9.580781010105261e-12
+    8.344081653569816e-11
+   -2.365457605223912e-13
+   -7.312922148044405e-13
+   -2.010161986942301e-11
+    8.183033127936467e-11
+ 9.1e+09     
+    8.180852620164647e-11
+   -2.009301882755185e-11
+     8.33997296969731e-11
+   -7.350091023383221e-13
+   -9.575397441357799e-12
+    8.340539514772103e-11
+   -2.460744148580022e-13
+   -7.359404850871998e-13
+   -2.009101781328401e-11
+    8.179563108842042e-11
+ 9.6e+09     
+    8.177577132698787e-11
+   -2.008382166083421e-11
+    8.336647258133166e-11
+   -7.441536228339887e-13
+   -9.569923269574751e-12
+     8.33721629147007e-11
+   -2.585651610995137e-13
+     -7.4507573643375e-13
+   -2.008180588401553e-11
+    8.176285355896449e-11
+ 1.01e+10    
+    8.174792028917332e-11
+   -2.007645849486229e-11
+    8.333741561548465e-11
+   -7.586154709100972e-13
+   -9.563862671183487e-12
+    8.334312820101245e-11
+   -2.742972074761646e-13
+   -7.595020363130991e-13
+   -2.007443986020481e-11
+    8.173507902329415e-11
+ 1.06e+10    
+    8.173315281006399e-11
+   -2.007420095708091e-11
+    8.331824228758473e-11
+   -7.755869500410977e-13
+    -9.55725195354874e-12
+    8.332398086247457e-11
+   -2.911196704470314e-13
+   -7.763624755504483e-13
+   -2.007229176000443e-11
+     8.17207933201098e-11
+ 1.11e+10    
+    8.171818741154732e-11
+   -2.007210171493726e-11
+    8.329942625232958e-11
+   -7.931942203357452e-13
+   -9.550762035409868e-12
+    8.330519333982237e-11
+   -3.083922170363285e-13
+   -7.938493062140319e-13
+   -2.007029077827254e-11
+    8.170624834642782e-11
+ 1.16e+10    
+    8.170307242864827e-11
+   -2.007017946927337e-11
+    8.328103310846179e-11
+   -8.114150880464532e-13
+   -9.544425271377978e-12
+    8.328683125279497e-11
+   -3.260724359361411e-13
+   -8.119398919906022e-13
+   -2.006845639579663e-11
+      8.1691496476457e-11
+ 1.21e+10    
+    8.168785177268277e-11
+   -2.006845124216517e-11
+    8.326311901095233e-11
+   -8.302269726961313e-13
+   -9.538271809133296e-12
+    8.326895074222396e-11
+   -3.441176403651804e-13
+   -8.306111731944049e-13
+    -2.00668064345903e-11
+    8.167658576718575e-11
+ 1.26e+10    
+    8.167256476178837e-11
+   -2.006693246418248e-11
+    8.324573123439858e-11
+    -8.49606946178798e-13
+   -9.532329617339462e-12
+     8.32515990395896e-11
+   -3.624850135951534e-13
+   -8.498397014476823e-13
+   -2.006535712438848e-11
+    8.166155967360182e-11
+ 1.31e+10    
+    8.165724607397265e-11
+   -2.006563708544693e-11
+    8.322890879887034e-11
+   -8.695317672316122e-13
+   -9.526624534530651e-12
+    8.323481509936617e-11
+   -3.811317509695412e-13
+   -8.696016698376714e-13
+   -2.006412319899358e-11
+     8.16464569177168e-11
+ 1.36e+10    
+    8.164192580121207e-11
+   -2.006457770248247e-11
+    8.321268313177533e-11
+   -8.899779099439757e-13
+   -9.521180334526958e-12
+    8.321863026729801e-11
+   -4.000151983669946e-13
+   -8.898729372801789e-13
+   -2.006311801321701e-11
+    8.163131148363841e-11
+ 1.41e+10    
+    8.162662958383995e-11
+   -2.006376569373738e-11
+    8.319707874349162e-11
+   -9.109215848403272e-13
+   -9.516018804765535e-12
+    8.320306896213556e-11
+   -4.190929870503665e-13
+   -9.106290455334286e-13
+   -2.006235367215337e-11
+    8.161615271245698e-11
+ 1.46e+10    
+    8.161137880608285e-11
+   -2.006321135808813e-11
+    8.318211389908288e-11
+   -9.323387504987137e-13
+   -9.511159834841434e-12
+    8.318814935285246e-11
+   -4.383231650880465e-13
+   -9.318452269771719e-13
+   -2.006184116620106e-11
+    8.160100547330593e-11
+ 1.51e+10    
+    8.159619083563655e-11
+    -2.00629240515728e-11
+    8.316780127199292e-11
+   -9.542051134781048e-13
+   -9.506621513133182e-12
+    8.317388401734738e-11
+   -4.576643256398297e-13
+    -9.53496400889631e-13
+   -2.006159050638699e-11
+    8.158589038977548e-11
+ 1.56e+10    
+    8.158107929254601e-11
+   -2.006291231905552e-11
+    8.315414856946167e-11
+   -9.764961135338911e-13
+   -9.502420230311296e-12
+    8.316028057197999e-11
+   -4.770757326635741e-13
+    -9.75557155510367e-13
+   -2.006161085596174e-11
+    8.157082410400556e-11
+ 1.61e+10    
+    8.156605433489407e-11
+   -2.006318401826465e-11
+    8.314115912203317e-11
+   -9.991868907256271e-13
+   -9.498570789023961e-12
+    8.314734226465193e-11
+   -4.965174447786841e-13
+   -9.980017125705997e-13
+   -2.006191065545105e-11
+    8.155581956367806e-11
+ 1.66e+10    
+    8.155112295110528e-11
+   -2.006374643490407e-11
+    8.312883243243388e-11
+   -1.022252229823412e-12
+   -9.495086519848999e-12
+    8.313506852646607e-11
+   -5.159504384163934e-13
+   -1.020803870226772e-12
+   -2.006249773932564e-11
+    8.154088631993629e-11
+ 1.71e+10    
+    8.153628925063462e-11
+   -2.006460638810369e-11
+    8.311716468089267e-11
+   -1.045666476677589e-12
+   -9.491979404169386e-12
+    8.312345547916775e-11
+   -5.353367316353338e-13
+   -1.043936919472781e-12
+    -2.00633794433709e-11
+    8.152603082667082e-11
+ 1.76e+10    
+    8.152155474664317e-11
+   -2.006577032643371e-11
+    8.310614918586702e-11
+   -1.069403419595662e-12
+   -9.489260205357861e-12
+    8.311249639733117e-11
+   -5.546395105707755e-13
+   -1.067373527824887e-12
+   -2.006456270272124e-11
+    8.151125673376433e-11
+ 1.81e+10    
+    8.150691862574197e-11
+    -2.00672444152096e-11
+    8.309577682029314e-11
+   -1.093436127062636e-12
+   -9.486938610299503e-12
+     8.31021821253207e-11
+   -5.738232609612358e-13
+     -1.0910855826966e-12
+   -2.006605414103297e-11
+    8.149656516868454e-11
+ 1.86e+10    
+     8.14923780011836e-11
+    -2.00690346163938e-11
+    8.308603638443675e-11
+   -1.117736730972439e-12
+   -9.485023384182451e-12
+    8.309250145024282e-11
+     -5.9285390787099e-13
+   -1.115043984970945e-12
+   -2.006786015199322e-11
+     8.14819550022695e-11
+ 1.91e+10    
+    8.147792814682237e-11
+   -2.007114676297854e-11
+    8.307691493722238e-11
+   -1.142276141421158e-12
+   -9.483522542384189e-12
+    8.308344143250602e-11
+    -6.11698967742578e-13
+   -1.139218380870341e-12
+   -2.006998697478258e-11
+    8.146742309575993e-11
+ 1.96e+10    
+    8.146356270995895e-11
+   -2.007358663022592e-11
+    8.306839808827526e-11
+   -1.167023675626031e-12
+   -9.482443544428162e-12
+    8.307498769623768e-11
+   -6.303277178213545e-13
+   -1.163576817275767e-12
+   -2.007244076563297e-11
+    8.145296452696541e-11
+ 2.01e+10    
+     8.14492739016658e-11
+   -2.007636000660032e-11
+    8.306047025314159e-11
+   -1.191946578559372e-12
+   -9.481793516405889e-12
+    8.306712468171758e-11
+   -6.487113895321995e-13
+   -1.188085301877492e-12
+    -2.00752276680329e-11
+     8.14385727941815e-11
+ 2.06e+10    
+    8.143505266350645e-11
+   -2.007947276792821e-11
+    8.305311487443614e-11
+   -1.217009406885811e-12
+   -9.481579510061927e-12
+    8.305983586232899e-11
+   -6.668233940189833e-13
+   -1.212707244728249e-12
+    -2.00783538847359e-11
+    8.142423999685094e-11
+ 2.11e+10    
+    8.142088880964707e-11
+   -2.008293095889427e-11
+    8.304631461140903e-11
+     -1.2421732400203e-12
+   -9.481808808779288e-12
+    8.305310392807063e-11
+   -6.846395903176023e-13
+     -1.2374027519606e-12
+   -2.008182575515906e-11
+    8.140995699220579e-11
+ 2.16e+10    
+    8.140677114324162e-11
+   -2.008674088688921e-11
+    8.304005150057104e-11
+   -1.267394672192925e-12
+   -9.482489293669524e-12
+    8.304691093751128e-11
+   -7.021386092803236e-13
+   -1.262127734956906e-12
+    -2.00856498424494e-11
+    8.139571352716035e-11
+ 2.21e+10    
+    8.139268754566469e-11
+   -2.009090923418985e-11
+    8.303430708969706e-11
+   -1.292624527181712e-12
+   -9.483629886103215e-12
+    8.304123843977742e-11
+   -7.193022498350591e-13
+   -1.286832789393597e-12
+   -2.008983303535164e-11
+    8.138149834466183e-11
+ 2.26e+10    
+    8.137862503669303e-11
+   -2.009544319574226e-11
+    8.302906254735327e-11
+   -1.317806221963233e-12
+   -9.485241087407873e-12
+    8.303606756735972e-11
+   -7.361159682145734e-13
+   -1.311461787690749e-12
+   -2.009438267076375e-11
+    8.136729926334137e-11
+ 2.31e+10    
+    8.136456980292606e-11
+   -2.010035065132455e-11
+    8.302429874993025e-11
+   -1.342873687007732e-12
+   -9.487335641272806e-12
+    8.303137910005489e-11
+   -7.525694857678552e-13
+   -1.335950115808773e-12
+   -2.009930668411235e-11
+    8.135310322898497e-11
+ 2.36e+10    
+    8.135050719095906e-11
+   -2.010564038268102e-11
+     8.30199963478629e-11
+    -1.36774872909481e-12
+   -9.489929350270406e-12
+    8.302715349952053e-11
+   -7.686575468031275e-13
+   -1.360222471033413e-12
+   -2.010461379579943e-11
+    8.133889633576986e-11
+ 2.41e+10    
+    8.133642166061726e-11
+   -2.011132234820976e-11
+    8.301613581258418e-11
+   -1.392337698277091e-12
+    -9.49304208413969e-12
+    8.302337091291383e-11
+   -7.843808639250142e-13
+   -1.384190122857421e-12
+   -2.011031374335548e-11
+    8.132466381466218e-11
+ 2.46e+10    
+    8.132229669252783e-11
+   -2.011740802992165e-11
+    8.301269746560323e-11
+      -1.416527296012e-12
+   -9.496699023694961e-12
+    8.302001114320316e-11
+   -7.997472946902734e-13
+   -1.407747525772559e-12
+   -2.011641757002302e-11
+    8.131038998575461e-11
+ 2.51e+10    
+    8.130811464318113e-11
+   -2.012391086894215e-11
+    8.300966149118287e-11
+   -1.440179342035658e-12
+   -9.500932188736664e-12
+    8.301705358268055e-11
+   -8.147732976857663e-13
+   -1.430768165902883e-12
+   -2.012293798131119e-11
+    8.129605817104039e-11
+ 2.56e+10    
+     8.12938565402009e-11
+   -2.013084680629268e-11
+    8.300700793418539e-11
+   -1.463124313256179e-12
+   -9.505782298449282e-12
+    8.301447710556048e-11
+   -8.294857163307153e-13
+   -1.453099530393244e-12
+   -2.012988978043413e-11
+    8.128165056411195e-11
+ 2.61e+10    
+    8.127950181128496e-11
+   -2.013823494320108e-11
+    8.300471668534073e-11
+   -1.485153498189299e-12
+   -9.511301003262387e-12
+    8.301225991542311e-11
+   -8.439239291338606e-13
+   -1.474557123728082e-12
+   -2.013729039070217e-11
+    8.126714805453475e-11
+ 2.66e+10    
+    8.126502794366027e-11
+   -2.014609832689501e-11
+    8.300276745685149e-11
+   -1.506009709379113e-12
+   -9.517553498930436e-12
+    8.301037934486873e-11
+   -8.581423770728101e-13
+   -1.494917542313701e-12
+   -2.014516046542252e-11
+    8.125253000750037e-11
+ 2.71e+10    
+    8.125041007929438e-11
+   -2.015446484904743e-11
+    8.300113975284179e-11
+   -1.525376720856215e-12
+   -9.524621471949359e-12
+    8.300881160924797e-11
+   -8.722134175954665e-13
+    -1.51391079551489e-12
+   -2.015352457035408e-11
+    8.123777400571998e-11
+ 2.76e+10    
+    8.123562056804214e-11
+   -2.016336820691716e-11
+    8.299981284083186e-11
+   -1.542868039105406e-12
+   -9.532606206704472e-12
+    8.300753152635868e-11
+   -8.862303367375483e-13
+    -1.53121238556097e-12
+   -2.016241189522479e-11
+     8.12228555720833e-11
+ 2.81e+10    
+    8.122062853218994e-11
+   -2.017284881036178e-11
+    8.299876573269436e-11
+   -1.558016407809623e-12
+   -9.541631475551527e-12
+    8.300651223343004e-11
+    -9.00310143354964e-13
+   -1.546436210261176e-12
+   -2.017185690157039e-11
+    8.120774791148191e-11
+ 2.86e+10    
+    8.120539954863631e-11
+   -2.018295440690118e-11
+    8.299797718551034e-11
+   -1.570266761120202e-12
+   -9.551845489689358e-12
+    8.300572496642383e-11
+    -9.14595428870172e-13
+   -1.559130230016866e-12
+   -2.018189973539529e-11
+    8.119242174210748e-11
+ 2.91e+10    
+    8.118989563685675e-11
+   -2.019374002664002e-11
+    8.299742573395871e-11
+   -1.578977346909383e-12
+   -9.563420670086622e-12
+    8.300513902067853e-11
+    -9.29254061582976e-13
+   -1.568778132202077e-12
+   -2.019258611623662e-11
+     8.11768453336585e-11
+ 2.96e+10    
+    8.117407585438941e-11
+   -2.020526661632715e-11
+    8.299708976512501e-11
+   -1.583436472810831e-12
+   -9.576549295268954e-12
+    8.300472208794801e-11
+   -9.444747883657916e-13
+   -1.574811934616591e-12
+    -2.02039662583268e-11
+    8.116098493285237e-11
+ 3.01e+10    
+     8.11578979319309e-11
+   -2.021759746917934e-11
+    8.299694764505298e-11
+   -1.582905381691341e-12
+   -9.591432294926495e-12
+    8.300444125331297e-11
+   -9.604560362606735e-13
+   -1.576642350208459e-12
+   -2.021609220642072e-11
+    8.114480582772268e-11
+ 3.06e+10    
+    8.114132147333176e-11
+   -2.023079137775841e-11
+    8.299697790777578e-11
+   -1.576699776982401e-12
+   -9.608257913936312e-12
+    8.300426499788018e-11
+    -9.77384668509487e-13
+   -1.573715025855038e-12
+   -2.022901284728826e-11
+    8.112827435513798e-11
+ 3.11e+10    
+    8.112431318162261e-11
+   -2.024489158782093e-11
+    8.299715953461341e-11
+    -1.56432054819634e-12
+   -9.627167382056447e-12
+    8.300416650310178e-11
+   -9.954018599238076e-13
+   -1.565599865087177e-12
+   -2.024276593535858e-11
+    8.111136113610318e-11
+ 3.16e+10    
+    8.110685415845964e-11
+   -2.025991050017902e-11
+    8.299747240106715e-11
+   -1.545633696818665e-12
+   -9.648207214317184e-12
+    8.300412825176776e-11
+   -1.014555729740045e-12
+    -1.55211502243909e-12
+   -2.025736697997365e-11
+     8.10940456405743e-11
+ 3.21e+10    
+    8.108894837496011e-11
+   -2.027581202632972e-11
+    8.299789805586686e-11
+   -1.521076050343543e-12
+   -9.671273444028825e-12
+    8.300414724165085e-11
+   -1.034746002751844e-12
+   -1.533474188203918e-12
+   -2.027279602472028e-11
+    8.107632173908303e-11
+ 3.26e+10    
+    8.107062997903323e-11
+   -2.029249643546191e-11
+    8.299842106613804e-11
+   -1.491828739648848e-12
+   -9.696061764478075e-12
+    8.300423913332511e-11
+   -1.055674570521741e-12
+   -1.510425305269467e-12
+   -2.028898521623603e-11
+    8.105820316667554e-11
+ 3.31e+10    
+    8.105196581259978e-11
+    -2.03097951656542e-11
+    8.299903106014399e-11
+   -1.459870061247963e-12
+   -9.722045843688282e-12
+    8.300443884389842e-11
+   -1.076824033709392e-12
+   -1.484327290639313e-12
+   -2.030581200821096e-11
+    8.103972699843902e-11
+ 3.36e+10    
+    8.103304961537449e-11
+   -2.032748287524993e-11
+    8.299972514202182e-11
+   -1.427823457809589e-12
+   -9.748506840714479e-12
+    8.300479540973511e-11
+   -1.097487044702208e-12
+   -1.457103950780559e-12
+   -2.032310346159662e-11
+    8.102095283207988e-11
+ 3.41e+10    
+    8.101398698122253e-11
+   -2.034530876079028e-11
+    8.300050961134045e-11
+   -1.398580504264867e-12
+    -9.77462344963708e-12
+    8.300536106741007e-11
+    -1.11685566005973e-12
+   -1.431039035853837e-12
+   -2.034065476609217e-11
+    8.100195607178575e-11
+ 3.46e+10    
+     8.09948746303573e-11
+   -2.036303997510212e-11
+    8.300139947329771e-11
+   -1.374788067489091e-12
+   -9.799605246950411e-12
+    8.300617774393392e-11
+   -1.134153575257743e-12
+   -1.408436602345666e-12
+   -2.035825960906193e-11
+    8.098281577461017e-11
+ 3.51e+10    
+    8.097578116450507e-11
+   -2.038050245287567e-11
+    8.300241483601972e-11
+   -1.358375325819004e-12
+   -9.822827437752069e-12
+    8.300726621960551e-11
+   -1.148769658721328e-12
+   -1.391239812003592e-12
+   -2.037574389365052e-11
+    8.096360016352736e-11
+ 3.56e+10    
+    8.095673619524805e-11
+   -2.039760471346019e-11
+    8.300357494799783e-11
+   -1.350288551120809e-12
+    -9.84392091186168e-12
+    8.300862214000917e-11
+   -1.160347091301216e-12
+   -1.380732600692084e-12
+   -2.039299173815505e-11
+    8.094435444502989e-11
+ 3.61e+10    
+    8.093773049971999e-11
+   -2.041433866424238e-11
+    8.300489213997849e-11
+   -1.350498071630503e-12
+   -9.862792658615238e-12
+    8.301021940717468e-11
+    -1.16880341254882e-12
+   -1.377414978389803e-12
+   -2.040995593774288e-11
+    8.092509473258261e-11
+ 3.66e+10    
+    8.091872480262591e-11
+    -2.04307618908108e-11
+    8.300636801470989e-11
+   -1.358218468560441e-12
+   -9.879583154012754e-12
+    8.301201807114513e-11
+   -1.174288083944707e-12
+   -1.381064711426785e-12
+   -2.042665207242477e-11
+    8.090580911856578e-11
+ 3.71e+10    
+    8.089966216971806e-11
+    -2.04469716637588e-11
+    8.300799288412931e-11
+   -1.372218722417281e-12
+   -9.894588844124265e-12
+    8.301397284209026e-11
+   -1.177105491332072e-12
+   -1.390927134225851e-12
+    -2.04431415992441e-11
+      8.0886464094106e-11
+ 3.76e+10    
+    8.088047951258459e-11
+   -2.046308020798882e-11
+    8.300974785797742e-11
+   -1.391110920804338e-12
+   -9.908180563499325e-12
+    8.301603956127477e-11
+   -1.177633973259087e-12
+   -1.405947846576379e-12
+   -2.045951144659383e-11
+    8.086701317476688e-11
+ 3.81e+10    
+     8.08611158347087e-11
+   -2.047919653868251e-11
+    8.301160817983381e-11
+   -1.413558094156189e-12
+   -9.920738243044612e-12
+    8.301817882925735e-11
+   -1.176261046217293e-12
+   -1.424979322168874e-12
+   -2.047585606532487e-11
+    8.084740496215678e-11
+ 3.86e+10    
+    8.084151686107683e-11
+   -2.049541593294024e-11
+    8.301354651981765e-11
+   -1.438391518379869e-12
+   -9.932609022887484e-12
+    8.302035726310463e-11
+   -1.173341863095352e-12
+   -1.446927377958037e-12
+   -2.049226480003298e-11
+    8.082758912052651e-11
+ 3.91e+10    
+    8.082163680769471e-11
+   -2.051181562657518e-11
+    8.301553549804859e-11
+   -1.464655867735499e-12
+   -9.944086637109628e-12
+    8.302254728274255e-11
+   -1.169178773497832e-12
+   -1.470833983695904e-12
+   -2.050881480713412e-11
+    8.080751995299019e-11
+ 3.96e+10    
+    8.080143833642468e-11
+   -2.052845457717979e-11
+    8.301754925716875e-11
+   -1.491608241179742e-12
+   -9.955406027552912e-12
+    8.302472621870963e-11
+   -1.164015983755263e-12
+   -1.495909609199159e-12
+   -2.052556833270372e-11
+    8.078715798161763e-11
+ 4.01e+10    
+    8.078089158164881e-11
+   -2.054537538594076e-11
+    8.301956422325253e-11
+   -1.518693398615594e-12
+    -9.96674695071925e-12
+    8.302687525120284e-11
+   -1.158043128782465e-12
+   -1.521532768199648e-12
+   -2.054257280636002e-11
+    8.076647017425324e-11
+ 4.06e+10    
+    8.075997284438763e-11
+   -2.056260705520503e-11
+    8.302155930351667e-11
+   -1.545510366490942e-12
+   -9.978241800547649e-12
+    8.302897843811174e-11
+   -1.151403018065199e-12
+   -1.547232028594084e-12
+   -2.055986243066631e-11
+    8.074542940864323e-11
+ 4.11e+10    
+    8.073866328984836e-11
+   -2.058016781207575e-11
+    8.302351575487102e-11
+    -1.57177904020842e-12
+   -9.989984601964402e-12
+    8.303102192534552e-11
+   -1.144200537432905e-12
+   -1.572661134330748e-12
+   -2.057746035128473e-11
+     8.07240136025823e-11
+ 4.16e+10    
+    8.071694780404331e-11
+    -2.05980676253404e-11
+    8.302541689591382e-11
+   -1.597310825640322e-12
+   -1.000203952591541e-11
+    8.303299334784478e-11
+   -1.136511072688021e-12
+   -1.597573552414335e-12
+   -2.059538086818141e-11
+    8.070220477453586e-11
+ 4.21e+10    
+    8.069481405892505e-11
+   -2.061631028495704e-11
+     8.30272477713973e-11
+    -1.62198462819468e-12
+   -1.001444820376355e-11
+    8.303488139390358e-11
+   -1.128387740816323e-12
+   -1.621799599776395e-12
+   -2.061363141960393e-11
+    8.067998817394752e-11
+ 4.26e+10    
+    8.067225178110514e-11
+   -2.063489504088474e-11
+    8.302899482908076e-11
+   -1.645728087347987e-12
+   -1.002723565562633e-11
+    8.303667549695268e-11
+   -1.119867245955443e-12
+   -1.645227331235926e-12
+   -2.063221423946996e-11
+    8.065735153952041e-11
+ 4.31e+10    
+    8.064925219643951e-11
+   -2.065381785469508e-11
+    8.303064563635332e-11
+   -1.668503353664696e-12
+   -1.004041491550854e-11
+    8.303836562146193e-11
+   -1.110974443320509e-12
+   -1.667787289074731e-12
+    -2.06511276808834e-11
+    8.063428449772387e-11
+ 4.36e+10    
+    8.062580761669029e-11
+   -2.067307233470241e-11
+    8.303218864507903e-11
+   -1.690296541563244e-12
+   -1.005399054546204e-11
+    8.303994211611589e-11
+   -1.101725802224522e-12
+   -1.689440708802115e-12
+   -2.067036724141077e-11
+    8.061077809099578e-11
+ 4.41e+10    
+    8.060191113646368e-11
+   -2.069265042357371e-11
+    8.303361300328353e-11
+   -1.711110035424702e-12
+   -1.006796125436027e-11
+     8.30413956140995e-11
+   -1.092131982389574e-12
+   -1.710170599575142e-12
+   -2.068992634046598e-11
+    8.058682441611154e-11
+ 4.46e+10    
+    8.057755641342703e-11
+   -2.071254289778588e-11
+    8.303490840785741e-11
+   -1.730956951085754e-12
+    -1.00823218203382e-11
+    8.304271696589378e-11
+   -1.082199721113205e-12
+   -1.729975111152659e-12
+   -2.070979689960071e-11
+    8.056241635153398e-11
+ 4.51e+10    
+     8.05527375103462e-11
+   -2.073273972681365e-11
+     8.30360649912053e-11
+   -1.749857195342517e-12
+   -1.009706448452878e-11
+    8.304389719433277e-11
+   -1.071933197657773e-12
+   -1.748862666829885e-12
+   -2.072996977050729e-11
+    8.053754735435828e-11
+ 4.56e+10    
+    8.052744878241176e-11
+   -2.075323032922685e-11
+    8.303707323504345e-11
+    -1.76783469433342e-12
+   -1.011217995009208e-11
+    8.304492746474773e-11
+   -1.061335007728046e-12
+   -1.766848432997982e-12
+   -2.075043504774088e-11
+    8.051221131050522e-11
+ 4.61e+10    
+    8.050168479747133e-11
+   -2.077400375373822e-11
+    8.303792390528231e-11
+   -1.784915468567245e-12
+   -1.012765809005136e-11
+    8.304579906535337e-11
+   -1.050406850781843e-12
+    -1.78395178586394e-12
+   -2.077118229528588e-11
+    8.048640242499982e-11
+ 4.66e+10    
+    8.047544027992983e-11
+   -2.079504880601515e-11
+    8.303860800315085e-11
+   -1.801126316165536e-12
+   -1.014348844236073e-11
+    8.304650339441015e-11
+   -1.039150007786157e-12
+    -1.80019451400589e-12
+   -2.079220070952347e-11
+    8.046011514216585e-11
+ 4.71e+10    
+    8.044871007167411e-11
+   -2.081635413666113e-11
+    8.303911672856893e-11
+   -1.816493930055148e-12
+   -1.015966055060233e-11
+    8.304703195203708e-11
+   -1.027565667407576e-12
+   -1.815599559419428e-12
+   -2.081347923554187e-11
+    8.043334408786939e-11
+ 4.76e+10    
+    8.042148910507707e-11
+   -2.083790830143839e-11
+    8.303944145275689e-11
+   -1.831044322601925e-12
+   -1.017616419347291e-11
+    8.304737633493746e-11
+   -1.015655143346004e-12
+   -1.830190149765989e-12
+   -2.083500664947261e-11
+    8.040608402799409e-11
+ 4.81e+10    
+    8.039377238459005e-11
+   -2.085969980184381e-11
+    8.303957369773192e-11
+   -1.844802466612669e-12
+   -1.019298953461968e-11
+    8.304752823313695e-11
+   -1.003420013958009e-12
+   -1.843989213054307e-12
+   -2.085677161622588e-11
+    8.037832983873362e-11
+ 4.86e+10    
+    8.036555497439238e-11
+    -2.08817171118521e-11
+    8.303950512089096e-11
+   -1.857792087087504e-12
+     -1.0210127215767e-11
+    8.304747942792535e-11
+   -9.908622071292447e-13
+   -1.857018994806206e-12
+   -2.087876272952085e-11
+    8.035007648548992e-11
+ 4.91e+10    
+    8.033683199023443e-11
+   -2.090394869499138e-11
+    8.303922750340578e-11
+   -1.870035556974054e-12
+   -1.022756841000291e-11
+    8.304722179055124e-11
+   -9.779840467354769e-13
+   -1.869300819316487e-12
+   -2.090096853921696e-11
+    8.032131900797232e-11
+ 4.96e+10    
+    8.030759859425006e-11
+   -2.092638301477984e-11
+    8.303873274138479e-11
+   -1.881553863601994e-12
+   -1.024530484701611e-11
+    8.304674728138303e-11
+   -9.647882725785362e-13
+   -1.880854952670249e-12
+   -2.092337756966289e-11
+    8.029205250978098e-11
+ 5.01e+10    
+    8.027784999171506e-11
+   -2.094900854056532e-11
+    8.303801283906111e-11
+   -1.892366622026064e-12
+   -1.026332881921492e-11
+    8.304604794927091e-11
+   -9.512780425161986e-13
+    -1.89170053657988e-12
+   -2.094597833165372e-11
+    8.026227215115967e-11
+ 5.06e+10    
+    8.024758142918185e-11
+   -2.097181375036838e-11
+    8.303705990349922e-11
+   -1.902492118701423e-12
+   -1.028163317476843e-11
+    8.304511593097794e-11
+   -9.374569227039808e-13
+   -1.901855571003273e-12
+   -2.096875932997957e-11
+    8.023197314402543e-11
+ 5.11e+10    
+    8.021678819347781e-11
+   -2.099478713175491e-11
+    8.303586614034962e-11
+   -1.911947373677501e-12
+   -1.030021130212239e-11
+     8.30439434506598e-11
+    -9.23328870430518e-13
+   -1.911336929465014e-12
+   -2.099170906792717e-11
+    8.020115074858095e-11
+ 5.16e+10    
+    8.018546561125513e-11
+   -2.101791718146957e-11
+    8.303442385042105e-11
+   -1.920748213228699e-12
+   -1.031905710909079e-11
+    8.304252281921488e-11
+   -9.088982125849189e-13
+   -1.920160395738042e-12
+    -2.10148160496997e-11
+    8.016980027102076e-11
+ 5.21e+10    
+    8.015360904887057e-11
+    -2.10411924043805e-11
+     8.30327254267671e-11
+   -1.928909347315548e-12
+   -1.033816499876709e-11
+    8.304084643362383e-11
+   -8.941696218969997e-13
+   -1.928340713704483e-12
+   -2.103806878152836e-11
+     8.01379170619954e-11
+ 5.26e+10    
+    8.012121391242062e-11
+   -2.106460131205376e-11
+    8.303076335220531e-11
+   -1.936444448053191e-12
+   -1.035752984380243e-11
+    8.303890677610646e-11
+   -8.791480924568543e-13
+   -1.935891644748138e-12
+   -2.106145577190442e-11
+     8.01054965155544e-11
+ 5.31e+10    
+    8.008827564786457e-11
+   -2.108813242124078e-11
+    8.302853019706436e-11
+   -1.943366226728264e-12
+   -1.037714696012004e-11
+    8.303669641321639e-11
+   -8.638389155275468e-13
+   -1.942826028625562e-12
+   -2.108496553133503e-11
+    8.007253406842729e-11
+ 5.36e+10    
+    8.005478974111993e-11
+   -2.111177425239033e-11
+    8.302601861718618e-11
+   -1.949686507764836e-12
+   -1.039701208081322e-11
+    8.303420799482683e-11
+   -8.482476562704252e-13
+   -1.949155845146669e-12
+   -2.110858657185177e-11
+    8.003902519948657e-11
+ 5.41e+10    
+    8.002075171812913e-11
+   -2.113551532832422e-11
+     8.30232213519953e-11
+   -1.955416298672144e-12
+   -1.041712133063224e-11
+    8.303143425294967e-11
+   -8.323801318532692e-13
+   -1.954892274780961e-12
+   -2.113230740640679e-11
+     8.00049654292984e-11
+ 5.46e+10    
+    7.998615714484761e-11
+   -2.115934417308691e-11
+    8.302013122263878e-11
+   -1.960565855482192e-12
+   -1.043747120143081e-11
+    8.302836800053865e-11
+   -8.162423911558619e-13
+   -1.960045757021942e-12
+   -2.115611654833419e-11
+    7.997035031974335e-11
+ 5.51e+10    
+    7.995100162713445e-11
+    -2.11832493110569e-11
+    8.301674113024493e-11
+   -1.965144743444957e-12
+   -1.045805852871254e-11
+     8.30250021301136e-11
+    -7.99840696200697e-13
+   -1.964626045784885e-12
+   -2.118000251086601e-11
+    7.993517547362437e-11
+ 5.56e+10    
+    7.991528081057268e-11
+   -2.120721926627765e-11
+    8.301304405411867e-11
+   -1.969161892995524e-12
+   -1.047888046938529e-11
+    8.302132961238139e-11
+   -7.831815053257837e-13
+   -1.968642261409305e-12
+   -2.120395380681542e-11
+    7.989943653424946e-11
+ 5.61e+10    
+    7.987899038017537e-11
+   -2.123124256204006e-11
+    8.300903305001285e-11
+   -1.972625651114002e-12
+   -1.049993448069699e-11
+    8.301734349470775e-11
+   -7.662714581155497e-13
+   -1.972102939114653e-12
+    -2.12279589484006e-11
+    7.986312918498873e-11
+ 5.66e+10    
+    7.984212606003036e-11
+   -2.125530772070777e-11
+    8.300470124835623e-11
+   -1.975543828291491e-12
+   -1.052121830042025e-11
+    8.301303689959335e-11
+   -7.491173619646506e-13
+   -1.975016073841343e-12
+   -2.125200644725249e-11
+    7.982624914878257e-11
+ 5.71e+10    
+    7.980468361283048e-11
+   -2.127940326371837e-11
+     8.30000418524824e-11
+   -1.977923741387477e-12
+   -1.054272992815226e-11
+    8.300840302300441e-11
+   -7.317261802499768e-13
+   -1.977389161613425e-12
+   -2.127608481455525e-11
+    7.978879218758163e-11
+ 5.76e+10    
+    7.976665883937408e-11
+   -2.130351771185777e-11
+    8.299504813689976e-11
+   -1.979772252626125e-12
+   -1.056446760780153e-11
+    8.300343513277178e-11
+   -7.141050219309809e-13
+   -1.979229237498942e-12
+   -2.130018256141556e-11
+    7.975075410177969e-11
+ 5.81e+10    
+    7.972804757794911e-11
+   -2.132763958561841e-11
+    8.298971344543435e-11
+   -1.981095805061589e-12
+   -1.058642981102729e-11
+    8.299812656682053e-11
+   -6.962611325474652e-13
+   -1.980542910410959e-12
+   -2.132428819929664e-11
+    7.971213072954686e-11
+ 5.86e+10    
+    7.968884570371425e-11
+   -2.135175740581601e-11
+    8.298403118949158e-11
+   -1.981900454804976e-12
+   -1.060861522172759e-11
+    8.299247073145399e-11
+   -6.782018864082372e-13
+   -1.981336394912691e-12
+   -2.134839024067935e-11
+    7.967291794617578e-11
+ 5.91e+10    
+    7.964904912798836e-11
+   -2.137585969428492e-11
+    8.297799484621091e-11
+   -1.982191900276023e-12
+    -1.06310227213911e-11
+    8.298646109956988e-11
+   -6.599347799216414e-13
+   -1.981615540302999e-12
+   -2.137247719977848e-11
+     7.96331116633401e-11
+ 5.96e+10    
+    7.960865379752678e-11
+   -2.139993497472922e-11
+    8.297159795666077e-11
+    -1.98197550880325e-12
+   -1.065365137529893e-11
+    8.298009120887257e-11
+      -6.414674258907e-13
+   -1.981385857123517e-12
+   -2.139653759343499e-11
+    7.959270782836869e-11
+ 6.01e+10    
+    7.956765569374839e-11
+   -2.142397177367958e-11
+    8.296483412401163e-11
+   -1.981256340734377e-12
+   -1.067650041947463e-11
+    8.297335466002657e-11
+   -6.228075487294243e-13
+    -1.98065254138542e-12
+   -2.142055994204494e-11
+    7.955170242344262e-11
+ 6.06e+10    
+    7.952605083195576e-11
+   -2.144795862154435e-11
+    8.295769701167397e-11
+   -1.980039171423387e-12
+   -1.069956924834244e-11
+    8.296624511485296e-11
+   -6.039629803996969e-13
+   -1.979420496649602e-12
+   -2.144453277064279e-11
+    7.951009146481812e-11
+ 6.11e+10    
+    7.948383526051396e-11
+   -2.147188405375612e-11
+    8.295018034151037e-11
+   -1.978328511171426e-12
+   -1.072285740303402e-11
+    8.295875629448132e-11
+   -5.849416570532466e-13
+   -1.977694354216526e-12
+   -2.146844461002408e-11
+    7.946787100201235e-11
+ 6.16e+10    
+    7.944100506003393e-11
+   -2.149573661196319e-11
+    8.294227789196923e-11
+   -1.976128623446117e-12
+   -1.074636456027698e-11
+     8.29508819775084e-11
+   -5.657516162336375e-13
+   -1.975478491550251e-12
+   -2.149228399794267e-11
+     7.94250371169706e-11
+ 6.21e+10    
+    7.939755634254547e-11
+   -2.151950484532195e-11
+    8.293398349624785e-11
+   -1.973443541501353e-12
+   -1.077009052176007e-11
+    8.294261599814021e-11
+   -5.464009945085313e-13
+   -1.972777049178563e-12
+   -2.151603948037555e-11
+    7.938158592324665e-11
+ 6.26e+10    
+    7.935348525066071e-11
+   -2.154317731180085e-11
+    8.292529104048604e-11
+   -1.970277083544901e-12
+    -1.07940352040688e-11
+    8.293395224436668e-11
+   -5.268980255758856e-13
+   -1.969593946133357e-12
+   -2.153969961282898e-11
+    7.933751356517264e-11
+ 6.31e+10    
+    7.930878795674941e-11
+   -2.156674257955566e-11
+    8.291619446192389e-11
+   -1.966632866669583e-12
+   -1.081819862900471e-11
+    8.292488465611003e-11
+   -5.072510385926687e-13
+   -1.965932894175086e-12
+   -2.156325296168956e-11
+    7.929281621703026e-11
+ 6.36e+10    
+    7.926346066212358e-11
+   -2.159018922833957e-11
+    8.290668774711515e-11
+   -1.962514319651047e-12
+   -1.084258091427732e-11
+    8.291540722341005e-11
+     -4.8746845677716e-13
+   -1.961797410862579e-12
+   -2.158668810561297e-11
+    7.924749008223809e-11
+ 6.41e+10    
+    7.921749959621542e-11
+    -2.16135058509067e-11
+    8.289676493008608e-11
+   -1.957924694724615e-12
+   -1.086718226461004e-11
+    8.290551398459168e-11
+   -4.675587961722922e-13
+   -1.957190831613852e-12
+    -2.16099936369476e-11
+    7.920153139254138e-11
+ 6.46e+10    
+    7.917090101579594e-11
+   -2.163668105451264e-11
+    8.288642009061209e-11
+   -1.952867078473786e-12
+   -1.089200296316084e-11
+    8.289519902447277e-11
+   -4.475306644990697e-13
+   -1.952116320866244e-12
+    -2.16331581631703e-11
+    7.915493640722646e-11
+ 6.51e+10    
+     7.91236612041899e-11
+   -2.165970346234538e-11
+    8.287564735237255e-11
+   -1.947344401961058e-12
+   -1.091704336317295e-11
+    8.288445647256419e-11
+   -4.273927600359878e-13
+   -1.946576882475321e-12
+   -2.165617030834401e-11
+    7.910770141234537e-11
+ 6.56e+10    
+    7.907577647053858e-11
+   -2.168256171506042e-11
+    8.286444088127633e-11
+   -1.941359450104183e-12
+    -1.09423038800065e-11
+    8.287328050131727e-11
+   -4.071538705299851e-13
+   -1.940575369329874e-12
+   -2.167901871460945e-11
+    7.905982271996283e-11
+ 6.61e+10    
+      7.9027243149052e-11
+   -2.170524447225283e-11
+    8.285279488365428e-11
+   -1.934914870497496e-12
+   -1.096778498328463e-11
+    8.286166532434835e-11
+   -3.868228719960109e-13
+   -1.934114492422435e-12
+   -2.170169204367409e-11
+    7.901129666744046e-11
+ 6.66e+10    
+    7.897805759832827e-11
+   -2.172774041399608e-11
+    8.284070360461237e-11
+   -1.928013181666518e-12
+   -1.099348718936171e-11
+    8.284960519472155e-11
+   -3.664087274420476e-13
+   -1.927196829326191e-12
+   -2.172417897831227e-11
+    7.896211961673181e-11
+ 6.71e+10    
+    7.892821620066948e-11
+   -2.175003824234812e-11
+    8.282816132628574e-11
+   -1.920656780861474e-12
+   -1.101941105392487e-11
+    8.283709440323491e-11
+    -3.45920485431051e-13
+   -1.919824832199386e-12
+   -2.174646822386978e-11
+    7.891228795371351e-11
+ 6.76e+10    
+    7.887771536145443e-11
+   -2.177212668288309e-11
+    8.281516236620354e-11
+   -1.912847951435714e-12
+   -1.104555716479359e-11
+    8.282412727672573e-11
+   -3.253672784936595e-13
+   -1.912000835376797e-12
+   -2.176854850977959e-11
+    7.886179808755168e-11
+ 6.81e+10    
+    7.882655150853409e-11
+   -2.179399448622234e-11
+    8.280170107563973e-11
+   -1.904588869881409e-12
+   -1.107192613490352e-11
+    8.281069817643359e-11
+   -3.047583212871977e-13
+   -1.903727062579257e-12
+   -2.179040859109733e-11
+    7.881064645011251e-11
+ 6.86e+10    
+    7.877472109167443e-11
+   -2.181563042955639e-11
+    8.278777183795768e-11
+   -1.895881612579383e-12
+   -1.109851859535621e-11
+    8.279680149631521e-11
+   -2.841029085482704e-13
+   -1.895005633844748e-12
+   -2.181203724999178e-11
+     7.87588294953817e-11
+ 6.91e+10    
+    7.872222058202195e-11
+   -2.183702331818141e-11
+    8.277336906707056e-11
+   -1.886728162228636e-12
+   -1.112533518872146e-11
+     8.27824316614831e-11
+   -2.634104128035697e-13
+   -1.885838572135331e-12
+    -2.18334232972877e-11
+    7.870634369895378e-11
+ 6.96e+10    
+     7.86690464716364e-11
+   -2.185816198702177e-11
+    8.275848720581663e-11
+   -1.877130414139373e-12
+   -1.115237656232721e-11
+    8.276758312658024e-11
+   -2.426902817582273e-13
+   -1.876227809768831e-12
+   -2.185455557397523e-11
+    7.865318555754791e-11
+ 7.01e+10    
+    7.861519527304239e-11
+   -2.187903530216227e-11
+    8.274312072446335e-11
+   -1.867090182276262e-12
+   -1.117964336176503e-11
+    8.275225037424084e-11
+   -2.219520354205181e-13
+    -1.86617519461771e-12
+   -2.187542295272248e-11
+    7.859935158856488e-11
+ 7.06e+10    
+    7.856066351883906e-11
+   -2.189963216235671e-11
+     8.27272641191525e-11
+   -1.856609205188779e-12
+   -1.120713622442545e-11
+    8.273642791354858e-11
+   -2.012052629216427e-13
+   -1.855682496174019e-12
+   -2.189601433940265e-11
+    7.854483832970091e-11
+ 7.11e+10    
+    7.850544776135199e-11
+    -2.19199415005535e-11
+    8.271091191042271e-11
+   -1.845689151802264e-12
+   -1.123485577313002e-11
+    8.272011027853256e-11
+   -1.804596190084599e-13
+    -1.84475141146155e-12
+   -2.191631867458359e-11
+    7.848964233859189e-11
+ 7.16e+10    
+    7.844954457234443e-11
+   -2.193995228540766e-11
+    8.269405864175341e-11
+   -1.834331627124074e-12
+    -1.12628026098511e-11
+    8.270329202668903e-11
+   -1.597248202138912e-13
+   -1.833383570864255e-12
+   -2.193632493505162e-11
+    7.843376019251583e-11
+ 7.21e+10    
+    7.839295054275147e-11
+   -2.195965352277955e-11
+    8.267669887812496e-11
+   -1.822538177849727e-12
+   -1.129097730952218e-11
+    8.268596773752912e-11
+   -1.390106407322622e-13
+   -1.821580543842295e-12
+   -2.195602213530007e-11
+    7.837718848815021e-11
+ 7.26e+10    
+    7.833566228249637e-11
+   -2.197903425723356e-11
+    8.265882720457876e-11
+   -1.810310297952237e-12
+   -1.131938041384854e-11
+    8.266813201115649e-11
+   -1.183269079225882e-13
+   -1.809343844617499e-12
+   -2.197539932902037e-11
+    7.831992384135689e-11
+ 7.31e+10    
+     7.82776764203389e-11
+      -2.199808357354e-11
+    8.264043822489656e-11
+   -1.797649434192208e-12
+     -1.1348012425261e-11
+    8.264977946686402e-11
+   -9.768349752264172e-14
+   -1.796674937795123e-12
+   -2.199444561059177e-11
+    7.826196288704644e-11
+ 7.36e+10    
+    7.821898960377864e-11
+   -2.201679059814431e-11
+    8.262152656019238e-11
+    -1.78455699164649e-12
+   -1.137687380083587e-11
+    8.263090474177509e-11
+   -7.709032851980657e-14
+   -1.783575243969379e-12
+   -2.201315011656113e-11
+    7.820330227907943e-11
+ 7.41e+10    
+    7.815959849902282e-11
+   -2.203514450065522e-11
+    8.260208684759343e-11
+   -1.771034339188606e-12
+   -1.140596494633202e-11
+    8.261150248948919e-11
+   -5.655735771772883e-14
+   -1.770046145289695e-12
+   -2.203150202710649e-11
+    7.814393869021444e-11
+ 7.46e+10    
+    7.809949979098362e-11
+   -2.205313449529066e-11
+    8.258211373894096e-11
+   -1.757082815010913e-12
+   -1.143528621020592e-11
+    8.259156737876151e-11
+   -3.609457399283893e-14
+   -1.756088991064072e-12
+   -2.204949056750251e-11
+    7.808386881212969e-11
+ 7.51e+10    
+    7.803869018336645e-11
+   -2.207074984236216e-11
+    8.256160189952312e-11
+    -1.74270373211929e-12
+   -1.146483787774961e-11
+    8.257109409223193e-11
+   -1.571199223026956e-14
+   -1.741705103340543e-12
+   -2.206710500956888e-11
+    7.802308935548455e-11
+ 7.56e+10    
+    7.797716639877717e-11
+   -2.208797984969482e-11
+    8.254054600678801e-11
+    -1.72789838388857e-12
+   -1.149462016516211e-11
+     8.25500773251217e-11
+    4.580352996423611e-15
+   -1.726895782508771e-12
+   -2.208433467311193e-11
+     7.79615970500343e-11
+ 7.61e+10    
+    7.791492517890937e-11
+   -2.210481387407737e-11
+    8.251894074915592e-11
+   -1.712668049615241e-12
+   -1.152463321374626e-11
+    8.252851178403982e-11
+    2.477241406929986e-14
+   -1.711662312937572e-12
+   -2.210116892736878e-11
+    7.789938864482405e-11
+ 7.66e+10    
+    7.785196328477481e-11
+    -2.21212413226796e-11
+    8.249678082476645e-11
+   -1.697014000128422e-12
+   -1.155487708407182e-11
+    8.250639218571856e-11
+    4.485413720914762e-14
+   -1.696005968645493e-12
+   -2.211759719239367e-11
+    7.783646090838821e-11
+ 7.71e+10    
+    7.778827749699484e-11
+   -2.213725165446804e-11
+    8.247406094034527e-11
+   -1.680937503413329e-12
+   -1.158535175022803e-11
+    8.248371325583926e-11
+    6.481546960848368e-14
+   -1.679928018977589e-12
+   -2.213360894049944e-11
+    7.777281062906889e-11
+ 7.76e+10    
+    7.772386461613951e-11
+   -2.215283438159976e-11
+    8.245077581000781e-11
+   -1.664439830317806e-12
+   -1.161605709401984e-11
+    8.246046972786335e-11
+     8.46463668503814e-14
+   -1.663429734377765e-12
+   -2.214919369763042e-11
+    7.770843461533265e-11
+ 7.81e+10    
+    7.765872146313668e-11
+   -2.216797907081149e-11
+    8.242692015412238e-11
+   -1.647522260246038e-12
+   -1.164699289929381e-11
+    8.243665634187996e-11
+     1.04336800481038e-13
+   -1.646512392131117e-12
+   -2.216434104476174e-11
+    7.764332969618898e-11
+ 7.86e+10    
+    7.759284487971809e-11
+   -2.218267534479688e-11
+    8.240248869822637e-11
+   -1.630186086958645e-12
+   -1.167815884620953e-11
+    8.241226784346633e-11
+    1.238767658715834e-13
+   -1.629177282225154e-12
+   -2.217904061924509e-11
+    7.757749272162119e-11
+ 7.91e+10    
+     7.75262317289332e-11
+   -2.219691288354924e-11
+    8.237747617187811e-11
+   -1.612432624397361e-12
+   -1.170955450556244e-11
+    8.238729898258911e-11
+     1.43256290215568e-13
+   -1.611425713203798e-12
+     -2.2193282116177e-11
+    7.751092056310075e-11
+ 7.96e+10    
+    7.745887889571147e-11
+    -2.22106814257243e-11
+    8.235187730762346e-11
+    -1.59426321253981e-12
+    -1.17411793331543e-11
+    8.236174451252143e-11
+    1.624654407474286e-13
+    -1.59325901810014e-12
+   -2.220705528973767e-11
+    7.744361011415198e-11
+ 8.01e+10    
+    7.739078328747331e-11
+   -2.222397076994507e-11
+    8.232568683990263e-11
+   -1.575679223330413e-12
+   -1.177303266415842e-11
+    8.233559918874306e-11
+    1.814943330837473e-13
+   -1.574678560390716e-12
+   -2.222034995449515e-11
+    7.737555829094794e-11
+ 8.06e+10    
+    7.732194183479843e-11
+   -2.223677077613198e-11
+     8.22988995040338e-11
+   -1.556682066654957e-12
+   -1.180511370752101e-11
+    8.230885776791625e-11
+    2.003331397664477e-13
+   -1.555685740027694e-12
+   -2.223315598673595e-11
+     7.73067620329892e-11
+ 8.11e+10    
+    7.725235149214537e-11
+   -2.224907136678412e-11
+    8.227151003517835e-11
+   -1.537273196341111e-12
+   -1.183742154042433e-11
+    8.228151500685597e-11
+    2.189720988666748e-13
+   -1.536281999484024e-12
+   -2.224546332573114e-11
+    7.723721830380549e-11
+ 8.16e+10    
+    7.718200923861977e-11
+   -2.226086252825969e-11
+    8.224351316732708e-11
+   -1.517454116226164e-12
+   -1.186995510271123e-11
+    8.225356566147978e-11
+    2.374015227713678e-13
+   -1.516468829860468e-12
+   -2.225726197501676e-11
+    7.716692409172395e-11
+ 8.21e+10    
+    7.711091207878517e-11
+   -2.227213431203533e-11
+    8.221490363231925e-11
+   -1.497226386264514e-12
+   -1.190271319139413e-11
+    8.222500448582968e-11
+    2.556118070294431e-13
+   -1.496247777040162e-12
+   -2.226854200365037e-11
+    7.709587641068659e-11
+ 8.26e+10    
+    7.703905704353047e-11
+   -2.228287683594201e-11
+    8.218567615884941e-11
+   -1.476591628649697e-12
+   -1.193569445519083e-11
+    8.219582623106718e-11
+    2.735934392787766e-13
+   -1.475620447844955e-12
+   -2.227929354743047e-11
+    7.702407230109297e-11
+ 8.31e+10    
+    7.696644119097867e-11
+   -2.229308028538957e-11
+    8.215582547151909e-11
+   -1.455551533996617e-12
+    -1.19688973890672e-11
+    8.216602564451856e-11
+    2.913370082561689e-13
+   -1.454588516283523e-12
+   -2.228950681012769e-11
+     7.69515088307253e-11
+ 8.36e+10    
+    7.689306160743464e-11
+    -2.23027349145646e-11
+    8.212534628988468e-11
+   -1.434107867544741e-12
+    -1.20023203288541e-11
+    8.213559746869541e-11
+    3.088332128541407e-13
+   -1.433153729769782e-12
+   -2.229917206466232e-11
+    7.687818309567811e-11
+ 8.41e+10    
+    7.681891540839049e-11
+   -2.231183104761802e-11
+    8.209423332752124e-11
+   -1.412262475396028e-12
+   -1.203596144586545e-11
+    8.210453644035927e-11
+    3.260728712097225e-13
+    -1.41131791541527e-12
+   -2.230827965428981e-11
+    7.680409222136107e-11
+ 8.46e+10    
+    7.674399973954985e-11
+   -2.232035907981209e-11
+    8.206248129107959e-11
+   -1.390017290761933e-12
+   -1.206981874158684e-11
+    8.207283728958885e-11
+    3.430469298133797e-13
+   -1.389082986319527e-12
+   -2.231681999374945e-11
+    7.672923336352747e-11
+ 8.51e+10    
+     7.66683117779149e-11
+   -2.232830947867373e-11
+    8.203008487940282e-11
+   -1.367374340245156e-12
+   -1.210389004238393e-11
+    8.204049473883915e-11
+    3.597464726346039e-13
+   -1.366450947889391e-12
+   -2.232478357039172e-11
+    7.665360370934082e-11
+ 8.56e+10    
+    7.659184873289102e-11
+    -2.23356727851067e-11
+    8.199703878260641e-11
+   -1.344335750110045e-12
+   -1.213817299430319e-11
+    8.200750350204688e-11
+    3.761627302203325e-13
+   -1.343423904154388e-12
+   -2.233216094529067e-11
+    7.657720047848795e-11
+ 8.61e+10    
+    7.651460784744475e-11
+   -2.234243961449358e-11
+    8.196333768120395e-11
+   -1.320903752583009e-12
+   -1.217266505787267e-11
+    8.197385828374267e-11
+    3.922870887935582e-13
+   -1.320004064112112e-12
+    -2.23389427543457e-11
+    7.650002092432485e-11
+ 8.66e+10    
+    7.643658639927088e-11
+   -2.234860065775721e-11
+    8.192897624520369e-11
+   -1.297080692151155e-12
+   -1.220736350297814e-11
+    8.193955377811494e-11
+    4.081110993181338e-13
+   -1.296193748061663e-12
+   -2.234511970931161e-11
+    7.642206233503765e-11
+ 8.71e+10    
+    7.635778170202209e-11
+   -2.235414668242606e-11
+     8.18939491332678e-11
+   -1.272869031846834e-12
+   -1.224226540381129e-11
+    8.190458466817806e-11
+    4.236264864894908e-13
+   -1.271995393937191e-12
+   -2.235068259887998e-11
+    7.634332203487391e-11
+ 8.76e+10    
+    7.627819110654542e-11
+   -2.235906853366917e-11
+    8.185825099184667e-11
+   -1.248271359521388e-12
+   -1.227736763387706e-11
+    8.186894562489557e-11
+     4.38825157715288e-13
+   -1.247411563626173e-12
+   -2.235562228968243e-11
+    7.626379738536301e-11
+ 8.81e+10    
+    7.619781200215461e-11
+   -2.236335713529712e-11
+    8.182187645433869e-11
+   -1.223290394099795e-12
+   -1.231266686105868e-11
+    8.183263130630686e-11
+    4.536992119577651e-13
+   -1.222444949265892e-12
+   -2.235992972728723e-11
+    7.618348578658643e-11
+ 8.86e+10    
+    7.611664181792207e-11
+   -2.236700349074025e-11
+    8.178482014022516e-11
+   -1.197928991843569e-12
+    -1.23481595427431e-11
+    8.179563635668521e-11
+      4.6824094858415e-13
+   -1.197098379550099e-12
+   -2.236359593717273e-11
+     7.61023846784693e-11
+ 8.91e+10    
+    7.603467802401017e-11
+   -2.236999868403491e-11
+    8.174707665429331e-11
+    -1.17219015253461e-12
+   -1.238384192106973e-11
+    8.175795540571927e-11
+    4.824428760465828e-13
+   -1.171374825951094e-12
+   -2.236661202569086e-11
+    7.602049154209365e-11
+ 8.96e+10    
+    7.595191813300431e-11
+   -2.237233388075033e-11
+    8.170864058579404e-11
+   -1.146077025639875e-12
+   -1.241971001821917e-11
+    8.171958306766908e-11
+    4.962977204781575e-13
+   -1.145277408948416e-12
+   -2.236896918098624e-11
+    7.593780390103385e-11
+ 9.01e+10    
+    7.586835970127832e-11
+   -2.237400032891427e-11
+    8.166950650765665e-11
+   -1.119592916450679e-12
+   -1.245575963181079e-11
+    8.168051394056269e-11
+     5.09798434219564e-13
+   -1.118809404195339e-12
+   -2.237065867390818e-11
+    7.585431932270921e-11
+ 9.06e+10    
+    7.578400033037409e-11
+   -2.237498935991158e-11
+    8.162966897568221e-11
+     -1.0927412921422e-12
+   -1.249198633037642e-11
+    8.164074260540582e-11
+    5.229382041635935e-13
+   -1.091974248625208e-12
+   -2.237167185889584e-11
+    7.577003541976145e-11
+ 9.11e+10    
+     7.56988376683948e-11
+   -2.237529238936851e-11
+    8.158912252780417e-11
+   -1.065525787783289e-12
+   -1.252838544896052e-11
+    8.160026362537249e-11
+    5.357104600154354e-13
+   -1.064775546527567e-12
+   -2.237200017483808e-11
+    7.568494985143057e-11
+ 9.16e+10    
+    7.561286941141644e-11
+   -2.237490091799913e-11
+    8.154786168330152e-11
+   -1.037950212277909e-12
+   -1.256495208480665e-11
+    8.155907154507098e-11
+    5.481088823826176e-13
+    -1.03721707550871e-12
+   -2.237163514592789e-11
+    7.559906032497171e-11
+ 9.21e+10    
+    7.552609330490575e-11
+    -2.23738065324578e-11
+    8.150588094206783e-11
+   -1.010018554226812e-12
+   -1.260168109315043e-11
+    8.151716088973977e-11
+    5.601274107234247e-13
+   -1.009302792421438e-12
+   -2.237056838247121e-11
+    7.551236459705373e-11
+ 9.26e+10    
+    7.543850714514852e-11
+   -2.237200090613692e-11
+    8.146317478386311e-11
+   -9.817349877167738e-13
+   -1.263856708313801e-11
+    8.147452616454758e-11
+    5.717602511676234e-13
+    -9.81036839192704e-13
+   -2.236879158168917e-11
+    7.542486047518251e-11
+ 9.31e+10    
+    7.535010878069902e-11
+   -2.236947579999551e-11
+    8.141973766766736e-11
+   -9.531038779896968e-13
+   -1.267560441390328e-11
+     8.14311618538654e-11
+     5.83001884106576e-13
+   -9.524235485387308e-13
+   -2.236629652851777e-11
+    7.533654581914031e-11
+ 9.36e+10    
+    7.526089611380682e-11
+   -2.236622306331203e-11
+    8.137556403091565e-11
+   -9.241297870338721e-13
+   -1.271278719070138e-11
+    8.138706242054346e-11
+    5.938470716883831e-13
+   -9.234674496210223e-13
+   -2.236307509634691e-11
+     7.52474185424074e-11
+ 9.41e+10    
+    7.517086710188333e-11
+   -2.236223463447569e-11
+    8.133064828889428e-11
+   -8.948174790638592e-13
+   -1.275010926124085e-11
+     8.13422223052483e-11
+    6.042908650719896e-13
+   -8.941732735493599e-13
+   -2.235911924778433e-11
+    7.515747661360964e-11
+ 9.46e+10    
+    7.508001975894445e-11
+   -2.235750254171342e-11
+     8.12849848340661e-11
+    -8.65171925862296e-13
+   -1.278756421215814e-11
+    8.129663592580255e-11
+    6.143286115377711e-13
+   -8.645459587925189e-13
+   -2.235442103538301e-11
+    7.506671805796004e-11
+ 9.51e+10    
+    7.498835215706593e-11
+   -2.235201890383827e-11
+    8.123856803546463e-11
+   -8.351983120096334e-13
+   -1.282514536560901e-11
+    8.125029767655904e-11
+    6.239559613567027e-13
+   -8.345906564485645e-13
+   -2.234897260235264e-11
+    7.497514095869829e-11
+ 9.56e+10    
+    7.489586242783655e-11
+   -2.234577593096557e-11
+    8.119139223810171e-11
+   -8.049020399724166e-13
+    -1.28628457760553e-11
+     8.12032019277862e-11
+    6.331688745149852e-13
+   -8.043127353774442e-13
+   -2.234276618326355e-11
+    7.488274345853684e-11
+ 9.61e+10    
+    7.480254876381323e-11
+   -2.233876592522275e-11
+    8.114345176242093e-11
+   -7.742887350437728e-13
+   -1.290065822719899e-11
+    8.115534302508456e-11
+    6.419636271847996e-13
+   -7.737177872030811e-13
+   -2.233579410472274e-11
+    7.478952376109652e-11
+ 9.66e+10    
+    7.470840941996782e-11
+   -2.233098128145281e-11
+    8.109474090377234e-11
+   -7.433642501139511e-13
+   -1.293857522911787e-11
+    8.110671528889508e-11
+    6.503368179959405e-13
+   -7.428116311256986e-13
+   -2.232804878607381e-11
+    7.469548013235087e-11
+ 9.71e+10    
+    7.461344271513401e-11
+   -2.232241448789531e-11
+    8.104525393192085e-11
+   -7.121346703039871e-13
+   -1.297658901554842e-11
+    8.105731301393191e-11
+    6.582853740961735e-13
+   -7.116003186028013e-13
+   -2.231952274004813e-11
+    7.460061090205691e-11
+ 9.76e+10    
+      7.4517647033446e-11
+   -2.231305812687655e-11
+    8.099498509059425e-11
+   -6.806063174091311e-13
+   -1.301469154138209e-11
+    8.100713046875217e-11
+    6.658065569759803e-13
+   -6.800901378381967e-13
+   -2.231020857341755e-11
+    7.450491446517619e-11
+ 9.81e+10    
+    7.442102082577147e-11
+   -2.230290487548033e-11
+    8.094392859709849e-11
+   -6.487857541325855e-13
+   -1.305287448038034e-11
+    8.095616189533086e-11
+    6.728979680509305e-13
+   -6.482876180759671e-13
+   -2.230009898766693e-11
+    7.440838928330754e-11
+ 9.86e+10    
+    7.432356261114593e-11
+   -2.229194750622788e-11
+    8.089207864193894e-11
+   -6.166797881735026e-13
+   -1.309112922305547e-11
+    8.090440150867498e-11
+    6.795575540219643e-13
+    -6.16199533720877e-13
+     -2.2289186779626e-11
+    7.431103388608647e-11
+ 9.91e+10    
+    7.422527097818468e-11
+   -2.228017888774436e-11
+    8.083942938852786e-11
+   -5.842954760596123e-13
+   -1.312944687481432e-11
+    8.085184349650097e-11
+     6.85783611973662e-13
+   -5.838329082382115e-13
+    -2.22774648421259e-11
+    7.421284687260901e-11
+ 9.96e+10    
+    7.412614458649708e-11
+   -2.226759198543393e-11
+    8.078597497292791e-11
+   -5.516401268133042e-13
+   -1.316781825428493e-11
+    8.079848201896898e-11
+    6.915747942313949e-13
+   -5.511950178398547e-13
+   -2.226492616464856e-11
+     7.41138269128122e-11
+ 1.001e+11   
+    7.402618216808903e-11
+   -2.225417986215385e-11
+    8.073170950365465e-11
+    -5.18721305351341e-13
+   -1.320623389192016e-11
+    8.074431120843484e-11
+    6.969301129643589e-13
+   -5.182933949601504e-13
+   -2.225156383395515e-11
+    7.401397274886685e-11
+ 1.006e+11   
+    7.392538252875563e-11
+   -2.223993567889608e-11
+     8.06766270615361e-11
+     -4.8554683568032e-13
+   -1.324468402880107e-11
+    8.068932516933416e-11
+    7.018489445033228e-13
+   -4.851358314746503e-13
+   -2.223737103476307e-11
+    7.391328319655392e-11
+ 1.011e+11   
+    7.382374454945887e-11
+   -2.222485269546928e-11
+    8.062072169966937e-11
+   -4.521248038279852e-13
+   -1.328315861573477e-11
+    8.063351797806919e-11
+    7.063310334118453e-13
+   -4.517303816916807e-13
+   -2.222234105039348e-11
+    7.381175714663645e-11
+ 1.016e+11   
+    7.372126718771019e-11
+    -2.22089242712036e-11
+    8.056398744339878e-11
+   -4.184635605436082e-13
+   -1.332164731257385e-11
+     8.05768836829999e-11
+    7.103764962678501e-13
+   -4.180853650790804e-13
+   -2.220646726344555e-11
+    7.370939356620932e-11
+ 1.021e+11   
+    7.361794947892195e-11
+   -2.219214386565976e-11
+     8.05064182904162e-11
+   -3.845717237019001e-13
+   -1.336013948784163e-11
+    8.051941630449076e-11
+    7.139858251668948e-13
+   -3.842093687342741e-13
+   -2.218974315647213e-11
+    7.360619150004601e-11
+ 1.026e+11   
+    7.351379053777248e-11
+   -2.217450503935214e-11
+      8.0448008210924e-11
+   -3.504581804714653e-13
+   -1.339862421861409e-11
+    8.046110983506209e-11
+      7.1715989094282e-13
+   -3.501112495773231e-13
+    -2.21721623126806e-11
+    7.350215007193776e-11
+ 1.031e+11   
+    7.340878955953354e-11
+   -2.215600145449496e-11
+    8.038875114787504e-11
+    -3.16132089166905e-13
+   -1.343709029068755e-11
+    8.040195823961916e-11
+    7.198999460760161e-13
+   -3.158001362567921e-13
+   -2.215371841664923e-11
+    7.339726848601503e-11
+ 1.036e+11   
+    7.330294582141441e-11
+   -2.213662687576335e-11
+    8.032864101732841e-11
+   -2.816028808385679e-13
+   -1.347552619905237e-11
+    8.034195545574055e-11
+    7.222076273315056e-13
+   -2.812854307719599e-13
+   -2.213440525505562e-11
+    7.329154602806355e-11
+ 1.041e+11   
+    7.319625868387752e-11
+   -2.211637517108222e-11
+    8.026767170886035e-11
+   -2.468802605481919e-13
+   -1.351392014865615e-11
+    8.028109539410475e-11
+    7.240849580688323e-13
+   -2.465768097840914e-13
+   -2.211421671743123e-11
+    7.318498206682196e-11
+ 1.046e+11   
+    7.308872759195333e-11
+   -2.209524031244253e-11
+     8.02058370861359e-11
+   -2.119742083109723e-13
+   -1.355226005550827e-11
+    8.021937193901203e-11
+    7.255343502308976e-13
+   -2.116842256128909e-13
+   -2.209314679695848e-11
+    7.307757605528987e-11
+ 1.051e+11   
+    7.298035207654685e-11
+   -2.207321637674374e-11
+    8.014313098753185e-11
+   -1.768949797684572e-13
+   -1.359053354806529e-11
+    8.015677894898486e-11
+    7.265586060595285e-13
+   -1.766179069340662e-13
+   -2.207118959126409e-11
+    7.296932753199609e-11
+ 1.056e+11   
+    7.287113175572881e-11
+   -2.205029754666629e-11
+    8.007954722691393e-11
+   -1.416531064952647e-13
+   -1.362872796897708e-11
+    8.009331025749983e-11
+    7.271609194321859e-13
+    -1.41388359118495e-13
+   -2.204833930327153e-11
+    7.286023612228777e-11
+ 1.061e+11   
+    7.276106633603063e-11
+    -2.20264781115909e-11
+    8.001507959450098e-11
+   -1.062593959721097e-13
+   -1.366683037715409e-11
+    8.002895967385468e-11
+    7.273448769087739e-13
+   -1.060063642552551e-13
+   -2.202459024208283e-11
+    7.275030153959227e-11
+ 1.066e+11   
+    7.265015561371622e-11
+   -2.200175246853888e-11
+    7.994972185788599e-11
+   -7.072493123860766e-14
+   -1.370482755018179e-11
+    7.996372098412162e-11
+    7.271144584365268e-13
+   -7.048298081954799e-14
+     -2.1999936823891e-11
+    7.263952358668277e-11
+ 1.071e+11   
+    7.253839947606491e-11
+   -2.197611512316186e-11
+    7.988346776314718e-11
+   -3.506107016042518e-14
+   -1.374270598709159e-11
+    7.989758795225678e-11
+    7.264740376821096e-13
+   -3.482954298141354e-14
+   -2.197437357293589e-11
+    7.252790215692843e-11
+ 1.076e+11   
+    7.242579790263339e-11
+   -2.194956069077944e-11
+    7.981631103612725e-11
+    7.205556341142627e-16
+   -1.378045191147669e-11
+     7.98305543213278e-11
+    7.254283820844462e-13
+    9.423404272352052e-16
+   -2.194789512249979e-11
+    7.241543723554276e-11
+ 1.081e+11   
+    7.231235096653033e-11
+   -2.192208389745912e-11
+    7.974824538385175e-11
+    3.660804220362846e-14
+   -1.381805127499188e-11
+    7.976261381490253e-11
+    7.239826524743483e-13
+     3.68207873384151e-14
+   -2.192049621596034e-11
+    7.230212890083033e-11
+ 1.086e+11   
+    7.219805883566165e-11
+   -2.189367958113842e-11
+    7.967926449605732e-11
+    7.258921511132751e-14
+   -1.385548976120957e-11
+    7.969376013855955e-11
+    7.221424024100727e-13
+     7.27936442339184e-14
+   -2.189217170788396e-11
+    7.218797732542439e-11
+ 1.091e+11   
+    7.208292177399763e-11
+   -2.186434269280529e-11
+     7.96093620469145e-11
+    1.086516316197638e-13
+   -1.389275278985356e-11
+    7.962398698154347e-11
+    7.199135770957755e-13
+    1.088484883224148e-13
+   -2.186291656515533e-11
+    7.207298277751554e-11
+ 1.096e+11   
+    7.196694014282744e-11
+   -2.183406829773931e-11
+    7.953853169688188e-11
+    1.447825832808346e-13
+   -1.392982552143052e-11
+    7.955328801862918e-11
+    7.173025119791213e-13
+    1.449726300908587e-13
+   -2.183272586820486e-11
+    7.195714562209765e-11
+ 1.101e+11   
+     7.18501144020011e-11
+   -2.180285157677692e-11
+    7.946676709471306e-11
+    1.809690989063299e-13
+   -1.396669286222062e-11
+    7.948165691205846e-11
+    7.143159309219506e-13
+    1.811531162769893e-13
+   -2.180159481223563e-11
+    7.184046632218884e-11
+ 1.106e+11   
+    7.173244511118993e-11
+    -2.17706878276839e-11
+    7.939406187966044e-11
+    2.171979479487498e-13
+   -1.400333946969347e-11
+     7.94090873137125e-11
+    7.109609440617641e-13
+    2.173767332012621e-13
+   -2.176951870853941e-11
+    7.172294544005768e-11
+ 1.111e+11   
+    7.161393293113561e-11
+   -2.173757246654158e-11
+    7.932040968380604e-11
+    2.534556442740419e-13
+   -1.403974975828038e-11
+    7.933557286741943e-11
+    7.072450452227347e-13
+     2.53630010541648e-13
+   -2.173649298587555e-11
+    7.160458363846254e-11
+ 1.116e+11   
+    7.149457862489216e-11
+   -2.170350102921087e-11
+    7.924580413459127e-11
+    2.897284503342061e-13
+   -1.407590790558211e-11
+    7.926110721143917e-11
+    7.031761090019012e-13
+    2.898992254853958e-13
+   -2.170251319189023e-11
+    7.148538168186984e-11
+ 1.121e+11   
+    7.137438305908326e-11
+   -2.166846917286002e-11
+    7.917023885749779e-11
+    3.260023817693303e-13
+   -1.411179785893661e-11
+    7.918568398110995e-11
+    6.987623874058594e-13
+    3.261704073092762e-13
+   -2.166757499460878e-11
+    7.136534043768532e-11
+ 1.126e+11   
+     7.12533472051446e-11
+   -2.163247267754738e-11
+    7.909370747893811e-11
+    3.622632123995722e-13
+   -1.414740334242597e-11
+    7.910929681169775e-11
+    6.940125061606708e-13
+    3.624293423612654e-13
+   -2.163167418398909e-11
+    7.124446087748363e-11
+ 1.131e+11   
+    7.113147214058472e-11
+   -2.159550744787647e-11
+    7.901620362929263e-11
+    3.984964796393199e-13
+   -1.418270786425859e-11
+    7.903193934139604e-11
+    6.889354605578729e-13
+    3.986615794674723e-13
+   -2.159480667353553e-11
+    7.112274407823738e-11
+ 1.136e+11   
+    7.100875905022098e-11
+   -2.155756951468442e-11
+    7.893772094612442e-11
+    4.346874903123537e-13
+   -1.421769472453117e-11
+    7.895360521450042e-11
+    6.835406109594084e-13
+      4.3485243572846e-13
+   -2.155696850196183e-11
+      7.1000191223539e-11
+ 1.141e+11   
+    7.088520922743805e-11
+   -2.151865503683139e-11
+    7.885825307761007e-11
+    4.708213269087387e-13
+   -1.425234702345841e-11
+    7.887428808481164e-11
+    6.778376778536956e-13
+     4.70987002781546e-13
+   -2.151815583494305e-11
+    7.087680360483494e-11
+ 1.146e+11   
+    7.076082407542738e-11
+   -2.147876030301146e-11
+    7.877779368609556e-11
+    5.068828542189557e-13
+   -1.428664766990793e-11
+    7.879398161913893e-11
+    6.718367365372348e-13
+    5.070501534101916e-13
+   -2.147836496689599e-11
+    7.075258262265008e-11
+ 1.151e+11   
+    7.063560510843777e-11
+   -2.143788173363686e-11
+    7.869633645187217e-11
+    5.428567263959264e-13
+   -1.432057939038039e-11
+    7.871267950104343e-11
+    6.655482113798911e-13
+    5.430265486202231e-13
+   -2.143759232283007e-11
+    7.062752978781033e-11
+ 1.156e+11   
+    7.050955395301308e-11
+   -2.139601588278334e-11
+    7.861387507710712e-11
+    5.787273944431345e-13
+   -1.435412473838111e-11
+    7.863037543474106e-11
+    6.589828696741919e-13
+    5.789006451099151e-13
+   -2.139583446026516e-11
+    7.050164672266883e-11
+ 1.161e+11   
+    7.038267234922147e-11
+   -2.135315944015915e-11
+     7.85304032899386e-11
+    6.144791140570319e-13
+   -1.438726610410944e-11
+    7.854706314913137e-11
+    6.521518150968298e-13
+    6.146567031211848e-13
+    -2.13530880711605e-11
+     7.03749351623083e-11
+ 1.166e+11   
+    7.025496215189202e-11
+   -2.130930923315501e-11
+    7.844591484875842e-11
+    6.500959539257172e-13
+   -1.441998572458484e-11
+    7.846273640206195e-11
+    6.450664807467722e-13
+    6.502787947349695e-13
+   -2.130934998394052e-11
+    7.024739695576155e-11
+ 1.171e+11   
+    7.012642533181802e-11
+   -2.126446222889697e-11
+    7.836040354662076e-11
+    6.855618043798312e-13
+   -1.445226569408775e-11
+    7.837738898470581e-11
+    6.377386217649036e-13
+    6.857508125301098e-13
+   -2.126461716552542e-11
+    7.011903406720111e-11
+ 1.176e+11   
+    6.999706397695913e-11
+   -2.121861553635962e-11
+    7.827386321582493e-11
+    7.208603864434212e-13
+   -1.448408797495009e-11
+    7.829101472608843e-11
+    6.301803075871202e-13
+    7.210564786245367e-13
+   -2.121888672340217e-11
+     6.99898485771183e-11
+ 1.181e+11   
+    6.986688029362922e-11
+   -2.117176640849764e-11
+    7.818628773262959e-11
+    7.559752612643693e-13
+   -1.451543440870018e-11
+    7.820360749778404e-11
+    6.224039137423443e-13
+    7.561793541326611e-13
+   -2.117215590774108e-11
+    6.985984268349597e-11
+ 1.186e+11   
+     6.97358766076473e-11
+   -2.112391224439316e-11
+    7.809767102211511e-11
+    7.908898399039191e-13
+   -1.454628672749766e-11
+    7.811516121870908e-11
+    6.144221132967451e-13
+    7.911028489446967e-13
+   -2.112442211350728e-11
+    6.972901870294628e-11
+ 1.191e+11   
+    6.960405536546901e-11
+   -2.107505059140715e-11
+    7.800800706311818e-11
+    8.255873934861139e-13
+   -1.457662656588159e-11
+    7.802566986006006e-11
+    6.062478678522658e-13
+    8.258102318991141e-13
+   -2.107568288259449e-11
+    6.959737907182133e-11
+ 1.196e+11   
+    6.947141913528834e-11
+   -2.102517914734404e-11
+    7.791728989332042e-11
+    8.600510636856142e-13
+   -1.460643547279441e-11
+    7.793512745034906e-11
+    5.978944182021418e-13
+    8.602846412738832e-13
+   -2.102593590596276e-11
+    6.946492634730562e-11
+ 1.201e+11   
+    6.933797060808525e-11
+    -2.09742957625843e-11
+    7.782551361438559e-11
+    8.942638735403867e-13
+   -1.463569492384031e-11
+    7.784352808050214e-11
+    5.893752745505415e-13
+    8.945090956209293e-13
+   -2.097517902574896e-11
+    6.933166320845093e-11
+ 1.206e+11   
+    6.920371259863809e-11
+   -2.092239844219343e-11
+    7.773267239716774e-11
+    9.282087385786421e-13
+   -1.466438633380425e-11
+    7.775086590904487e-11
+    5.807042063899228e-13
+    9.284665049011281e-13
+   -2.092341023735401e-11
+    6.919759245716797e-11
+ 1.211e+11   
+    6.906864804647091e-11
+   -2.086948534799455e-11
+    7.763876048699056e-11
+    9.618684782388608e-13
+   -1.469249106936751e-11
+    7.765713516733879e-11
+    5.718952319678267e-13
+    9.621396819283663e-13
+   -2.087062769150279e-11
+    6.906271701918188e-11
+ 1.216e+11   
+    6.893278001673941e-11
+   -2.081555480057085e-11
+    7.754377220889178e-11
+     9.95225827551766e-13
+   -1.471999046195902e-11
+    7.756233016481742e-11
+    5.629626074211413e-13
+    9.955113540652888e-13
+   -2.081682969621993e-11
+    6.892703994488757e-11
+ 1.221e+11   
+    6.879611170103974e-11
+   -2.076060528119254e-11
+    7.744770197292233e-11
+    1.028263449075644e-12
+    -1.47468658207949e-11
+    7.746644529423082e-11
+    5.539208155404197e-13
+    1.028564175191219e-12
+   -2.076201471875109e-11
+     6.87905644101606e-11
+ 1.226e+11   
+    6.865864641812315e-11
+   -2.070463543363852e-11
+    7.735054427934749e-11
+    1.060963945062132e-12
+   -1.477309844598774e-11
+    7.736947503684047e-11
+    5.447845541718582e-13
+    1.061280737879846e-12
+   -2.070618138736294e-11
+    6.865329371706849e-11
+ 1.231e+11   
+    6.852038761452429e-11
+    -2.06476440659111e-11
+    7.725229372382608e-11
+    1.093309869807532e-12
+   -1.479866964171014e-11
+    7.727141396756379e-11
+    5.355687243181465e-13
+     1.09364358578155e-12
+   -2.064932849305342e-11
+    6.851523129448502e-11
+ 1.236e+11   
+    6.838133886505929e-11
+   -2.058963015177964e-11
+    7.715294500244171e-11
+    1.125283742174934e-12
+   -1.482356072940422e-11
+    7.717225675999145e-11
+    5.262884179090663e-13
+    1.125635226180183e-12
+   -2.059145499108322e-11
+    6.837638069858964e-11
+ 1.241e+11   
+    6.824150387320101e-11
+   -2.053059283216827e-11
+    7.705249291662532e-11
+    1.156868058262824e-12
+     -1.4847753060945e-11
+    7.707199819128066e-11
+    5.169589052458805e-13
+    1.157238142683836e-12
+   -2.053256000236435e-11
+    6.823674561324556e-11
+ 1.246e+11   
+    6.810088647131571e-11
+   -2.047053141633959e-11
+     7.69509323778495e-11
+    1.188045304164734e-12
+   -1.487122803171971e-11
+    7.697063314684308e-11
+    5.075956221931649e-13
+    1.188434808022275e-12
+   -2.047264281463061e-11
+     6.80963298502274e-11
+ 1.251e+11   
+    6.795949062072602e-11
+   -2.040944538283499e-11
+     7.68482584121104e-11
+    1.218797968793803e-12
+   -1.489396709356868e-11
+    7.686815662480314e-11
+    4.982141570862648e-13
+    1.219207696903696e-12
+   -2.041170288337918e-11
+    6.795513734928899e-11
+ 1.256e+11   
+    6.781732041159438e-11
+   -2.034733438015765e-11
+    7.674446616411527e-11
+    1.249108556738297e-12
+   -1.491595176754033e-11
+    7.676456374018018e-11
+    4.888302373881564e-13
+    1.249539298912112e-12
+   -2.034973983256367e-11
+    6.781317217805594e-11
+ 1.261e+11   
+    6.767438006260721e-11
+   -2.028419822713893e-11
+    7.663955090111005e-11
+     1.27895960109794e-12
+    -1.49371636563866e-11
+    7.665984972871446e-11
+    4.794597161256515e-13
+    1.279412131380688e-12
+   -2.028675345496601e-11
+    6.767043853170821e-11
+ 1.266e+11   
+    6.753067392042606e-11
+   -2.022003691298016e-11
+    7.653350801632873e-11
+    1.308333676252614e-12
+   -1.495758445671536e-11
+    7.655400995029253e-11
+    4.701185581193921e-13
+     1.30880875220662e-12
+   -2.022274371222839e-11
+    6.752694073244569e-11
+ 1.271e+11   
+    6.738620645889598e-11
+   -2.015485059688249e-11
+     7.64263330319366e-11
+    1.337213410524333e-12
+   -1.497719597075706e-11
+    7.644703989191833e-11
+    4.608228260436403e-13
+    1.337711772558723e-12
+   -2.015771073452721e-11
+    6.738268322870561e-11
+ 1.276e+11   
+    6.724098227797798e-11
+    -2.00886396072756e-11
+    7.631802160147834e-11
+    1.365581498667027e-12
+   -1.499598011763042e-11
+    7.633893517014172e-11
+    4.515886663306462e-13
+    1.366103869410336e-12
+   -2.009165481978724e-11
+    6.723767059410256e-11
+ 1.281e+11   
+    6.709500610237006e-11
+   -2.002140444054308e-11
+    7.620856951167958e-11
+    1.393420714141429e-12
+   -1.501391894407792e-11
+    7.622969153287482e-11
+    4.424322949631784e-13
+    1.393967797875886e-12
+   -2.002457643244868e-11
+    6.709190752607426e-11
+ 1.286e+11   
+    6.694828277980792e-11
+   -1.995314575923307e-11
+    7.609797268355695e-11
+    1.420713921105254e-12
+   -1.503099463449915e-11
+      7.6119304860526e-11
+    4.333699831749336e-13
+    1.421286403244387e-12
+   -1.995647620169132e-11
+     6.69453988441931e-11
+ 1.291e+11   
+    6.680081727899342e-11
+   -1.988386438967537e-11
+    7.598622717276329e-11
+    1.447444086053377e-12
+   -1.504718952027137e-11
+    7.600777116635143e-11
+    4.244180431080095e-13
+    1.448042632686979e-12
+    -1.98873549190858e-11
+    6.679814948812024e-11
+ 1.296e+11   
+     6.66526146871335e-11
+    -1.98135613189701e-11
+    7.587332916905329e-11
+    1.473594289063615e-12
+   -1.506248608820707e-11
+     7.58950865959425e-11
+    4.155928134428872e-13
+    1.474219546551532e-12
+   -1.981721353560376e-11
+    6.665016451516071e-11
+ 1.301e+11   
+    6.650368020703897e-11
+   -1.974223769124625e-11
+    7.575927499477518e-11
+    1.499147734525239e-12
+   -1.507686698802666e-11
+    7.578124742575454e-11
+    4.069106450777019e-13
+    1.499800329167623e-12
+   -1.974605315793065e-11
+    6.650144909739783e-11
+ 1.306e+11   
+    6.635401915375934e-11
+   -1.966989480317902e-11
+    7.564406110229581e-11
+    1.524087761343817e-12
+   -1.509031503880626e-11
+    7.566625006056069e-11
+    3.983878868474912e-13
+    1.524768299110986e-12
+   -1.967387504401577e-11
+    6.635200851835501e-11
+ 1.311e+11   
+    6.620363695071016e-11
+   -1.959653409865367e-11
+    7.552768407023781e-11
+    1.548397852474097e-12
+   -1.510281323416975e-11
+    7.555009102973369e-11
+    3.900408713790158e-13
+    1.549106918804957e-12
+    -1.96006805977818e-11
+    6.620184816914962e-11
+ 1.316e+11   
+    6.605253912524801e-11
+   -1.952215716252027e-11
+    7.541014059843084e-11
+    1.572061643750166e-12
+   -1.511434474620659e-11
+    7.543276698223663e-11
+    3.818859010963386e-13
+    1.572799803426674e-12
+   -1.952647136293544e-11
+     6.60509735441105e-11
+ 1.321e+11   
+    6.590073130364848e-11
+   -1.944676571335939e-11
+    7.529142750140386e-11
+    1.595062931880546e-12
+   -1.512489292789403e-11
+    7.531427468017411e-11
+    3.739392344438273e-13
+    1.595830728982538e-12
+   -1.945124901579452e-11
+     6.58993902357926e-11
+ 1.326e+11   
+    6.574821920545205e-11
+   -1.937036159518874e-11
+    7.517154170035262e-11
+     1.61738568154346e-12
+   -1.513444131391903e-11
+    7.519461099082399e-11
+    3.662170723701046e-13
+    1.618183639474352e-12
+   -1.937501535704663e-11
+    6.574710392936437e-11
+ 1.331e+11   
+     6.55950086371157e-11
+   -1.929294676800026e-11
+    7.505048021340433e-11
+    1.639014031467546e-12
+    -1.51429736197581e-11
+     7.50737728769621e-11
+    3.587355451446709e-13
+    1.639842653067759e-12
+   -1.929777230237072e-11
+    6.559412039630863e-11
+ 1.336e+11   
+     6.54411054849268e-11
+   -1.921452329707009e-11
+    7.492824014402575e-11
+    1.659932299396362e-12
+   -1.515047373883104e-11
+     7.49517573853468e-11
+    3.515106995484104e-13
+    1.660792067147366e-12
+    -1.92195218718114e-11
+    6.544044548738187e-11
+ 1.341e+11   
+    6.528651570713295e-11
+   -1.913509334092396e-11
+     7.48048186674444e-11
+    1.680124985830736e-12
+     -1.5156925737567e-11
+    7.482856163322893e-11
+    3.445584865218681e-13
+      1.6810163621381e-12
+   -1.914026617782895e-11
+    6.528608512479644e-11
+ 1.346e+11   
+    6.513124532521224e-11
+    -1.90546591378715e-11
+    7.468021301490585e-11
+    1.699576776423053e-12
+   -1.516231384821042e-11
+    7.470418279270411e-11
+    3.378947493161033e-13
+    1.700500204004906e-12
+   -1.906000741192536e-11
+    6.513104529355513e-11
+ 1.351e+11   
+    6.497530041425911e-11
+   -1.897322299101238e-11
+    7.455442045561201e-11
+     1.71827254291993e-12
+   -1.516662245919929e-11
+    7.457861807273675e-11
+    3.315352122436636e-13
+    1.719228445278594e-12
+   -1.897874782973824e-11
+    6.497533203188728e-11
+ 1.356e+11   
+    6.481868709238956e-11
+   -1.889078725159107e-11
+    7.442743827611899e-11
+    1.736197342506295e-12
+   -1.516983610287103e-11
+    7.445186469868135e-11
+    3.254954700761455e-13
+    1.737186124506256e-12
+   -1.889648973449879e-11
+    6.481895142072605e-11
+ 1.361e+11   
+    6.466141150914128e-11
+   -1.880735430061433e-11
+     7.42992637570747e-11
+    1.753336415440047e-12
+   -1.517193944036757e-11
+    7.432391988912795e-11
+     3.19790978180276e-13
+    1.754358463983757e-12
+   -1.881323545876138e-11
+    6.466190957217274e-11
+ 1.366e+11   
+    6.450347983277278e-11
+   -1.872292652859414e-11
+    7.416989414702203e-11
+    1.769675180819446e-12
+   -1.517291724345623e-11
+    7.419478082985027e-11
+     3.14437043487291e-13
+    1.770730865628917e-12
+   -1.872898734425754e-11
+    6.450421261686879e-11
+ 1.371e+11   
+    6.434489823642169e-11
+   -1.863750631331732e-11
+    7.403932663312944e-11
+    1.785199230365678e-12
+   -1.517275437308386e-11
+    7.406444464465663e-11
+    3.094488163382094e-13
+    1.786288904862729e-12
+   -1.864374771978556e-11
+    6.434586669023059e-11
+ 1.376e+11   
+    6.418567288303933e-11
+   -1.855109599550606e-11
+    7.390755830860172e-11
+    1.799894320043352e-12
+   -1.517143575445478e-11
+    7.393290836295723e-11
+    3.048412833385005e-13
+    1.801018322349433e-12
+   -1.855751887700665e-11
+    6.418687791746541e-11
+ 1.381e+11   
+     6.40258099090444e-11
+    -1.84636978522553e-11
+    7.377458613653441e-11
+     1.81374635939812e-12
+   -1.516894634832219e-11
+    7.380016888377793e-11
+    3.006292612979825e-13
+    1.814905013424766e-12
+   -1.847030304400871e-11
+    6.402725239730366e-11
+ 1.386e+11   
+    6.386531540661556e-11
+   -1.837531406810655e-11
+    7.364040691002932e-11
+    1.826741398421667e-12
+   -1.516527111833179e-11
+    7.366622293604197e-11
+    2.968273923357426e-13
+    1.827935015088742e-12
+   -1.838210235653657e-11
+    6.386699618438687e-11
+ 1.391e+11   
+    6.370419540456126e-11
+   -1.828594670363892e-11
+    7.350501720827566e-11
+    1.838865611811104e-12
+   -1.516039499410201e-11
+    7.353106703483568e-11
+    2.934501402720695e-13
+    1.840094490361783e-12
+   -1.829291882672406e-11
+    6.370611527022541e-11
+ 1.396e+11   
+    6.354245584769027e-11
+   -1.819559766142912e-11
+    7.336841334838898e-11
+     1.85010528042524e-12
+   -1.515430282978643e-11
+    7.339469743343771e-11
+    2.905117884008347e-13
+    1.851369709859775e-12
+   -1.820275430921614e-11
+    6.354461556266472e-11
+ 1.401e+11   
+    6.338010257461098e-11
+   -1.810426864925789e-11
+    7.323059133273922e-11
+    1.860446769804944e-12
+   -1.514697935788189e-11
+    7.325711007084762e-11
+    2.880264387380614e-13
+    1.861747030416139e-12
+   -1.811161046454335e-11
+    6.338250286378788e-11
+ 1.406e+11   
+    6.321714129388819e-11
+    -1.80119611404101e-11
+     7.30915467914999e-11
+    1.869876505535614e-12
+   -1.513840913794349e-11
+     7.31183005145494e-11
+    2.860080128793871e-13
+    1.871212870561973e-12
+   -1.801948871959314e-11
+    6.321978284617241e-11
+ 1.411e+11   
+    6.305357755848536e-11
+   -1.791867633093923e-11
+    7.295127492014892e-11
+    1.878380945322576e-12
+   -1.512857649996469e-11
+    7.297826389824714e-11
+    2.844702545525684e-13
+    1.879753682698556e-12
+   -1.792639022505798e-11
+    6.305646102744385e-11
+ 1.416e+11   
+    6.288941673841566e-11
+   -1.782441509374447e-11
+    7.280977041165764e-11
+    1.885946547553388e-12
+   -1.511746548211222e-11
+    7.283699485428235e-11
+    2.834267339996083e-13
+    1.887355921771205e-12
+    -1.78323158096991e-11
+     6.28925427430385e-11
+ 1.421e+11   
+    6.272466399154103e-11
+   -1.772917792933227e-11
+    7.266702738307688e-11
+    1.892559736210509e-12
+   -1.510505976250876e-11
+    7.269448744047728e-11
+    2.828908542851068e-13
+    1.894006010274503e-12
+   -1.773726593130477e-11
+    6.272803311711572e-11
+ 1.426e+11   
+    6.255932423243938e-11
+   -1.763296491311084e-11
+    7.252303929623405e-11
+    1.898206861901321e-12
+   -1.509134258477912e-11
+    7.255073506108706e-11
+    2.828758596815104e-13
+    1.899690299391093e-12
+   -1.764124062418926e-11
+     6.25629370315481e-11
+ 1.431e+11   
+    6.239340209928225e-11
+   -1.753577563908848e-11
+    7.237779887225195e-11
+    1.902874158877272e-12
+   -1.507629667702943e-11
+    7.240573038160855e-11
+    2.833948462021196e-13
+    1.904395026091118e-12
+   -1.754423944310004e-11
+    6.239725909292027e-11
+ 1.436e+11   
+    6.222690191865614e-11
+   -1.743760915983108e-11
+    7.223129799960718e-11
+    1.906547697812682e-12
+   -1.505990416396374e-11
+    7.225946523710247e-11
+    2.844607744638252e-13
+    1.908106266005845e-12
+   -1.744626140339259e-11
+    6.223100359747696e-11
+ 1.441e+11   
+    6.205982766826709e-11
+   -1.733846392256337e-11
+    7.208352763543165e-11
+    1.909213334204425e-12
+   -1.504214647183671e-11
+    7.211193053381225e-11
+    2.860864849414682e-13
+    1.910809881896228e-12
+   -1.734730491735491e-11
+    6.206417449395823e-11
+ 1.446e+11   
+    6.189218293747756e-11
+   -1.723833770127047e-11
+    7.193447769976082e-11
+    1.910856652180001e-12
+    -1.50230042259115e-11
+    7.196311614371657e-11
+    2.882847157876738e-13
+    1.912491467550172e-12
+   -1.724736772654239e-11
+    6.189677534427054e-11
+ 1.451e+11   
+    6.172397088562807e-11
+   -1.713722752470261e-11
+    7.178413696247082e-11
+    1.911462903592918e-12
+    -1.50024571401489e-11
+     7.18130107917836e-11
+    2.910681232876014e-13
+    1.913136286926684e-12
+   -1.714644683001766e-11
+    6.172880928194498e-11
+ 1.456e+11   
+    6.155519419810329e-11
+   -1.703512960016855e-11
+    7.163249292259193e-11
+    1.911016942206391e-12
+    -1.49804838988121e-11
+    7.166160193563053e-11
+    2.944493051121543e-13
+    1.912729208402969e-12
+   -1.704453840838114e-11
+    6.156027896834003e-11
+ 1.461e+11   
+    6.138585504010413e-11
+   -1.693203923301334e-11
+    7.147953167976955e-11
+    1.909503152835734e-12
+    -1.49570620297066e-11
+     7.15088756373054e-11
+    2.984408264498107e-13
+    1.911254633959668e-12
+   -1.694163774350162e-11
+    6.139118654656062e-11
+ 1.466e+11   
+    6.121595500811979e-11
+   -1.682795074171904e-11
+    7.132523779757531e-11
+    1.906905375317568e-12
+   -1.493216776879843e-11
+    7.135481642698172e-11
+    3.030552491476194e-13
+     1.90869642318449e-12
+   -1.683773913386569e-11
+    6.122153359307045e-11
+ 1.471e+11   
+    6.104549507907494e-11
+   -1.672285736855063e-11
+    7.116959415849428e-11
+    1.903206823178733e-12
+   -1.490577591594479e-11
+    7.119940715828279e-11
+    3.083051639487712e-13
+    1.905037811967978e-12
+   -1.673283580548166e-11
+    6.105132106698898e-11
+ 1.476e+11   
+    6.087447555716594e-11
+   -1.661675118570913e-11
+    7.101258181029924e-11
+    1.898389996911304e-12
+   -1.487785968150845e-11
+     7.10426288550445e-11
+    3.142032259273324e-13
+    1.900261325787716e-12
+   -1.662691981828997e-11
+    6.088054925707583e-11
+ 1.481e+11   
+    6.070289601840601e-11
+   -1.650962299697782e-11
+    7.085417980369778e-11
+     1.89243659177926e-12
+   -1.484839052366477e-11
+    7.088446054934117e-11
+    3.207621932140586e-13
+    1.894348687509955e-12
+   -1.651998196807138e-11
+    6.070921772642675e-11
+ 1.486e+11   
+    6.053075525291568e-11
+   -1.640146223485824e-11
+    7.069436502105351e-11
+    1.885327400095311e-12
+   -1.481733797623015e-11
+    7.072487911058553e-11
+    3.279949690716639e-13
+    1.887280719662467e-12
+   -1.641201168384855e-11
+    6.053732525491541e-11
+ 1.491e+11   
+    6.035805120501927e-11
+   -1.629225685324662e-11
+    7.053311199608864e-11
+    1.877042207970918e-12
+   -1.478466946688052e-11
+    7.056385906563686e-11
+    3.359146473881635e-13
+    1.879037241151256e-12
+   -1.630299692082796e-11
+    6.036486977944426e-11
+ 1.496e+11   
+    6.018478091123631e-11
+   -1.618199321572854e-11
+    7.037039272450014e-11
+    1.867559686548065e-12
+   -1.475035012570384e-11
+     7.04013724098106e-11
+    3.445345616179968e-13
+    1.869596958451007e-12
+   -1.619292404895852e-11
+    6.019184833208716e-11
+ 1.501e+11   
+    6.001094043626853e-11
+   -1.607065597960116e-11
+    7.020617646548909e-11
+    1.856857277767558e-12
+    -1.47143425840456e-11
+    7.023738840880593e-11
+    3.538683372137216e-13
+    1.858937351321466e-12
+   -1.608177773721947e-11
+    6.001825697623359e-11
+ 1.506e+11   
+    5.983652480713152e-11
+   -1.595822797579526e-11
+    7.004042953423466e-11
+      1.8449110747898e-12
+   -1.467660676370847e-11
+    7.007187339158902e-11
+    3.639299475194544e-13
+    1.847034553166825e-12
+   -1.596954083380234e-11
+     5.98440907408686e-11
+ 1.511e+11   
+    5.966152794560045e-11
+    -1.58446900849191e-11
+    6.987311508548773e-11
+    1.831695697242389e-12
+    -1.46370996566373e-11
+    6.990479053438265e-11
+    3.747337731103285e-13
+    1.833863226189448e-12
+   -1.585619424241803e-11
+    5.966934355317521e-11
+ 1.516e+11   
+    5.948594259918555e-11
+   -1.573002110970497e-11
+    6.970419288846499e-11
+    1.817184161490715e-12
+   -1.459577509528887e-11
+    6.973609963596515e-11
+    3.862946645173109e-13
+      1.8193964315812e-12
+   -1.574171679499421e-11
+    5.949400816965819e-11
+ 1.521e+11   
+    5.930976027088439e-11
+   -1.561419764419868e-11
+    6.953361909338531e-11
+    1.801347746255577e-12
+   -1.455258351403273e-11
+    6.956575688460034e-11
+    3.986280082399542e-13
+    1.803605495026512e-12
+   -1.562608512111346e-11
+    5.931807610604419e-11
+ 1.526e+11   
+     5.91329711480204e-11
+   -1.549719394013941e-11
+    6.936134599010053e-11
+    1.784155853930802e-12
+   -1.450747170198826e-11
+    6.939371461704654e-11
+    4.117497958913542e-13
+    1.786459867907506e-12
+   -1.550927351462858e-11
+    5.914153756626512e-11
+ 1.531e+11   
+      5.8955564030511e-11
+   -1.537898177100787e-11
+    6.918732175932887e-11
+    1.765575868063923e-12
+   -1.446038254788818e-11
+    6.921992107018092e-11
+    4.256766963152772e-13
+    1.767926984656665e-12
+   -1.539125379795131e-11
+    5.896438137086931e-11
+ 1.536e+11   
+    5.877752625898041e-11
+   -1.525953029439039e-11
+    6.901149021728114e-11
+    1.745573007553574e-12
+   -1.441125477767985e-11
+    6.904432012596926e-11
+    4.404261304232823e-13
+    1.747972116812403e-12
+   -1.527199518461428e-11
+     5.87865948852658e-11
+ 1.541e+11   
+    5.859884364318237e-11
+   -1.513880591333146e-11
+    6.883379055449472e-11
+      1.7241101782274e-12
+   -1.436002268574789e-11
+    6.886685105066408e-11
+    4.560163484493511e-13
+    1.726558224460812e-12
+   -1.515146414084756e-11
+    5.860816394828098e-11
+ 1.546e+11   
+    5.841950039128114e-11
+   -1.501677213753558e-11
+    6.865415706998074e-11
+    1.701147822580564e-12
+   -1.430661586084535e-11
+     6.86874482292439e-11
+    4.724665092775279e-13
+    1.703645805810918e-12
+   -1.502962424694371e-11
+    5.842907280155633e-11
+ 1.551e+11   
+    5.823947904059125e-11
+   -1.489338944534264e-11
+    6.847251890191628e-11
+    1.676643768573614e-12
+   -1.425095890799542e-11
+    6.850604089643286e-11
+    4.897967613887857e-13
+    1.679192745841957e-12
+   -1.490643605941764e-11
+    5.824930402040606e-11
+ 1.556e+11   
+    5.805876039048841e-11
+    -1.47686151476038e-11
+    6.828879975641888e-11
+    1.650553078558167e-12
+   -1.419297116790852e-11
+    6.832255286571847e-11
+    5.080283249140666e-13
+    1.653154165059948e-12
+   -1.478185697500806e-11
+    5.806883844682388e-11
+ 1.561e+11   
+    5.787732343825503e-11
+   -1.464240325467469e-11
+    6.810291763612821e-11
+    1.622827899516431e-12
+   -1.413256643566538e-11
+    6.813690225816687e-11
+    5.271835742074077e-13
+    1.625482269575331e-12
+   -1.465584109779631e-11
+    5.788765512542333e-11
+ 1.566e+11   
+    5.769514531875331e-11
+   -1.451470434795901e-11
+    6.791478457063871e-11
+    1.593417316007204e-12
+   -1.406965268074279e-11
+    6.794900123304331e-11
+     5.47286120200618e-13
+    1.596126203875887e-12
+   -1.452833911083154e-11
+    5.770573124318115e-11
+ 1.571e+11   
+    5.751220124889193e-11
+   -1.438546545758062e-11
+    6.772430635110217e-11
+    1.562267207361794e-12
+   -1.400413177073042e-11
+     6.77587557225507e-11
+     5.68360891764252e-13
+    1.565031907860648e-12
+   -1.439929815385548e-11
+    5.752304207396397e-11
+ 1.576e+11   
+    5.732846447797838e-11
+   -1.425462994797559e-11
+    6.753138227169169e-11
+    1.529320110892911e-12
+   -1.393589920145707e-11
+    6.756606517337929e-11
+    5.904342151299983e-13
+    1.532141979872456e-12
+   -1.426866170890544e-11
+    5.733956092891666e-11
+ 1.581e+11   
+     5.71439062451468e-11
+   -1.412213741337134e-11
+    6.733590488092668e-11
+    1.494515093055168e-12
+   -1.386484383657232e-11
+    6.737082229804954e-11
+    6.135338903414591e-13
+    1.497395547705321e-12
+   -1.413636949576776e-11
+    5.715525911390634e-11
+ 1.586e+11   
+    5.695849574518456e-11
+   -1.398792358537539e-11
+    6.713775974628175e-11
+    1.457787630778167e-12
+   -1.379084766007028e-11
+    6.717291283948414e-11
+     6.37689263537274e-13
+    1.460728149758524e-12
+   -1.400235737948634e-11
+    5.697010589533819e-11
+ 1.591e+11   
+    5.677220010419242e-11
+   -1.385192025508223e-11
+    6.693682523590584e-11
+    1.419069505346643e-12
+   -1.371378554559901e-11
+    6.697221535259646e-11
+    6.629312937703434e-13
+    1.422071628775277e-12
+     -1.3866557292345e-11
+    5.678406847577606e-11
+ 1.596e+11   
+    5.658498436664687e-11
+   -1.371405521237932e-11
+    6.673297232170068e-11
+    1.378288711518153e-12
+   -1.363352504688585e-11
+     6.67686010071705e-11
+    6.892926128810002e-13
+    1.381354040792058e-12
+   -1.372889717298199e-11
+    5.659711198093184e-11
+ 1.601e+11   
+    5.639681149555842e-11
+   -1.357425220534407e-11
+    6.652606440848959e-11
+    1.335369384788191e-12
+   -1.354992621408185e-11
+    6.656193341672809e-11
+    7.168075768116955e-13
+    1.338499582257648e-12
+    -1.35893009255414e-11
+    5.640919945971446e-11
+ 1.606e+11   
+    5.620764238755452e-11
+   -1.343243092291344e-11
+     6.63159571944749e-11
+    1.290231749967088e-12
+   -1.346284144125735e-11
+    6.635206849858726e-11
+     7.45512306591702e-13
+    1.293428538464628e-12
+   -1.344768840201632e-11
+    5.622029189915946e-11
+ 1.611e+11   
+     5.60174359048372e-11
+   -1.328850700421751e-11
+    6.610249856868052e-11
+    1.242792094530795e-12
+   -1.337211535086025e-11
+     6.61388543707976e-11
+    7.754447170531133e-13
+     1.24605725675205e-12
+   -1.330397541119183e-11
+    5.603034825618906e-11
+ 1.616e+11   
+    5.582614892609041e-11
+   -1.314239207824399e-11
+    6.588552855157496e-11
+    1.192962770421637e-12
+   -1.327758472139156e-11
+    6.592213129213233e-11
+     8.06644531191391e-13
+    1.196298148171001e-12
+   -1.315807375782962e-11
+    5.583932550827049e-11
+ 1.621e+11   
+    5.563373641853275e-11
+   -1.299399383774256e-11
+    6.566487928557615e-11
+    1.140652228289088e-12
+    -1.31790784651003e-11
+     6.57017316518378e-11
+    8.391532779090181e-13
+      1.1440597215751e-12
+   -1.300989131600463e-11
+    5.564717872515986e-11
+ 1.626e+11   
+    5.544015153340754e-11
+     -1.2843216151489e-11
+    6.544037508265585e-11
+    1.085765088351183e-12
+   -1.307641766300451e-11
+    6.547748001635139e-11
+    8.730142707558662e-13
+    1.089246654347292e-12
+   -1.285933214070993e-11
+     5.54538611640224e-11
+ 1.631e+11   
+    5.524534572728894e-11
+    -1.26899592192474e-11
+    6.521183253671083e-11
+    1.028202252323756e-12
+   -1.296941566500822e-11
+    6.524919324062336e-11
+    9.082725651243034e-13
+    1.031759904176949e-12
+   -1.270629662205184e-11
+    5.525932439029956e-11
+ 1.636e+11   
+    5.504926891165428e-11
+   -1.253411977394136e-11
+     6.49790607088141e-11
+    9.678610610436648e-13
+   -1.285787826335623e-11
+    6.501668065218715e-11
+    9.449748912373102e-13
+    9.714968665316572e-13
+   -1.255068168655601e-11
+    5.506351842677024e-11
+ 1.641e+11   
+    5.485186963320749e-11
+   -1.237559133568663e-11
+    6.474186139389233e-11
+     9.04635502573176e-13
+   -1.274160394805157e-11
+    6.477974431648104e-11
+    9.831695601822295e-13
+    9.083515825999827e-13
+   -1.239238105021308e-11
+    5.486639193327734e-11
+ 1.646e+11   
+    5.465309528743153e-11
+   -1.221426452241187e-11
+    6.450002947765727e-11
+    8.384164757022786e-13
+   -1.262038425322887e-11
+    6.453817939225616e-11
+    1.022906340148157e-12
+     8.42215002610679e-13
+   -1.223128552799607e-11
+    5.466789241960416e-11
+ 1.651e+11   
+     5.44528923678301e-11
+   -1.205002742182247e-11
+    6.425335339286977e-11
+    7.690921137865856e-13
+   -1.249400420366523e-11
+    6.429177458615666e-11
+    1.064236300029267e-12
+    7.729753094787035e-13
+    -1.20672834046009e-11
+    5.446796649394293e-11
+ 1.656e+11   
+    5.425120675320713e-11
+   -1.188276602940847e-11
+    6.400161568417829e-11
+    6.965481738682196e-13
+   -1.236224287080134e-11
+    6.404031271567818e-11
+    1.107211617526659e-12
+    7.005183077055929e-13
+    -1.19002608710992e-11
+    5.426656014930917e-11
+ 1.661e+11   
+    5.404798403520112e-11
+   -1.171236475704089e-11
+    6.374459369069507e-11
+    6.206684958822935e-13
+   -1.222487404759515e-11
+    6.378357138970064e-11
+    1.151885348981664e-12
+    6.247278823390483e-13
+   -1.173010253205275e-11
+    5.406361909010919e-11
+ 1.666e+11   
+    5.384316988807396e-11
+   -1.153870701644418e-11
+    6.348206035535159e-11
+    5.413355365518762e-13
+   -1.208166705137669e-11
+     6.35213238156182e-11
+    1.198311158288463e-12
+    5.454865325918107e-13
+   -1.155669198737306e-11
+    5.385908910085787e-11
+ 1.671e+11   
+    5.363671048245507e-11
+    -1.13616758814546e-11
+    6.321378516966236e-11
+     4.58430982218884e-13
+   -1.193238766347508e-11
+    6.325333974168949e-11
+    1.246543002433848e-12
+    4.626759843534439e-13
+    -1.13799124928345e-11
+    5.365291645875052e-11
+ 1.676e+11   
+    5.342855294438193e-11
+   -1.118115483243494e-11
+     6.29395352619212e-11
+    3.718364443660455e-13
+   -1.177679921380277e-11
+    6.297938654266546e-11
+    1.296634771517412e-12
+    3.761778853562176e-13
+   -1.119964770261853e-11
+    5.344504839142014e-11
+ 1.681e+11   
+     5.32186458604896e-11
+   -1.099702858554398e-11
+    6.265907663600495e-11
+     2.81434240959296e-13
+   -1.161466381769951e-11
+    6.269923045584526e-11
+    1.348639881461007e-12
+    2.858745861096027e-13
+   -1.101578249658407e-11
+    5.323543358074389e-11
+ 1.686e+11   
+    5.300693982964453e-11
+   -1.080918400867864e-11
+    6.237217556675114e-11
+    1.871082658933386e-13
+   -1.144574377115993e-11
+     6.24126379735674e-11
+    1.402610818120507e-12
+    1.916500088910053e-13
+   -1.082820389410087e-11
+     5.30240227129926e-11
+ 1.691e+11   
+    5.279338806063029e-11
+   -1.061751112487284e-11
+    6.207860015642868e-11
+    8.874494783801109e-14
+   -1.126980310909101e-11
+     6.21193773966499e-11
+    1.458598632094485e-12
+    9.339060607519452e-14
+   -1.063680205522511e-11
+    5.281076907493589e-11
+ 1.696e+11   
+    5.257794701470399e-11
+   -1.042190420266718e-11
+    6.177812205494622e-11
+   -1.376570145126812e-14
+   -1.108660932938519e-11
+    6.181922055145167e-11
+    1.516652384234777e-12
+   -9.013592126907135e-15
+   -1.044147136875673e-11
+    5.259562919473312e-11
+ 1.701e+11   
+    5.236057709092973e-11
+   -1.022226293150545e-11
+    6.147051834423049e-11
+   -1.205289507062466e-13
+   -1.089593528335571e-11
+    6.151194467102654e-11
+    1.576818542703765e-12
+   -1.156678418819433e-13
+   -1.024211162524453e-11
+    5.237856352552671e-11
+ 1.706e+11   
+    5.214124335117875e-11
+   -1.001849367853574e-11
+    6.115557358460721e-11
+    -2.31644127601151e-13
+    -1.06975612304788e-11
+    6.119733443820339e-11
+    1.639140333361068e-12
+    -2.26671464888935e-13
+   -1.003862927133821e-11
+    5.215953716864275e-11
+ 1.711e+11   
+    5.191991628055329e-11
+   -9.810510821306485e-12
+    6.083308201799307e-11
+   -3.472033169376675e-13
+   -1.049127705234411e-11
+    6.087518418545622e-11
+    1.703657046349505e-12
+   -3.421165473399053e-13
+    -9.83093873999491e-12
+    5.193852063217076e-11
+ 1.716e+11   
+    5.169657257775919e-11
+   -9.598238148750022e-12
+    6.050284991932007e-11
+   -4.672899854716418e-13
+   -1.027688461731287e-11
+    6.054530024302564e-11
+    1.770403302930666e-12
+   -4.620865655887423e-13
+   -9.618963848973589e-12
+    5.171549061947506e-11
+ 1.721e+11   
+    5.147119596864208e-11
+    -9.38161032059312e-12
+     6.01646980838385e-11
+   -5.919775425491718e-13
+   -1.005420028357249e-11
+    6.020750342297137e-11
+    1.839408287898542e-12
+   -5.866549476981493e-13
+   -9.402639257772276e-12
+    5.149043084087221e-11
+ 1.726e+11   
+    5.124377803472361e-11
+   -9.160574372892166e-12
+    5.981846443382904e-11
+   -7.213278481128419e-13
+   -9.823057524155437e-12
+    5.986163162273972e-11
+     1.91069495428355e-12
+   -7.158835824291176e-13
+   -9.181911970749084e-12
+    5.126333284034308e-11
+ 1.731e+11   
+    5.101431904715946e-11
+    -8.93509125487385e-12
+     5.94640067238819e-11
+    -8.55389682189935e-13
+   -9.583309653055861e-12
+     5.95075425274619e-11
+    1.984279208478101e-12
+   -8.498212897813946e-13
+   -8.956742871644393e-12
+    5.103419682773039e-11
+ 1.736e+11   
+    5.078282879513016e-11
+   -8.705137379661806e-12
+    5.910120531927398e-11
+   -9.941971925505838e-13
+   -9.334832626954066e-12
+    5.914511638556016e-11
+    2.060169085362465e-12
+   -9.885022697737091e-13
+   -8.727108272119467e-12
+    5.080303250546923e-11
+ 1.741e+11   
+    5.054932739629335e-11
+   -8.470706168876635e-12
+    5.872996601728946e-11
+   -1.137768339858584e-12
+   -9.077527892299976e-12
+     5.87742588275812e-11
+    2.138363924476037e-12
+   -1.131944548784764e-12
+   -8.493001454351505e-12
+    5.056985987751903e-11
+ 1.746e+11   
+    5.031384607564782e-11
+   -8.231809568603321e-12
+    5.835022287661783e-11
+   -1.286103362150609e-12
+   -8.811325242769012e-12
+     5.83949036934303e-11
+    2.218853559640446e-12
+    -1.28014844528909e-12
+   -8.254434185214043e-12
+    5.033471002688167e-11
+ 1.751e+11   
+    5.007642789799588e-11
+   -7.988479511867471e-12
+    5.796194101539796e-11
+   -1.439183282884549e-12
+   -8.536185647496836e-12
+    5.800701582865998e-11
+    2.301617535749012e-12
+   -1.433095079232303e-12
+    -8.01143817723981e-12
+    5.009762584694203e-11
+ 1.756e+11   
+    4.983712843825319e-11
+   -7.740769300705009e-12
+    5.756511933425669e-11
+   -1.596968488914323e-12
+   -8.252104006213561e-12
+    5.761059380619621e-11
+    2.386624367542127e-12
+   -1.590744951406648e-12
+   -7.764066469486121e-12
+    4.985866271091379e-11
+ 1.761e+11   
+    4.959601637314424e-11
+   -7.488754879205726e-12
+    5.715979311690725e-11
+   -1.759397406540512e-12
+   -7.959111783573327e-12
+    5.720567252613401e-11
+    2.473830856099601e-12
+      -1.753036620974e-12
+   -7.512394699736434e-12
+     4.96178890629817e-11
+ 1.766e+11   
+    4.935317397745789e-11
+   -7.232535967696085e-12
+     5.67460364578047e-11
+   -1.926385305081406e-12
+   -7.657279471856027e-12
+    5.679232564315572e-11
+    2.563181479392152e-12
+    -1.91988551059703e-12
+   -7.256522238244112e-12
+    4.937538691434854e-11
+ 1.771e+11   
+    4.910869750802836e-11
+   -6.972237027609159e-12
+    5.632396446414101e-11
+   -2.097823258166954e-12
+   -7.346718828926191e-12
+    5.637066776887762e-11
+    2.654607873524014e-12
+   -2.091182869388296e-12
+    -6.99657315260185e-12
+    4.913125222740035e-11
+ 1.776e+11   
+    4.886269745904552e-11
+    -6.70800802665726e-12
+    5.589373517831321e-11
+   -2.273577293012292e-12
+    -7.02758483715129e-12
+    5.594085639530534e-11
+    2.748028421167611e-12
+     -2.2667949239471e-12
+    -6.73269697339053e-12
+    4.888559517162749e-11
+ 1.781e+11   
+     4.86152986732034e-11
+   -6.440024974780614e-12
+    5.545555116709556e-11
+   -2.453487757244761e-12
+   -6.700077329001374e-12
+    5.550309348564337e-11
+    2.843347963145528e-12
+   -2.446562247075664e-12
+   -6.465069231114038e-12
+    4.863854023585313e-11
+ 1.786e+11   
+     4.83666402946259e-11
+   -6.168490203087297e-12
+    5.500966072525273e-11
+   -2.637368931332921e-12
+   -6.364442226499995e-12
+    5.505762668019218e-11
+    2.940457648054015e-12
+      -2.630299372231e-12
+   -6.193891736649205e-12
+    4.839022618273354e-11
+ 1.791e+11   
+    4.811687555145796e-11
+   -5.893632360624477e-12
+    5.455635864435895e-11
+   -2.825008912293337e-12
+   -6.020972344665072e-12
+    5.460475006810081e-11
+     3.03923493329731e-12
+   -2.817794679381954e-12
+   -5.919392580079871e-12
+    4.814080583345003e-11
+ 1.796e+11   
+    4.786617135850506e-11
+   -5.615706107428383e-12
+    5.409598650224377e-11
+   -3.016169791124636e-12
+   -5.670007713647364e-12
+    5.414480448035881e-11
+    3.139543748835585e-12
+   -3.008810574669758e-12
+   -5.641825826370161e-12
+    4.789044567299657e-11
+ 1.801e+11   
+     4.76147077333218e-11
+   -5.334991486804468e-12
+    5.362893243478232e-11
+   -3.210588142431631e-12
+   -5.311935380489595e-12
+    5.367817726571024e-11
+    3.241234832426058e-12
+   -3.203083982196062e-12
+   -5.361470890846329e-12
+    4.763932526946467e-11
+ 1.806e+11   
+     4.73626770226458e-11
+   -5.051792965196569e-12
+     5.31556303596697e-11
+   -3.407975840125178e-12
+   -4.947188659222692e-12
+    5.320530151909169e-11
+    3.344146242159115e-12
+    -3.40032716149115e-12
+   -5.078631582870042e-12
+    4.738763650422112e-11
+ 1.811e+11   
+    4.711028294004091e-11
+   -4.766438134196416e-12
+    5.267655863128568e-11
+   -3.608021208268702e-12
+   -4.576245807275483e-12
+    5.272665474166769e-11
+    3.448104048758599e-12
+    -3.60022885902268e-12
+   -4.793634812302624e-12
+     4.71355826137837e-11
+ 1.816e+11   
+    4.685773941997682e-11
+   -4.479276076096712e-12
+    5.219223811660073e-11
+   -3.810390511651234e-12
+    -4.19962811670711e-12
+    5.224275692246725e-11
+    3.552923206532829e-12
+   -3.802455796862677e-12
+   -4.506828960272002e-12
+    4.688337704850108e-11
+ 1.821e+11   
+    4.660526929837135e-11
+   -4.190675401768108e-12
+    5.170322969416888e-11
+     -4.0147297875885e-12
+   -3.817897420275925e-12
+     5.17541680438389e-11
+    3.658408598187799e-12
+    -4.00665449706426e-12
+   -4.218581923239354e-12
+    4.663124215777859e-11
+ 1.826e+11   
+    4.635310283492976e-11
+   -3.901021977338735e-12
+    5.121013119136008e-11
+   -4.220667020681459e-12
+   -3.431653024428598e-12
+    5.126148502643318e-11
+    3.764356245160633e-12
+   -4.212453437564294e-12
+   -3.929278847296996e-12
+    4.637940771656754e-11
+ 1.831e+11   
+    4.610147609879197e-11
+   -3.610716364069497e-12
+    5.071357378907048e-11
+   -4.427814669425317e-12
+   -3.041528093422924e-12
+    5.076533814423225e-11
+    3.870554672001835e-12
+   -4.419465536642987e-12
+   -3.639319577978885e-12
+    4.612810931330705e-11
+ 1.836e+11   
+    4.585062924688313e-11
+   -3.320171003881398e-12
+    5.021421793832425e-11
+   -4.635772574737111e-12
+   -2.648185520320112e-12
+    5.026638695697278e-11
+    3.976786411082139e-12
+   -4.627290972017081e-12
+   -3.349115859801775e-12
+      4.5877586625869e-11
+ 1.841e+11   
+    4.560080473595218e-11
+   -3.029807191453717e-12
+     4.97127488501873e-11
+   -4.844131329803195e-12
+   -2.252313330568055e-12
+    4.976531582784487e-11
+    4.082829633205037e-12
+   -4.835520364942911e-12
+   -3.059088329935983e-12
+    4.562808162033718e-11
+ 1.846e+11   
+     4.53522455289821e-11
+   -2.740051883572124e-12
+    4.920987164119708e-11
+   -5.052476297047961e-12
+   -1.854619671159839e-12
+    4.926282912284898e-11
+    4.188459891707318e-12
+   -5.043738413825046e-12
+   -2.769663363581149e-12
+    4.537983671987946e-11
+ 1.851e+11   
+    4.510519339414307e-11
+   -2.451334409965291e-12
+    4.870630624566725e-11
+   -5.260392680184196e-12
+   -1.455827441191492e-12
+    4.875964623424975e-11
+    4.293451974072746e-12
+    -5.25152817447244e-12
+   -2.481269848924584e-12
+    4.513309301238015e-11
+ 1.856e+11   
+    4.485988747000241e-11
+   -2.164083173498401e-12
+    4.820278225364422e-11
+   -5.467472511515419e-12
+   -1.056668616349125e-12
+    4.825649665459625e-11
+    4.397581868274423e-12
+   -5.458476410988659e-12
+   -2.194336006044419e-12
+    4.488808860585828e-11
+ 1.861e+11   
+    4.461656342278615e-11
+   -1.878722476388445e-12
+    4.770003391875589e-11
+   -5.673325287027587e-12
+   -6.578783112005196e-13
+    4.775411548868597e-11
+    4.500628871454409e-12
+   -5.664180881535928e-12
+   -1.909286434606318e-12
+    4.464505731929587e-11
+ 1.866e+11   
+    4.437545379964435e-11
+   -1.595669716665572e-12
+    4.719879573630129e-11
+   -5.877595412590799e-12
+   -2.601886251367368e-13
+    4.725324007808836e-11
+    4.602377881745707e-12
+   -5.868261207926476e-12
+   -1.626539704879473e-12
+    4.440422804375505e-11
+ 1.871e+11   
+     4.41367905165162e-11
+   -1.315333423763027e-12
+    4.669979923821002e-11
+   -6.079990669628525e-12
+    1.356775893151265e-13
+    4.675460875139714e-11
+    4.702621836195614e-12
+   -6.070376039583974e-12
+   -1.346506977012989e-12
+    4.416582533712111e-11
+ 1.876e+11   
+    4.390080988755383e-11
+   -1.038112940674489e-12
+    4.620377180135688e-11
+   -6.280319689386363e-12
+    5.290124202621072e-13
+    4.625896214940321e-11
+    4.801163758687991e-12
+   -6.270249011067504e-12
+   -1.069591982882936e-12
+     4.39300719227199e-11
+ 1.881e+11   
+    4.366775499354818e-11
+   -7.644002929416076e-13
+    4.571143707549786e-11
+   -6.478496666739655e-12
+     9.19125900159454e-13
+     4.57670417954065e-11
+    4.897816122776013e-12
+   -6.467696572855884e-12
+   -7.961905205531604e-13
+    4.369719250506731e-11
+ 1.886e+11   
+    4.343785197598192e-11
+   -4.945802595682994e-13
+    4.522350979873057e-11
+   -6.674365634612866e-12
+    1.305341988286874e-12
+    4.527956201912602e-11
+     4.99239233211909e-12
+   -6.662608629222097e-12
+   -5.266802265625744e-13
+    4.346741163561688e-11
+ 1.891e+11   
+    4.321123322945753e-11
+   -2.290114957000046e-13
+    4.474066190476733e-11
+   -6.867236990918981e-12
+    1.686989280233299e-12
+    4.479712825037823e-11
+    5.084690874613475e-12
+   -6.854752472216503e-12
+   -2.613889486434942e-13
+    4.324092370684838e-11
+ 1.896e+11   
+     4.29878961827724e-11
+    3.202046075663818e-14
+     4.42634491788762e-11
+   -7.055785183234586e-12
+    2.063411875695647e-12
+    4.432019320440324e-11
+    5.174500481501985e-12
+   -7.043391078488209e-12
+   -5.725240377520166e-16
+    4.301782616145786e-11
+ 1.901e+11   
+    4.276783996443654e-11
+    2.883111468014769e-13
+    4.379229777329178e-11
+   -7.239011985567669e-12
+    2.434012552531314e-12
+    4.384919388426651e-11
+    5.261645035895737e-12
+   -7.227343869455136e-12
+    2.555440952833776e-13
+    4.279811056615665e-11
+ 1.906e+11   
+    4.255118195280651e-11
+    5.396624069137936e-13
+    4.332763497732965e-11
+   -7.416821666983137e-12
+    2.798272377835801e-12
+    4.338466545869103e-11
+    5.346007420505533e-12
+   -7.405828795890552e-12
+     5.06722089618782e-13
+     4.25817906968375e-11
+ 1.911e+11   
+    4.233808959851375e-11
+    7.858438212643019e-13
+    4.286996532057035e-11
+   -7.589466369564387e-12
+    3.155725150041267e-12
+    4.292716891223113e-11
+    5.427501061429597e-12
+   -7.578805665067723e-12
+    7.527196911080713e-13
+    4.236897784492912e-11
+ 1.916e+11   
+    4.212870094550961e-11
+    1.026628426727189e-12
+    4.241980036545348e-11
+    -7.75708105665871e-12
+    3.505936310101158e-12
+    4.247720951719665e-11
+    5.506042795167082e-12
+   -7.746486838145208e-12
+    9.933179514274378e-13
+     4.21598149594556e-11
+ 1.921e+11   
+    4.192311021487908e-11
+     1.26182360512815e-12
+    4.197759381999785e-11
+    -7.91964429659253e-12
+    3.848504109231269e-12
+    4.203522108178106e-11
+    5.581550861105752e-12
+   -7.908982614774547e-12
+    1.228332578858405e-12
+    4.195441522753643e-11
+ 1.926e+11   
+    4.172137777465042e-11
+    1.491276116058966e-12
+     4.15437304686369e-11
+   -8.077058359085701e-12
+    4.183066920283591e-12
+    4.160157474166768e-11
+    5.653951482457567e-12
+   -8.066276914058681e-12
+    1.457614693910286e-12
+     4.17528523709329e-11
+ 1.931e+11   
+    4.152353953257735e-11
+    1.714868109651975e-12
+     4.11185342518108e-11
+   -8.229207666137515e-12
+    4.509307689858514e-12
+    4.117658753979199e-11
+    5.723183324343994e-12
+   -8.218292813814506e-12
+    1.681048178615455e-12
+    4.155516925800629e-11
+ 1.936e+11   
+    4.132961232631006e-11
+     1.93251305663853e-12
+    4.070227608507194e-11
+   -8.375986723160191e-12
+    4.826955400168598e-12
+    4.076052738772456e-11
+    5.789199142443949e-12
+   -8.364940828835689e-12
+    1.898547015042721e-12
+    4.136138596588531e-11
+ 1.941e+11   
+     4.11395968469559e-11
+    2.144152899914676e-12
+    4.029517869076057e-11
+   -8.517311220500441e-12
+    5.135784895545793e-12
+    4.035361589830279e-11
+    5.851965968026797e-12
+   -8.506142466813308e-12
+    2.110053159917709e-12
+     4.11715046222597e-11
+ 1.946e+11   
+    4.095347942946994e-11
+    2.349755953883503e-12
+    3.989741962933482e-11
+   -8.653121558369988e-12
+    5.435615869356803e-12
+    3.995603038871904e-11
+    5.911464680972054e-12
+   -8.641839696239649e-12
+    2.315534749753706e-12
+    4.098551219220071e-11
+ 1.951e+11   
+    4.077123338668297e-11
+    2.549315103969338e-12
+    3.950913360375274e-11
+    -8.78338317610431e-12
+    5.726311354895571e-12
+    3.956790570407372e-11
+    5.967689334567463e-12
+    -8.77199787239942e-12
+    2.514984419191766e-12
+    4.080338227940182e-11
+ 1.956e+11   
+    4.059282018004553e-11
+    2.742846078155263e-12
+    3.913041458716096e-11
+   -8.908085558350078e-12
+    6.007775868882878e-12
+    3.918933612726644e-11
+    6.020646370820715e-12
+   -8.896605830629076e-12
+    2.708417616092111e-12
+    4.062507650709038e-11
+ 1.961e+11   
+    4.041819054168131e-11
+    2.930385700399654e-12
+    3.876131800202511e-11
+   -9.027240696449277e-12
+    6.279953286975761e-12
+    3.882037746034334e-11
+    6.070353780043747e-12
+   -9.015674784881467e-12
+     2.89587086986905e-12
+    4.045054573200287e-11
+ 1.966e+11   
+    4.024728558527127e-11
+    3.111990103186231e-12
+    3.840186302315619e-11
+   -9.140881330316661e-12
+    6.542824508260251e-12
+    3.846104928366376e-11
+    6.116840229041242e-12
+   -9.129236733070273e-12
+    3.077400008697128e-12
+    4.027973119375918e-11
+ 1.971e+11   
+    4.008003791129341e-11
+      3.2877329062906e-12
+    3.805203500814948e-11
+   -9.249059111504512e-12
+    6.796404958424461e-12
+    3.811133736662386e-11
+    6.160144172487278e-12
+   -9.237342670854244e-12
+    3.253078339652197e-12
+    4.011256563464322e-11
+ 1.976e+11   
+    3.991637269963272e-11
+    3.457703380823893e-12
+    3.771178803015538e-11
+   -9.351842753036114e-12
+    7.040741978092364e-12
+    3.777119619150972e-11
+    6.200312958776934e-12
+   -9.340060747725523e-12
+    3.422994813380866e-12
+    3.994897439616178e-11
+ 1.981e+11   
+    3.975620877847285e-11
+    3.622004621325815e-12
+    3.738104747756493e-11
+   -9.449316200783854e-12
+    7.275912140106645e-12
+    3.744055154906852e-11
+    6.237401940226104e-12
+   -9.437474428842888e-12
+    3.587252196893303e-12
+    3.978887648736088e-11
+ 1.986e+11   
+    3.959945965792718e-11
+    3.780751748545913e-12
+    3.705971268314725e-11
+   -9.541576848144523e-12
+    7.502018536410795e-12
+    3.711930316565178e-11
+    6.271473596483677e-12
+   -9.529680696092964e-12
+    3.745965277316197e-12
+     3.96321856161143e-11
+ 1.991e+11   
+    3.944603451797384e-11
+     3.93407016361988e-12
+    3.674765954694008e-11
+   -9.628733809751845e-12
+    7.719188071487236e-12
+    3.680732732504085e-11
+    6.302596679005783e-12
+   -9.616788308630448e-12
+    3.899259117288633e-12
+    3.947881117418965e-11
+ 1.996e+11   
+    3.929583914199303e-11
+    4.082093871594342e-12
+    3.644474312070589e-11
+   -9.710906266617741e-12
+    7.927568795183858e-12
+    3.650447945225281e-11
+    6.330845383345441e-12
+   -9.698916136763358e-12
+    4.047267379876407e-12
+    3.932865916793241e-11
+ 2.001e+11   
+    3.914877678913351e-11
+    4.224963889181043e-12
+    3.615080012602443e-11
+   -9.788221892690906e-12
+    8.127327303388933e-12
+     3.62105966311859e-11
+    6.356298554873122e-12
+   -9.776191579418373e-12
+    4.190130737800584e-12
+    3.918163308801533e-11
+ 2.006e+11   
+    3.900474900064661e-11
+    4.362826748491817e-12
+    3.586565138258463e-11
+   -9.860815370736075e-12
+    8.318646230571845e-12
+    3.592550003258927e-11
+    6.379038932407116e-12
+   -9.848749072881055e-12
+    4.327995378662924e-12
+    3.903763471346192e-11
+ 2.011e+11   
+    3.886365633711599e-11
+    4.495833105477391e-12
+    3.558910412768925e-11
+    -9.92882700346899e-12
+    8.501721853832943e-12
+    3.564899723334525e-11
+    6.399152433149447e-12
+   -9.916728696410065e-12
+    4.461011614838915e-12
+    3.889656484687997e-11
+ 2.016e+11   
+    3.872539904512973e-11
+     4.62413645895851e-12
+    3.532095421221995e-11
+   -9.992401423998561e-12
+    8.676761823918124e-12
+     3.53808844123083e-11
+    6.416727481319131e-12
+   -9.980274878440057e-12
+    4.589332603889386e-12
+    3.875832397942769e-11
+ 2.021e+11   
+    3.858987765335782e-11
+    4.747891983556796e-12
+    3.506098816223975e-11
+    -1.00516864078569e-11
+    8.843983034733239e-12
+    3.512094841187593e-11
+    6.431854381974019e-12
+   -1.003953520536445e-11
+    4.713113182773746e-12
+    3.862281288544572e-11
+ 2.026e+11   
+    3.845699349920818e-11
+     4.86725547753323e-12
+    3.480898509896608e-11
+   -1.010683178727183e-11
+    9.003609639308013e-12
+    3.486896865802385e-11
+    6.444624740723913e-12
+   -1.009465933331649e-11
+     4.83250881685668e-12
+    3.848993314789365e-11
+ 2.031e+11   
+    3.832664918823735e-11
+    4.982382424547353e-12
+    3.456471851300696e-11
+   -1.015798846688509e-11
+    9.155871216932006e-12
+    3.462471893469187e-11
+    6.455130929362689e-12
+   -1.014579800196828e-11
+    4.947674662713348e-12
+     3.83595876167355e-11
+ 2.036e+11   
+    3.819874898929595e-11
+    5.093427166656209e-12
+    3.432795789149873e-11
+   -1.020530753886393e-11
+     9.30100109335164e-12
+     3.43879690111508e-11
+    6.463465596886281e-12
+   -1.019310214815305e-11
+    5.058764742048716e-12
+    3.823168080322609e-11
+ 2.041e+11   
+    3.807319916900704e-11
+    5.200542184478224e-12
+    3.409847019912411e-11
+   -1.024893949429633e-11
+    9.439234813467298e-12
+    3.415848612331877e-11
+    6.469721224903896e-12
+   -1.023672211609407e-11
+    5.165931222657024e-12
+    3.810611921367043e-11
+ 2.046e+11   
+    3.794990826962527e-11
+    5.303877479334797e-12
+    3.387602121593856e-11
+   -1.028903352690432e-11
+    9.570808763902603e-12
+    3.393603631194167e-11
+    6.473989726089341e-12
+   -1.027680696019348e-11
+    5.269323801236531e-12
+    3.798281162668148e-11
+ 2.051e+11   
+    3.782878733461865e-11
+    5.403580051334318e-12
+    3.366037673651173e-11
+   -1.032573692444202e-11
+    9.695958941113858e-12
+    3.372038562213277e-11
+    6.476362084039992e-12
+   -1.031350383568821e-11
+    5.369089182030684e-12
+    3.786166931826082e-11
+ 2.056e+11   
+    3.770975008648223e-11
+    5.499793466757208e-12
+     3.34513036361354e-11
+   -1.035919454265593e-11
+     9.81491985934176e-12
+    3.351130117000925e-11
+    6.476928032708331e-12
+   -1.034695747200433e-11
+    5.465370644659474e-12
+    3.774260623919271e-11
+ 2.061e+11   
+    3.759271306133985e-11
+    5.592657507707672e-12
+    3.324857081078568e-11
+   -1.038954835635194e-11
+    9.927923591653759e-12
+    3.330855208310173e-11
+    6.475775773427925e-12
+   -1.037730972332277e-11
+    5.558307694114413e-12
+    3.762553914929654e-11
+ 2.066e+11   
+    3.747759570484758e-11
+    5.682307896794798e-12
+    3.305194999819384e-11
+   -1.041693708192324e-11
+    1.003519893654698e-11
+    3.311191032188009e-11
+    6.472991727466672e-12
+   -1.040469919068425e-11
+     5.64803578568781e-12
+    3.751038771303725e-11
+ 2.071e+11   
+    3.736432043378882e-11
+     5.76887608956444e-12
+    3.286121648781207e-11
+   -1.044149586562052e-11
+    1.013697070205415e-11
+    3.292115139017237e-11
+    6.468660321992935e-12
+   -1.042926090989864e-11
+    5.734686117565203e-12
+    3.739707456087628e-11
+ 2.076e+11   
+    3.725281266756936e-11
+    5.852489127497867e-12
+    3.267614972769086e-11
+   -1.046335603187783e-11
+    1.023345909897704e-11
+     3.27360549424849e-11
+    6.462863807326435e-12
+    -1.04511260995573e-11
+    5.818385483905502e-12
+    3.728552532056134e-11
+ 2.081e+11   
+    3.714300083359089e-11
+    5.933269544599476e-12
+    3.249653383634599e-11
+   -1.048264488611827e-11
+    1.032487923473935e-11
+    3.255640529629515e-11
+    6.455682103359696e-12
+   -1.047042196356419e-11
+    5.899256181438551e-12
+    3.717566862232913e-11
+ 2.086e+11   
+     3.70348163502218e-11
+    6.011335320889432e-12
+    3.232215802761643e-11
+   -1.049948556664484e-11
+    1.041144069937022e-11
+    3.238199185731308e-11
+    6.447192673069563e-12
+   -1.048727154278286e-11
+    5.977415962904528e-12
+    3.706743608173267e-11
+ 2.091e+11   
+    3.692819359079966e-11
+    6.086799876480569e-12
+    3.215281695632662e-11
+   -1.051399694045001e-11
+    1.049334723527444e-11
+    3.221260946552139e-11
+    6.437470421087693e-12
+   -1.050179361062845e-11
+    6.052978031021664e-12
+    3.696076226352582e-11
+ 2.096e+11   
+       3.682306983181e-11
+    6.159772100328446e-12
+    3.198831099229255e-11
+   -1.052629353804627e-11
+    1.057079648269052e-11
+    3.204805866953027e-11
+    6.426587615359559e-12
+   -1.051410260770247e-11
+    6.126051067077945e-12
+    3.685558462974392e-11
+ 2.101e+11   
+    3.671938518808524e-11
+    6.230356408186889e-12
+    3.182844642987079e-11
+   -1.053648552271189e-11
+    1.064397979306124e-11
+     3.18881459364458e-11
+     6.41461382998985e-12
+   -1.052430861086198e-11
+    6.196739288687381e-12
+    3.675184347482511e-11
+ 2.106e+11   
+    3.661708253758107e-11
+     6.29865282476323e-12
+    3.167303563986574e-11
+   -1.054467868985655e-11
+    1.071308210292341e-11
+    3.173268380406576e-11
+    6.401615907446887e-12
+   -1.053251733242482e-11
+    6.265142531709762e-12
+    3.664948185032483e-11
+ 2.111e+11   
+    3.651610743799817e-11
+    6.364757085534571e-12
+    3.152189717019387e-11
+   -1.055097449252537e-11
+    1.077828186134635e-11
+    3.158149098180218e-11
+    6.387657938374592e-12
+    -1.05388301455289e-11
+    6.331356351802496e-12
+    3.654844548149281e-11
+ 2.116e+11   
+     3.64164080372529e-11
+    6.428760754149302e-12
+    3.137485580126883e-11
+   -1.055547008938077e-11
+    1.083975100439778e-11
+    3.143439240629716e-11
+    6.372801257342174e-12
+   -1.054334413198129e-11
+    6.395472141534323e-12
+    3.644868267771353e-11
+ 2.121e+11   
+    3.631793497954198e-11
+    6.490751351791037e-12
+    3.123174256163597e-11
+    -1.05582584118101e-11
+    1.089765497058168e-11
+    3.129121925725947e-11
+    6.357104452940567e-12
+   -1.054615214924591e-11
+    6.457577259442619e-12
+    3.635014423855568e-11
+ 2.126e+11   
+     3.62206413085125e-11
+    6.550812495314999e-12
+    3.109239470894408e-11
+   -1.055942824711391e-11
+    1.095215275165949e-11
+    3.115180893861387e-11
+    6.340623390716236e-12
+   -1.054734291352194e-11
+    6.517755167849473e-12
+    3.625278335694111e-11
+ 2.131e+11   
+    3.612448236883071e-11
+    6.609024041377047e-12
+    3.095665568091564e-11
+   -1.055906433501918e-11
+    1.100339697373077e-11
+    3.101600502962661e-11
+    6.323411247513834e-12
+   -1.054700109615659e-11
+    6.576085576661309e-12
+    3.615655552072662e-11
+ 2.136e+11   
+    3.602941570724503e-11
+    6.665462234160142e-12
+    3.082437502056531e-11
+   -1.055724747504037e-11
+    1.105153400390453e-11
+    3.088365721025809e-11
+    6.305518555878438e-12
+   -1.054520743091418e-11
+    6.632644590760037e-12
+    3.606141841379361e-11
+ 2.141e+11   
+     3.59354009740614e-11
+    6.720199854658322e-12
+    3.069540827951853e-11
+    -1.05540546424713e-11
+     1.10967040783285e-11
+    3.075462116459831e-11
+    6.286993257248023e-12
+   -1.054203882988371e-11
+    6.687504858949946e-12
+    3.596733181756422e-11
+ 2.146e+11   
+    3.584239982578905e-11
+    6.773306369803161e-12
+    3.056961690290996e-11
+   -1.054955911103708e-11
+    1.113904144776366e-11
+     3.06287584658673e-11
+     6.26788076274424e-12
+    -1.05375685060523e-11
+    6.740735722747974e-12
+    3.587425751370058e-11
+ 2.151e+11   
+    3.575037582957379e-11
+    6.824848080013845e-12
+    3.044686809898995e-11
+   -1.054383058045996e-11
+    1.117867453728734e-11
+    3.050593644611064e-11
+    6.248224020446397e-12
+   -1.053186610079887e-11
+    6.792403363601388e-12
+    3.578215918860555e-11
+ 2.156e+11   
+    3.565929436991349e-11
+    6.874888264016232e-12
+    3.032703469623889e-11
+   -1.053693530740599e-11
+    1.121572611708028e-11
+    3.038602805339282e-11
+    6.228063588109368e-12
+   -1.052499781477274e-11
+     6.84257094738015e-12
+    3.569100234021756e-11
+ 2.161e+11   
+    3.556912255803896e-11
+    6.923487320012118e-12
+    3.020999499048468e-11
+   -1.052893623846891e-11
+    1.125031348160028e-11
+    3.026891169898576e-11
+    6.207437710358995e-12
+   -1.051702654081402e-11
+    6.891298765227817e-12
+    3.560075418748418e-11
+ 2.166e+11   
+    3.547982914425468e-11
+    6.970702902488906e-12
+    3.009563258424033e-11
+   -1.051989314402674e-11
+     1.12825486347673e-11
+     3.01544710967713e-11
+    6.186382399471202e-12
+   -1.050801199774955e-11
+    6.938644370061936e-12
+    3.551138358280635e-11
+ 2.171e+11   
+    3.539138443344923e-11
+    7.016590054139375e-12
+    2.998383622021797e-11
+   -1.050986275196469e-11
+    1.131253847908045e-11
+    3.004259509681658e-11
+     6.16493151891104e-12
+    -1.04980108640582e-11
+    6.984662708195759e-12
+    3.542286092766442e-11
+ 2.176e+11   
+    3.530376020392129e-11
+    7.061201332519686e-12
+    2.987449961074407e-11
+   -1.049889888040503e-11
+    1.134038500685958e-11
+    2.993317751484776e-11
+    6.143116868875872e-12
+   -1.048707691054481e-11
+    7.029406245709944e-12
+    3.533515809156964e-11
+ 2.181e+11   
+     3.52169296296067e-11
+    7.104586931206675e-12
+      2.9767521264583e-11
+   -1.048705256871341e-11
+    1.136618549205052e-11
+    2.982611695913096e-11
+    6.120968273152541e-12
+   -1.047526113129263e-11
+    7.072925089336094e-12
+     3.52482483344268e-11
+ 2.186e+11   
+    3.513086720574628e-11
+    7.146794795328149e-12
+    2.966280431248496e-11
+   -1.047437220617093e-11
+    1.139003268125867e-11
+    2.972131665607802e-11
+    6.098513666662595e-12
+   -1.046261187228236e-11
+    7.115267101726667e-12
+    3.516210623234624e-11
+ 2.191e+11   
+    3.504554867799423e-11
+    7.187870731435103e-12
+    2.956025633259654e-11
+   -1.046090365780458e-11
+    1.141201498287632e-11
+    2.961868427571577e-11
+    6.075779183129983e-12
+    -1.04491749571706e-11
+    7.156478011080198e-12
+    3.507670760690469e-11
+ 2.196e+11   
+    3.496095097493481e-11
+    7.227858511760761e-12
+    2.945978917671513e-11
+    -1.04466903869635e-11
+    1.143221665335148e-11
+    2.951813175800132e-11
+    6.052789242364422e-12
+   -1.043499380981423e-11
+     7.19660151516705e-12
+    3.499202945782097e-11
+ 2.201e+11   
+    3.487705214394912e-11
+    7.266799972973869e-12
+    2.936131879822684e-11
+   -1.043177357431065e-11
+    1.145071797980893e-11
+      2.9419575140823e-11
+     6.02956663670947e-12
+   -1.042010957321102e-11
+    7.235679379863239e-12
+    3.490804989898848e-11
+ 2.206e+11   
+    3.479383129035438e-11
+    7.304735109582706e-12
+    2.926476508243958e-11
+   -1.041619223297395e-11
+    1.146759545837812e-11
+    2.932293439039982e-11
+    6.006132616256854e-12
+   -1.040456122459917e-11
+    7.273751532348181e-12
+    3.482474809778467e-11
+ 2.211e+11   
+    3.471126851972162e-11
+    7.341702162183442e-12
+    2.917005167990964e-11
+    -1.03999833196639e-11
+    1.148292196770938e-11
+     2.92281332346771e-11
+    5.982506972478965e-12
+   -1.038838568652394e-11
+    7.310856149160208e-12
+    3.474210421756346e-11
+ 2.216e+11   
+    3.462934488326678e-11
+    7.377737700773285e-12
+    2.907710584325964e-11
+   -1.038318184162288e-11
+    1.149676693727483e-11
+    2.913509900021717e-11
+    5.958708119978192e-12
+   -1.037161793373515e-11
+    7.347029739329606e-12
+    3.466009936322365e-11
+ 2.221e+11   
+    3.454804232620086e-11
+    7.412876703368273e-12
+    2.898585826789534e-11
+    -1.03658209593189e-11
+    1.150919651014767e-11
+    2.904376245299259e-11
+    5.934753176096023e-12
+    -1.03542910958293e-11
+    7.382307222828847e-12
+    3.457871552973912e-11
+ 2.226e+11   
+    3.446734363892082e-11
+    7.447152630176869e-12
+    2.889624293695006e-11
+   -1.034793208483966e-11
+    1.152027370003964e-11
+    2.895405764340941e-11
+    5.910658038165893e-12
+   -1.033643655559185e-11
+    7.416722004590174e-12
+    3.449793555353037e-11
+ 2.231e+11   
+    3.438723241091751e-11
+    7.480597493585877e-12
+    2.880819697071469e-11
+   -1.032954497597952e-11
+    1.153005854245221e-11
+    2.886592175581992e-11
+    5.886437458231551e-12
+   -1.031808404303209e-11
+    7.450306044347031e-12
+    3.441774306655416e-11
+ 2.236e+11   
+    3.430769298727807e-11
+    7.513241924215862e-12
+    2.872166048075043e-11
+   -1.031068782604294e-11
+    1.153860823986049e-11
+    2.877929496272063e-11
+    5.862105115088453e-12
+    -1.02992617251343e-11
+    7.483089922555433e-12
+    3.433812245298596e-11
+ 2.241e+11   
+    3.422871042765698e-11
+     7.54511523330001e-12
+    2.863657642882663e-11
+    -1.02913873494138e-11
+    1.154597730090405e-11
+    2.869412028377819e-11
+    5.837673683537167e-12
+    -1.02799962913748e-11
+    7.515102902649116e-12
+    3.425905880837098e-11
+ 2.246e+11   
+    3.415027046759509e-11
+    7.576245471633436e-12
+    2.855289049078006e-11
+   -1.027166886296298e-11
+    1.155221767360696e-11
+    2.861034344977889e-11
+     5.81315490076849e-12
+   -1.026031303507738e-11
+    7.546372989874021e-12
+    3.418053790112008e-11
+ 2.251e+11   
+    3.407235948206453e-11
+    7.606659485331017e-12
+    2.847055092534963e-11
+   -1.025155636338434e-11
+     1.15573788726861e-11
+    2.852791277155529e-11
+    5.788559629825008e-12
+   -1.024023593069725e-11
+    7.576926986940372e-12
+    3.410254613622954e-11
+ 2.256e+11   
+    3.399496445112323e-11
+    7.636382968621122e-12
+    2.838950844800628e-11
+    -1.02310726005643e-11
+    1.156150810104283e-11
+    2.844677901391004e-11
+    5.763897920109498e-12
+   -1.021978770713855e-11
+    7.606790546718346e-12
+    3.402507052110616e-11
+ 2.261e+11   
+    3.391807292756451e-11
+    7.665440513889585e-12
+    2.830971610976644e-11
+    -1.02102391471023e-11
+    1.156465036555721e-11
+    2.836689527452418e-11
+    5.739179064931658e-12
+   -1.019898991722338e-11
+    7.635988222191879e-12
+    3.394809863338448e-11
+ 2.266e+11   
+    3.384167300645159e-11
+    7.693855659176725e-12
+    2.823112918095211e-11
+   -1.018907646410787e-11
+    1.156684858732813e-11
+    2.828821686781265e-11
+    5.714411656103507e-12
+   -1.017786300343801e-11
+    7.664543513871678e-12
+    3.387161859062393e-11
+ 2.271e+11   
+    3.376575329643204e-11
+    7.721650933314879e-12
+    2.815370503983741e-11
+    -1.01676039634091e-11
+    1.156814370651825e-11
+    2.821070121366685e-11
+    5.689603635611402e-12
+   -1.015642636009059e-11
+     7.69247891485527e-12
+     3.37956190217806e-11
+ 2.276e+11   
+    3.369030289272962e-11
+    7.748847898881852e-12
+    2.807740306610383e-11
+   -1.014584006630963e-11
+    1.156857478197722e-11
+    2.813430773100578e-11
+    5.664762344406927e-12
+   -1.013469839201877e-11
+    7.719815953708395e-12
+    3.372008904035206e-11
+ 2.281e+11   
+    3.361531135171745e-11
+     7.77546719313059e-12
+    2.800218453900996e-11
+   -1.012380225903712e-11
+    1.156817908582663e-11
+    2.805899773604153e-11
+    5.639894568372582e-12
+   -1.011269656998884e-11
+    7.746575235327883e-12
+    3.364501821909726e-11
+ 2.286e+11   
+    3.354076866697977e-11
+     7.80152856704394e-12
+    2.792801254016919e-11
+   -1.010150714502559e-11
+    1.156699219319631e-11
+    2.798473434515138e-11
+    5.615006581528195e-12
+   -1.009043748293059e-11
+    7.772776479933614e-12
+    3.357039656623931e-11
+ 2.291e+11   
+    3.346666524677412e-11
+    7.827050922648377e-12
+    2.785485186081776e-11
+    -1.00789704941771e-11
+    1.156504806730676e-11
+    2.791148238224007e-11
+    5.590104186553888e-12
+   -1.006793688715154e-11
+    7.798438560323993e-12
+    3.349621450306265e-11
+ 2.296e+11   
+     3.33929918928109e-11
+    7.852052348710055e-12
+    2.778266891344829e-11
+   -1.005620728924492e-11
+    1.156237914009538e-11
+    2.783920829046559e-11
+    5.565192752713474e-12
+   -1.004520975267453e-11
+    7.823579537517066e-12
+    3.342246284282139e-11
+ 2.301e+11   
+    3.331973978027052e-11
+    7.876550154924344e-12
+    2.771143164767616e-11
+   -1.003323176948068e-11
+    1.155901638858275e-11
+    2.776788004819639e-11
+    5.540277251267353e-12
+   -1.002227030684023e-11
+     7.84821669488821e-12
+    3.334913277087894e-11
+ 2.306e+11   
+    3.324690043898402e-11
+    7.900560904698656e-12
+    2.764110947020289e-11
+   -1.001005747168531e-11
+    1.155498940717672e-11
+    2.769746708906357e-11
+     5.51536228847037e-12
+   -9.999132075314692e-12
+    7.872366570903892e-12
+    3.327621582600451e-11
+ 2.311e+11   
+    3.317446573570506e-11
+    7.924100446619081e-12
+    2.757167316873483e-11
+   -9.986697268799738e-12
+    1.155032647610667e-11
+    2.762794022596692e-11
+    5.490452136252187e-12
+   -9.975807920637916e-12
+    7.896044990541963e-12
+     3.32037038827552e-11
+ 2.316e+11   
+    3.310242785740771e-11
+    7.947183944681578e-12
+    2.750309483971727e-11
+   -9.963163406169036e-12
+    1.154505462617997e-11
+    2.755927157889317e-11
+    5.465550760681859e-12
+   -9.952310078447469e-12
+    7.919267095478119e-12
+    3.313158913487652e-11
+ 2.321e+11   
+    3.303077929554557e-11
+    7.969825907359759e-12
+    2.743534781973838e-11
+   -9.939467535608668e-12
+    1.153919970004526e-11
+    2.749143450640226e-11
+    5.440661848319333e-12
+   -9.928650191505541e-12
+    7.942047373110922e-12
+    3.305986407965888e-11
+ 2.326e+11   
+    3.295951283121352e-11
+    7.992040215574014e-12
+     2.73684066204612e-11
+   -9.915620747398079e-12
+    1.153278641014455e-11
+    2.742440354063918e-11
+    5.415788830556951e-12
+   -9.904839341654781e-12
+    7.964399684490011e-12
+    3.298852150318994e-11
+ 2.331e+11   
+    3.288862152115536e-11
+    8.013840149618856e-12
+    2.730224686694042e-11
+   -9.891633600321861e-12
+    1.152583839352901e-11
+    2.735815432572751e-11
+    5.390934906055027e-12
+   -9.880888079823158e-12
+    7.986337291203715e-12
+    3.291755446644707e-11
+ 2.336e+11   
+    3.281809868456522e-11
+    8.035238415100297e-12
+    2.723684523918261e-11
+   -9.867516149874228e-12
+    1.151837826370735e-11
+    2.729266355940381e-11
+    5.366103061374249e-12
+   -9.856806454193922e-12
+    8.007872881277387e-12
+    3.284695629217719e-11
+ 2.341e+11   
+    3.274793789063228e-11
+     8.05624716792795e-12
+    2.717217941681095e-11
+   -9.843277974737313e-12
+    1.151042765969047e-11
+    2.722790893775368e-11
+    5.341296089906705e-12
+   -9.832604036650535e-12
+    8.029018594128261e-12
+    3.277672055251445e-11
+ 2.346e+11   
+    3.267813294678223e-11
+    8.076878038402395e-12
+    2.710822802669705e-11
+   -9.818928201639662e-12
+    1.150200729238798e-11
+    2.716386910291219e-11
+    5.316516609205467e-12
+   -9.808289947603614e-12
+    8.049786044615644e-12
+    3.270684105728899e-11
+ 2.351e+11   
+    3.260867788757225e-11
+    8.097142154433838e-12
+    2.704497059342607e-11
+    -9.79447552869591e-12
+    1.149313698850633e-11
+    2.710052359359467e-11
+    5.291767076810598e-12
+   -9.783872879300281e-12
+    8.070186346223779e-12
+    3.263731184298351e-11
+ 2.356e+11   
+    3.253956696419699e-11
+    8.117050163924248e-12
+    2.698238749246482e-11
+   -9.769928247322936e-12
+    1.148383573209134e-11
+    2.703785279832703e-11
+    5.267049804666907e-12
+   -9.759361117712176e-12
+    8.090230133408161e-12
+    3.256812716229646e-11
+ 2.361e+11   
+     3.24707946345682e-11
+    8.136612256341299e-12
+    2.692045990590358e-11
+   -9.745294262825068e-12
+    1.147412170385093e-11
+    2.697583791124801e-11
+    5.242366972225772e-12
+   -9.734762563092792e-12
+    8.109927583134767e-12
+    3.249928147427244e-11
+ 2.366e+11   
+    3.240235555393048e-11
+    8.155838183510163e-12
+    2.685916978065024e-11
+   -9.720581113733422e-12
+    1.146401231838777e-11
+     2.69144608903597e-11
+    5.217720638320667e-12
+   -9.710084749291762e-12
+    8.129288435637199e-12
+    3.243076943496557e-11
+ 2.371e+11   
+    3.233424456598003e-11
+     8.17473727964644e-12
+    2.679849978895461e-11
+   -9.695795989982076e-12
+    1.145352425946399e-11
+    2.685370441810637e-11
+    5.193112751902193e-12
+   -9.685334861906486e-12
+    8.148322014415612e-12
+     3.23625858886002e-11
+ 2.376e+11   
+    3.226645669445376e-11
+    8.193318480651726e-12
+     2.67384332911478e-11
+   -9.670945749997596e-12
+    1.144267351341419e-11
+    2.679355186416496e-11
+    5.168545161715291e-12
+    -9.66051975534887e-12
+    8.167037245498624e-12
+    3.229472585919831e-11
+ 2.381e+11   
+    3.219898713515958e-11
+    8.211590342690768e-12
+     2.66789543004846e-11
+   -9.646036936775142e-12
+    1.143147540081719e-11
+    2.673398725033645e-11
+    5.144019624998006e-12
+   -9.635645968899819e-12
+    8.185442675987224e-12
+    3.222718454264362e-11
+ 2.386e+11   
+    3.213183124841883e-11
+    8.229561060069004e-12
+    2.662004744997981e-11
+   -9.621075793008772e-12
+      1.1419944606529e-11
+    2.667499521742772e-11
+    5.119537815276893e-12
+   -9.610719741819672e-12
+    8.203546491899256e-12
+     3.21599572991545e-11
+ 2.391e+11   
+    3.206498455189585e-11
+    8.247238482426649e-12
+    2.656169796113586e-11
+   -9.596068275341356e-12
+    1.140809520817643e-11
+     2.66165609940232e-11
+    5.095101329331277e-12
+   -9.585747027578799e-12
+    8.221356535331252e-12
+     3.20930396461403e-11
+ 2.396e+11   
+    3.199844271378947e-11
+     8.26463013126644e-12
+    2.650389161445997e-11
+   -9.571020067792826e-12
+    1.139594070320144e-11
+    2.655867036704288e-11
+    5.070711693394214e-12
+   -9.560733507268453e-12
+    8.238880320953771e-12
+    3.202642725141606e-11
+ 2.401e+11   
+    3.193220154636315e-11
+    8.281743215828874e-12
+    2.644661472167682e-11
+   -9.545936594424441e-12
+    1.138349403454486e-11
+    2.650130965399366e-11
+    5.046370368654842e-12
+   -9.535684602248434e-12
+    8.256125051855061e-12
+    3.196011592675325e-11
+ 2.406e+11   
+    3.186625699979356e-11
+    8.298584648331168e-12
+    2.638985409954272e-11
+   -9.520823031291015e-12
+    1.137076761504887e-11
+    2.644446567682008e-11
+    5.022078756123065e-12
+   -9.510605486083939e-12
+    8.273097634748661e-12
+    3.189410162174584e-11
+ 2.411e+11   
+    3.180060515631663e-11
+    8.315161058583164e-12
+    2.633359704517482e-11
+   -9.495684317730882e-12
+    1.135777335065579e-11
+    2.638812573726788e-11
+    4.997838200913801e-12
+   -9.485501095821059e-12
+    8.289804694558551e-12
+    3.182838041797114e-11
+ 2.416e+11   
+    3.173524222465252e-11
+    8.331478807995332e-12
+    2.627783131281009e-11
+   -9.470525167038552e-12
+    1.134452266247409e-11
+      2.6332277593675e-11
+    4.973649996004649e-12
+   -9.460376142646448e-12
+    8.306252588396583e-12
+    3.176294852342759e-11
+ 2.421e+11   
+    3.167016453469268e-11
+    8.347544002991681e-12
+    2.622254509191428e-11
+   -9.445350076564133e-12
+     1.13310265077788e-11
+    2.627690943911111e-11
+    4.949515385517655e-12
+   -9.435235121974125e-12
+    8.322447418945802e-12
+    3.169780226723212e-11
+ 2.426e+11   
+    3.160536853243231e-11
+     8.36336250784273e-12
+    2.616772698656321e-11
+   -9.420163337277914e-12
+    1.131729540000858e-11
+    2.622200988078741e-11
+    4.925435567572004e-12
+    -9.41008232299872e-12
+    8.338395047263956e-12
+    3.163293809456092e-11
+ 2.431e+11   
+    3.154085077513316e-11
+    8.378939956931439e-12
+    2.611336599602437e-11
+    -9.39496904283775e-12
+     1.13033394278184e-11
+    2.616756792066458e-11
+    4.901411696751985e-12
+   -9.384921837752373e-12
+    8.354101105020776e-12
+    3.156835256181915e-11
+ 2.436e+11   
+    3.147660792670339e-11
+     8.39428176646671e-12
+    2.605945149646806e-11
+   -9.369771098193329e-12
+    1.128916827324232e-11
+    2.611357293718969e-11
+     4.87744488623103e-12
+   -9.359757569699177e-12
+    8.369571006183507e-12
+    3.150404233202579e-11
+ 2.441e+11   
+    3.141263675327985e-11
+     8.40939314565817e-12
+    2.600597322374237e-11
+   -9.344573227758721e-12
+    1.127479122901713e-11
+    2.606001466809422e-11
+    4.853536209589316e-12
+    -9.33459324189876e-12
+    8.384809958164202e-12
+    3.144000417039971e-11
+ 2.446e+11   
+    3.134893411900303e-11
+    8.424279107366816e-12
+     2.59529212571488e-11
+   -9.319378983183014e-12
+    1.126021721511501e-11
+    2.600688319419209e-11
+    4.829686702360795e-12
+   -9.309432404768543e-12
+     8.39982297244364e-12
+    3.137623494013683e-11
+ 2.451e+11   
+    3.128549698197108e-11
+    8.438944478245253e-12
+    2.590028600415878e-11
+   -9.294191750745418e-12
+    1.124545479452935e-11
+    2.595416892411691e-11
+    4.805897363341616e-12
+     -9.2842784434715e-12
+    8.414614874685632e-12
+    3.131273159836598e-11
+ 2.456e+11   
+    3.122232239036399e-11
+    8.453393908382648e-12
+    2.584805818601367e-11
+   -9.269014758400498e-12
+    1.123051218835458e-11
+    2.590186257994186e-11
+    4.782169155689642e-12
+   -9.259134584953882e-12
+     8.42919031435696e-12
+     3.12494911922732e-11
+ 2.461e+11   
+    3.115940747872797e-11
+    8.467631880468765e-12
+    2.579622882415575e-11
+   -9.243851082496015e-12
+    1.121539729019977e-11
+    2.584995518362848e-11
+    4.758503007842827e-12
+    -9.23400390465739e-12
+     8.44355377386644e-12
+    3.118651085538618e-11
+ 2.466e+11   
+    3.109674946441082e-11
+    8.481662718491349e-12
+    2.574478922743741e-11
+   -9.218703654185396e-12
+    1.120011767997051e-11
+    2.579843804425406e-11
+    4.734899814280974e-12
+   -9.208889332924929e-12
+     8.45770957723941e-12
+    3.112378780400834e-11
+ 2.471e+11   
+    3.103434564414056e-11
+    8.495490595982856e-12
+    2.569373098006196e-11
+    -9.19357526555312e-12
+    1.118468063705383e-11
+    2.574730274596823e-11
+     4.71136043615438e-12
+   -9.183793661121043e-12
+      8.4716618983411e-12
+    3.106131933379621e-11
+ 2.476e+11   
+    3.097219339073882e-11
+    8.509119543830086e-12
+    2.564304593020896e-11
+   -9.168468575472147e-12
+    1.116909315293595e-11
+    2.569654113663406e-11
+    4.687885701799487e-12
+     -9.1587195474843e-12
+    8.485414768664741e-12
+    3.099910281647109e-11
+ 2.481e+11   
+    3.091029014996359e-11
+    8.522553457663099e-12
+    2.559272617930226e-11
+   -9.143386115209268e-12
+    1.115336194328326e-11
+    2.564614531711069e-11
+    4.664476407160868e-12
+   -9.133669522727925e-12
+    8.498972084699252e-12
+    3.093713569665919e-11
+ 2.486e+11   
+    3.084863343747267e-11
+    8.535796104837435e-12
+    2.554276407187886e-11
+   -9.118330293793404e-12
+    1.113749345951248e-11
+      2.5596107631136e-11
+    4.641133316136223e-12
+   -9.108645995404078e-12
+    8.512337614891361e-12
+    3.087541548885306e-11
+ 2.491e+11   
+    3.078722083590431e-11
+     8.54885113102558e-12
+    2.549315218602105e-11
+    -9.09330340316135e-12
+    1.112149389987567e-11
+    2.554642065577209e-11
+    4.617857160859863e-12
+   -9.083651257045673e-12
+     8.52551500621773e-12
+    3.081393977448959e-11
+ 2.496e+11   
+    3.072604999206702e-11
+    8.561722066431976e-12
+    2.544388332431478e-11
+   -9.068307623092713e-12
+    1.110536922008333e-11
+    2.549707719237606e-11
+    4.594648641938238e-12
+   -9.058687487097646e-12
+    8.538507790381694e-12
+      3.0752706199137e-11
+ 2.501e+11   
+    3.066511861423596e-11
+    8.574412331647481e-12
+    2.539495050530106e-11
+   -9.043345025946488e-12
+    1.108912514348756e-11
+    2.544807025806331e-11
+    4.571508428650031e-12
+   -9.033756757650486e-12
+    8.551319389650316e-12
+    3.069171246978902e-11
+ 2.506e+11   
+    3.060442446954951e-11
+     8.58692524315752e-12
+    2.534634695538728e-11
+   -9.018417581209668e-12
+    1.107276717084565e-11
+     2.53993930776307e-11
+    4.548437159121207e-12
+   -9.008861037985513e-12
+    8.563953122345969e-12
+    3.063095635225866e-11
+ 2.511e+11   
+    3.054396538150267e-11
+    8.599264018519546e-12
+    2.529806610118954e-11
+   -8.993527159867247e-12
+    1.105630058968307e-11
+    2.535103907590884e-11
+    4.525435440484801e-12
+   -8.984002198942517e-12
+    8.576412208007804e-12
+    3.057043566866914e-11
+ 2.516e+11   
+     3.04837392275329e-11
+    8.611431781223665e-12
+    2.525010156227586e-11
+   -8.968675538603369e-12
+     1.10397304832739e-11
+    2.530300187051708e-11
+    4.502503849033779e-12
+   -8.959182017117664e-12
+    8.588699772238266e-12
+     3.05101482950377e-11
+ 2.521e+11   
+     3.04237439366954e-11
+    8.623431565251946e-12
+    2.520244714428548e-11
+    -8.94386440384073e-12
+    1.102306173925476e-11
+    2.525527526499179e-11
+    4.479642930374465e-12
+   -8.934402178901104e-12
+    8.600818851247932e-12
+    3.045009215894869e-11
+ 2.526e+11   
+    3.036397748742407e-11
+     8.63526631935043e-12
+    2.515509683239795e-11
+   -8.919095355626555e-12
+    1.100629905788838e-11
+    2.520785324226546e-11
+    4.456853199586247e-12
+   -8.909664284360267e-12
+    8.612772396114795e-12
+    3.039026523731279e-11
+ 2.531e+11   
+    3.030443790537533e-11
+    8.646938911027598e-12
+    2.510804478512909e-11
+   -8.894369911371641e-12
+    1.098944695999116e-11
+    2.516072995847196e-11
+    4.434135141393627e-12
+   -8.884969850976941e-12
+    8.624563276770428e-12
+    3.033066555420898e-11
+ 2.536e+11   
+    3.024512326135174e-11
+    8.658452130294225e-12
+    2.506128532843163e-11
+   -8.869689509448646e-12
+    1.097250979453817e-11
+    2.511389973705642e-11
+    4.411489210354166e-12
+   -8.860320317243534e-12
+    8.636194285728801e-12
+    3.027129117880766e-11
+ 2.541e+11   
+    3.018603166930398e-11
+    8.669808693157252e-12
+    2.501481295008063e-11
+    -8.84505551265569e-12
+    1.095549174595913e-11
+    2.506735706316895e-11
+    4.388915831067427e-12
+   -8.835717046124646e-12
+    8.647668141569306e-12
+    3.021214022337067e-11
+ 2.546e+11   
+     3.01271612844071e-11
+    8.681011244881925e-12
+    2.496862229432357e-11
+   -8.820469211550071e-12
+    1.093839684113635e-11
+    2.502109657832314e-11
+     4.36641539840635e-12
+    -8.81116132838909e-12
+    8.658987492189211e-12
+    3.015321084132727e-11
+ 2.551e+11   
+    3.006851030121024e-11
+    8.692062363034684e-12
+    2.492270815677766e-11
+   -8.795931827657278e-12
+    1.092122895611737e-11
+    2.497511307530173e-11
+    4.343988277774901e-12
+    -8.78665438581717e-12
+    8.670154917837927e-12
+    3.009450122542387e-11
+ 2.556e+11   
+     3.00100769518578e-11
+    8.702964560319628e-12
+     2.48770654795576e-11
+   -8.771444516560108e-12
+    1.090399182255181e-11
+    2.492940149329223e-11
+    4.321634805392905e-12
+   -8.762197374287996e-12
+    8.681172933944921e-12
+    3.003600960594454e-11
+ 2.561e+11   
+    2.995185950437921e-11
+    8.713720287221517e-12
+    2.483168934661841e-11
+   -8.747008370871045e-12
+    1.088668903386357e-11
+    2.488395691323704e-11
+    4.299355288609629e-12
+   -8.737791386750476e-12
+    8.692043993755337e-12
+     2.99777342490014e-11
+ 2.566e+11   
+    2.989385626104662e-11
+    8.724331934466435e-12
+     2.47865749792976e-11
+   -8.722624423092659e-12
+     1.08693240511672e-11
+    2.483877455338337e-11
+    4.277150006247361e-12
+   -8.713437456081863e-12
+    8.702770490784012e-12
+    2.991967345489278e-11
+ 2.571e+11   
+    2.983606555679856e-11
+    8.734801835312589e-12
+    2.474171773204519e-11
+   -8.698293648369288e-12
+    1.085190020893838e-11
+    2.479384976502016e-11
+    4.255019208974703e-12
+   -8.689136557838307e-12
+    8.713354761099831e-12
+    2.986182555652779e-11
+ 2.576e+11   
+     2.97784857577281e-11
+      8.7451322676819e-12
+    2.469711308832652e-11
+   -8.674016967133078e-12
+    1.083442072044666e-11
+    2.474917802838809e-11
+      4.2329631197106e-12
+   -8.664889612898968e-12
+    8.723799085452057e-12
+    2.980418891791539e-11
+ 2.581e+11   
+    2.972111525963384e-11
+    8.755325456143676e-12
+    2.465275665668834e-11
+   -8.649795247647899e-12
+    1.081688868295897e-11
+    2.470475494875214e-11
+     4.21098193405793e-12
+   -8.640697490008838e-12
+    8.734105691248964e-12
+    2.974676193271717e-11
+ 2.586e+11   
+    2.966395248663292e-11
+    8.765383573760684e-12
+    2.460864416697573e-11
+   -8.625629308453631e-12
+    1.079930708272156e-11
+    2.466057625262506e-11
+     4.18907582076682e-12
+   -8.616561008221544e-12
+    8.744276754399579e-12
+     2.96895430228619e-11
+ 2.591e+11   
+    2.960699588983449e-11
+    8.775308743807479e-12
+     2.45647714666904e-11
+   -8.601519920713872e-12
+    1.078167879972862e-11
+    2.461663778413201e-11
+    4.167244922227093e-12
+   -8.592480939245468e-12
+    8.754314401028148e-12
+    2.963253063722069e-11
+ 2.596e+11   
+     2.95502439460723e-11
+    8.785103041371181e-12
+    2.452113451748095e-11
+   -8.577467810469567e-12
+    1.076400661228374e-11
+    2.457293550150697e-11
+    4.145489354987823e-12
+   -8.568458009696251e-12
+    8.764220709071649e-12
+    2.957572325034217e-11
+ 2.601e+11   
+     2.94936951566958e-11
+    8.794768494843014e-12
+    2.447772939175632e-11
+   -8.553473660801387e-12
+    1.074629320136207e-11
+    2.452946547371184e-11
+    4.123809210304195e-12
+   -8.544492903257674e-12
+    8.773997709768418e-12
+     2.95191193612456e-11
+ 2.606e+11   
+    2.943734804641781e-11
+    8.804307087310673e-12
+    2.443455226941467e-11
+   -8.529538113901838e-12
+    1.072854115478005e-11
+    2.448622387717097e-11
+    4.102204554710022e-12
+   -8.520586262752534e-12
+     8.78364738904802e-12
+    2.946271749227125e-11
+ 2.611e+11   
+    2.938120116221855e-11
+    8.813720757858533e-12
+    2.439159943467945e-11
+   -8.505661773061824e-12
+    1.071075297117784e-11
+    2.444320699261292e-11
+    4.080675430613568e-12
+   -8.496738692127713e-12
+    8.793171688829779e-12
+    2.940651618798722e-11
+ 2.616e+11   
+    2.932525307230446e-11
+     8.82301140278502e-12
+     2.43488672730369e-11
+   -8.481845204571184e-12
+    1.069293106382199e-11
+    2.440041120201268e-11
+    4.059221856916883e-12
+   -8.472950758353585e-12
+    8.802572508237971e-12
+    2.935051401415076e-11
+ 2.621e+11   
+    2.926950236512041e-11
+    8.832180876743433e-12
+    2.430635226826807e-11
+   -8.458088939537378e-12
+    1.067507776423426e-11
+    2.435783298562894e-11
+    4.037843829655485e-12
+   -8.449222993241522e-12
+    8.811851704741668e-12
+     2.92947095567241e-11
+ 2.626e+11   
+    2.921394764841562e-11
+    8.841230993814513e-12
+     2.42640509995692e-11
+    -8.43439347562328e-12
+    1.065719532565123e-11
+    2.431546891912912e-11
+    4.016541322657911e-12
+   -8.425555895179993e-12
+    8.821011095226428e-12
+    2.923910142094286e-11
+ 2.631e+11   
+    2.915858754836028e-11
+    8.850163528516671e-12
+     2.42219601387558e-11
+   -8.410759278706134e-12
+    1.063928592632212e-11
+     2.42733156707979e-11
+    3.995314288223205e-12
+   -8.401949930792791e-12
+    8.830052457003428e-12
+    2.918368823043625e-11
+ 2.636e+11   
+    2.910342070871387e-11
+    8.858980216760865e-12
+    2.418007644754491e-11
+   -8.387186784460457e-12
+    1.062135167264858e-11
+    2.423136999882379e-11
+    3.974162657813979e-12
+   -8.378405536520126e-12
+    8.838977528764214e-12
+    2.912846862639811e-11
+ 2.641e+11   
+    2.904844579004255e-11
+    8.867682756755923e-12
+    2.413839677491163e-11
+    -8.36367639986547e-12
+    1.060339460217304e-11
+    2.418962874865937e-11
+    3.953086342764412e-12
+   -8.354923120125505e-12
+    8.847788011485708e-12
+    2.907344126680847e-11
+ 2.646e+11   
+    2.899366146898564e-11
+    8.876272809869571e-12
+    2.409691805451484e-11
+    -8.34022850464047e-12
+    1.058541668642021e-11
+    2.414808885045125e-11
+    3.932085235000811e-12
+   -8.331503062129336e-12
+    8.856485569291081e-12
+    2.901860482570242e-11
+ 2.651e+11   
+    2.893906643756934e-11
+    8.884752001450703e-12
+    2.405563730218892e-11
+   -8.316843452608715e-12
+    1.056741983359664e-11
+    2.410674731653459e-11
+    3.911159207773547e-12
+   -8.308145717171997e-12
+    8.865071830272285e-12
+    2.896395799248771e-11
+ 2.656e+11   
+    2.888465940256759e-11
+    8.893121921618333e-12
+    2.401455161349803e-11
+   -8.293521572992382e-12
+    1.054940589115388e-11
+    2.406560123899143e-11
+    3.890308116398007e-12
+   -8.284851415307318e-12
+    8.873548387279289e-12
+    2.890949947130842e-11
+ 2.661e+11   
+    2.883043908490807e-11
+    8.901384126020724e-12
+    2.397365816134942e-11
+   -8.270263171640135e-12
+    1.053137664821935e-11
+    2.402464778726625e-11
+    3.869531799003949e-12
+   -8.261620463229407e-12
+     8.88191679867967e-12
+    2.885522798045491e-11
+ 2.666e+11   
+    2.877640421912289e-11
+    8.909540136569391e-12
+    2.393295419366268e-11
+   -8.247068532189646e-12
+    1.051333383789984e-11
+    2.398388420583843e-11
+    3.848830077290751e-12
+   -8.238453145433536e-12
+    8.890178589093078e-12
+     2.88011422518168e-11
+ 2.671e+11   
+    2.872255355284262e-11
+    8.917591442152496e-12
+    2.389243703109322e-11
+   -8.223937917165759e-12
+    1.049527913946258e-11
+    2.394330781194784e-11
+    3.828202757287468e-12
+    -8.21534972531392e-12
+     8.89833525010522e-12
+    2.874724103038108e-11
+ 2.676e+11   
+    2.866888584633289e-11
+    8.925539499329942e-12
+    2.385210406480569e-11
+   -8.200871569017379e-12
+    1.047721418039719e-11
+    2.390291599337059e-11
+    3.807649630116601e-12
+   -8.192310446198997e-12
+    8.906388240963568e-12
+    2.869352307377092e-11
+ 2.681e+11   
+    2.861539987207159e-11
+    8.933385733014229e-12
+    2.381195275429747e-11
+   -8.177869711093898e-12
+    1.045914053836501e-11
+    2.386270620624471e-11
+    3.787170472759378e-12
+   -8.169335532326929e-12
+    8.914338989259383e-12
+    2.863998715182656e-11
+ 2.686e+11   
+    2.856209441436726e-11
+    8.941131537140596e-12
+    2.377198062526804e-11
+   -8.154932548563557e-12
+    1.044105974303702e-11
+    2.382267597294071e-11
+    3.766765048821426e-12
+   -8.146425189763104e-12
+    8.922188891597929e-12
+    2.858663204622576e-11
+ 2.691e+11   
+    2.850896826901548e-11
+    8.948778275327498e-12
+    2.373218526753366e-11
+    -8.13206026927507e-12
+     1.04229732778275e-11
+    2.378282287997823e-11
+    3.746433109298193e-12
+   -8.123579607260643e-12
+    8.929939314260328e-12
+    2.853345655014357e-11
+ 2.696e+11   
+     2.84560202429937e-11
+    8.956327281531865e-12
+    2.369256433298571e-11
+   -8.109253044564207e-12
+    1.040488258152576e-11
+    2.374314457598495e-11
+    3.726174393337915e-12
+   -8.100798957066196e-12
+    8.937591593859104e-12
+    2.848045946794929e-11
+ 2.701e+11   
+    2.840324915419263e-11
+    8.963779860699591e-12
+    2.365311553358992e-11
+    -8.08651103000787e-12
+    1.038678904982974e-11
+    2.370363876969714e-11
+    3.705988629001538e-12
+   -8.078083395673112e-12
+    8.945147037989821e-12
+     2.84276396149408e-11
+ 2.706e+11   
+    2.835065383118337e-11
+    8.971137289414487e-12
+    2.361383663942666e-11
+   -8.063834366126213e-12
+    1.036869403678684e-11
+     2.36643032280003e-11
+    3.685875534018397e-12
+   -8.055433064522546e-12
+    8.952606925880416e-12
+    2.837499581711327e-11
+ 2.711e+11   
+    2.829823311301888e-11
+    8.978400816546621e-12
+    2.357472547677016e-11
+    -8.04122317903558e-12
+    1.035059885614425e-11
+    2.362513577400912e-11
+    3.665834816536582e-12
+   -8.032848090655654e-12
+    8.959972509040478e-12
+    2.832252691096332e-11
+ 2.716e+11   
+    2.824598584906861e-11
+     8.98557166390212e-12
+    2.353577992620562e-11
+   -8.018677581053064e-12
+    1.033250478261342e-11
+    2.358613428518449e-11
+     3.64586617586683e-12
+   -8.010328587317404e-12
+    8.967245011911564e-12
+    2.827023174332545e-11
+ 2.721e+11   
+    2.819391089888569e-11
+    8.992651026875324e-12
+    2.349699792078322e-11
+   -7.996197671255432e-12
+    1.031441305305133e-11
+    2.354729669148742e-11
+    3.625969303219175e-12
+    -7.98787465451457e-12
+    8.974425632520029e-12
+    2.821810917124082e-11
+ 2.726e+11   
+    2.814200713210456e-11
+    8.999640075104693e-12
+     2.34583774442084e-11
+   -7.973783535992844e-12
+    1.029632486756357e-11
+    2.350862097356915e-11
+    3.606143882431884e-12
+   -7.965486379528819e-12
+    8.981515543133357e-12
+    2.816615806185662e-11
+ 2.731e+11   
+    2.809027342836876e-11
+    9.006539953133473e-12
+    2.341991652906718e-11
+   -7.951435249359948e-12
+    1.027824139053108e-11
+    2.347010516099544e-11
+     3.58638959069111e-12
+   -7.943163837387445e-12
+    8.988515890920929e-12
+    2.811437729235516e-11
+ 2.736e+11   
+    2.803870867728694e-11
+    9.013351781075194e-12
+     2.33816132550856e-11
+   -7.929152873626077e-12
+      1.0260163751565e-11
+    2.343174733050581e-11
+    3.566706099241064e-12
+   -7.920907091292178e-12
+     8.99542779862079e-12
+    2.806276574991138e-11
+ 2.741e+11   
+    2.798731177841707e-11
+    9.020076655286203e-12
+    2.334346574742367e-11
+   -7.906936459625223e-12
+    1.024209304639264e-11
+    2.339354560430609e-11
+    3.547093074084049e-12
+   -7.898716193009237e-12
+    9.002252365211376e-12
+    2.801132233167766e-11
+ 2.746e+11   
+    2.793608164127582e-11
+    9.026715649043525e-12
+    2.330547217500148e-11
+    -7.88478604710837e-12
+    1.022403033767707e-11
+    2.335549814839323e-11
+     3.52755017666961e-12
+   -7.876591183220888e-12
+    9.008990666590263e-12
+    2.796004594479446e-11
+ 2.751e+11   
+    2.788501718537425e-11
+    9.033269813230606e-12
+    2.326763074885832e-11
+   -7.862701665059555e-12
+     1.02059766557747e-11
+    2.331760317091329e-11
+     3.50807706457201e-12
+   -7.854532091840616e-12
+    9.015643756259726e-12
+    2.790893550642617e-11
+ 2.756e+11   
+    2.783411734027646e-11
+    9.039740177029313e-12
+    2.322993972054395e-11
+   -7.840683331976831e-12
+    1.018793299943291e-11
+     2.32798589205508e-11
+    3.488673392156162e-12
+   -7.832538938294052e-12
+    9.022212666018812e-12
+    2.785798994382069e-11
+ 2.761e+11   
+    2.778338104568178e-11
+    9.046127748619894e-12
+    2.319239738054144e-11
+   -7.818731056119806e-12
+    1.016990033643119e-11
+    2.324226368494954e-11
+    3.469338811231041e-12
+   -7.810611731765947e-12
+    9.028698406663004e-12
+    2.780720819439157e-11
+ 2.766e+11   
+    2.773280725152837e-11
+    9.052433515887343e-12
+    2.315500205672066e-11
+   -7.796844835726177e-12
+    1.015187960416823e-11
+    2.320481578916444e-11
+    3.450072971690314e-12
+   -7.788750471416059e-12
+    9.035101968690484e-12
+     2.77565892058216e-11
+ 2.771e+11   
+    2.768239491811701e-11
+    9.058658447135278e-12
+    2.311775211282298e-11
+   -7.775024659197151e-12
+     1.01338717101981e-11
+    2.316751359414382e-11
+     3.43087552213992e-12
+   -7.766955146564295e-12
+    9.041424323015927e-12
+    2.770613193618693e-11
+ 2.776e+11   
+    2.763214301625526e-11
+    9.064803491806779e-12
+    2.308064594697636e-11
+   -7.753270505254776e-12
+    1.011587753271823e-11
+    2.313035549524211e-11
+    3.411746110512226e-12
+   -7.745225736847744e-12
+    9.047666421690471e-12
+    2.765583535410028e-11
+ 2.781e+11   
+    2.758205052741902e-11
+     9.07086958121169e-12
+    2.304368199024071e-11
+   -7.731582343071357e-12
+    1.009789792101205e-11
+    2.309333992076233e-11
+    3.392684384666724e-12
+   -7.723562212349794e-12
+    9.053829198628669e-12
+     2.76056984388724e-11
+ 2.786e+11   
+    2.753211644393164e-11
+    9.076857629259855e-12
+     2.30068587051819e-11
+   -7.709960132373705e-12
+    1.007993369584741e-11
+    2.305646533052815e-11
+    3.373689992976707e-12
+     -7.7019645337038e-12
+    9.059913570341435e-12
+    2.755572018069058e-11
+ 2.791e+11   
+    2.748233976915956e-11
+    9.082768533201083e-12
+    2.297017458447715e-11
+    -7.68840382352226e-12
+    1.006198564983586e-11
+    2.301973021448534e-11
+     3.35476258490183e-12
+   -7.680432652172471e-12
+    9.065920436674453e-12
+    2.750589958081287e-11
+ 2.796e+11   
+    2.743271951772243e-11
+    9.088603174369522e-12
+    2.293362814954827e-11
+   -7.666913357567495e-12
+    1.004405454775318e-11
+    2.298313309133307e-11
+     3.33590181154686e-12
+   -7.658966509703365e-12
+    9.071850681552938e-12
+    2.745623565177805e-11
+ 2.801e+11   
+    2.738325471571812e-11
+    9.094362418933971e-12
+    2.289721794922427e-11
+   -7.645488666284376e-12
+    1.002614112682341e-11
+    2.294667250718267e-11
+     3.31710732620574e-12
+   -7.637566038963775e-12
+    9.077705173729838e-12
+    2.740672741762859e-11
+ 2.806e+11   
+     2.73339444009598e-11
+    9.100047118651578e-12
+    2.286094255843296e-11
+   -7.624129672186169e-12
+    1.000824609697029e-11
+    2.291034703424583e-11
+    3.298378784891879e-12
+   -7.616231163354208e-12
+    9.083484767538904e-12
+    2.735737391414666e-11
+ 2.811e+11   
+    2.728478762322582e-11
+    9.105658111625439e-12
+      2.2824800576921e-11
+   -7.602836288519842e-12
+    9.990370141037045e-12
+    2.287415526955228e-11
+    3.279715846853531e-12
+   -7.594961797003066e-12
+    9.089190303651933e-12
+    2.730817418910288e-11
+ 2.816e+11   
+    2.723578344452048e-11
+    9.111196223066208e-12
+    2.278879062800223e-11
+   -7.581608419242364e-12
+    9.972513914976277e-12
+    2.283809583369342e-11
+     3.26111817507501e-12
+   -7.573757844743841e-12
+    9.094822609837966e-12
+    2.725912730251489e-11
+ 2.821e+11   
+    2.718693093934477e-11
+     9.11666226605499e-12
+    2.275291135733438e-11
+   -7.560445958981036e-12
+    9.954678048013609e-12
+     2.28021673695961e-11
+    3.242585436763863e-12
+   -7.552619202074581e-12
+    9.100382501725609e-12
+    2.721023232691645e-11
+ 2.826e+11   
+     2.71382291949762e-11
+    9.122057042308272e-12
+    2.271716143172352e-11
+   -7.539348792978394e-12
+    9.936863142785462e-12
+    2.276636854132357e-11
+    3.224117303823183e-12
+   -7.531545755102888e-12
+    9.105870783566807e-12
+    2.716148834763563e-11
+ 2.831e+11   
+    2.708967731175744e-11
+    9.127381342944698e-12
+     2.26815395379565e-11
+   -7.518316797021849e-12
+    9.919069775453553e-12
+    2.273069803290355e-11
+    3.205713453310291e-12
+   -7.510537380475791e-12
+     9.11128824900137e-12
+    2.711289446308063e-11
+ 2.836e+11   
+    2.704127440339142e-11
+    9.132635949250881e-12
+     2.26460443816608e-11
+    -7.49734983736117e-12
+    9.901298495797953e-12
+    2.269515454718471e-11
+    3.187373567880683e-12
+   -7.489593945296959e-12
+    9.116635681822068e-12
+    2.706444978503359e-11
+ 2.841e+11   
+    2.699301959724387e-11
+    9.137821633447962e-12
+    2.261067468619189e-11
+   -7.476447770612809e-12
+     9.88354982729068e-12
+    2.265973680472017e-11
+    3.169097336218472e-12
+    -7.46871530703103e-12
+    9.121913856739182e-12
+    2.701615343895003e-11
+ 2.846e+11   
+    2.694491203465055e-11
+    9.142939159456258e-12
+    2.257542919154783e-11
+   -7.455610443653536e-12
+     9.86582426715086e-12
+    2.262444354267807e-11
+    3.150884453452543e-12
+   -7.447901313397417e-12
+    9.127123540143796e-12
+    2.696800456426429e-11
+ 2.851e+11   
+    2.689695087122993e-11
+    9.147989283658488e-12
+     2.25403066533106e-11
+   -7.434837693503897e-12
+    9.848122286383502e-12
+    2.258927351377874e-11
+    3.132734621559009e-12
+   -7.427151802253753e-12
+    9.132265490868877e-12
+    2.692000231469907e-11
+ 2.856e+11   
+    2.684913527719991e-11
+    9.152972755660031e-12
+    2.250530584161507e-11
+   -7.414129347202609e-12
+    9.830444329804049e-12
+    2.255422548526013e-11
+    3.114647549750339e-12
+   -7.406466601470193e-12
+    9.137340460948532e-12
+    2.687214585858021e-11
+ 2.861e+11   
+    2.680146443769733e-11
+    9.157890319046536e-12
+     2.24704255401435e-11
+    -7.39348522167221e-12
+    9.812790816048692e-12
+    2.251929823786756e-11
+    3.096622954850469e-12
+   -7.385845528795528e-12
+    9.142349196372702e-12
+    2.682443437915262e-11
+ 2.866e+11   
+    2.675393755309997e-11
+    9.162742712136076e-12
+    2.243566454514699e-11
+   -7.372905123578505e-12
+    9.795162137573544e-12
+    2.248449056487229e-11
+    3.078660561657144e-12
+   -7.365288391716076e-12
+    9.147292437838806e-12
+    2.677686707490031e-11
+ 2.871e+11   
+    2.670655383935095e-11
+    9.167530668728403e-12
+    2.240102166449396e-11
+   -7.352388849182235e-12
+    9.777558660643151e-12
+    2.244980127111447e-11
+    3.060760103290898e-12
+   -7.344794987308294e-12
+    9.152170921497804e-12
+    2.672944315986734e-11
+ 2.876e+11   
+    2.665931252828305e-11
+    9.172254918846687e-12
+    2.236649571674314e-11
+   -7.331936184186703e-12
+    9.759980725309663e-12
+    2.241522917207329e-11
+    3.042921321531054e-12
+   -7.324365102085602e-12
+    9.156985379695146e-12
+    2.668216186397959e-11
+ 2.881e+11   
+    2.661221286794466e-11
+    9.176916189474813e-12
+    2.233208553024361e-11
+   -7.311546903579359e-12
+    9.742428645384266e-12
+    2.238077309296215e-11
+    3.025143967139301e-12
+   -7.303998511841051e-12
+    9.161736541705076e-12
+     2.66350224333674e-11
+ 2.886e+11   
+    2.656525412292418e-11
+    9.181515205286395e-12
+    2.229778994226016e-11
+   -7.291220771470431e-12
+    9.724902708402185e-12
+    2.234643186785057e-11
+    3.007427800170484e-12
+   -7.283694981485367e-12
+    9.166425134458592e-12
+    2.658802413068725e-11
+ 2.891e+11   
+    2.651843557467444e-11
+    9.186052689367201e-12
+    2.226360779812337e-11
+   -7.270957540928045e-12
+    9.707403175581371e-12
+    2.231220433880995e-11
+    2.989772590271072e-12
+   -7.263454264882334e-12
+    9.171051883263196e-12
+    2.654116623544255e-11
+ 2.896e+11   
+    2.647175652183467e-11
+    9.190529363928623e-12
+    2.222953795040636e-11
+   -7.250756953810865e-12
+    9.689930281778046e-12
+    2.227808935508618e-11
+    2.972178116965723e-12
+   -7.243276104681974e-12
+    9.175617512514803e-12
+    2.649444804430328e-11
+ 2.901e+11   
+    2.642521628055121e-11
+    9.194945951012871e-12
+    2.219557925812477e-11
+   -7.230618740599261e-12
+    9.672484235437246e-12
+    2.224408577229569e-11
+    2.954644169931803e-12
+   -7.223160232151702e-12
+    9.180122746400329e-12
+    2.644786887142273e-11
+ 2.906e+11   
+    2.637881418479499e-11
+     9.19930317318821e-12
+    2.216173058596268e-11
+   -7.210542620225692e-12
+    9.655065218542714e-12
+    2.221019245164803e-11
+    2.937170549262093e-12
+   -7.203106367006324e-12
+    9.184568309591674e-12
+    2.640142804875213e-11
+ 2.911e+11   
+    2.633254958667541e-11
+     9.20360175423465e-12
+    2.212799080352291e-11
+   -7.190528299903785e-12
+    9.637673386564037e-12
+    2.217640825919128e-11
+    2.919757065716131e-12
+    -7.18311421723842e-12
+    9.188954927928582e-12
+    2.635512492635151e-11
+ 2.916e+11   
+     2.62864218567509e-11
+    9.207842419818099e-12
+    2.209435878460043e-11
+   -7.170575474959301e-12
+    9.620308868403599e-12
+    2.214273206508268e-11
+    2.902403540960058e-12
+   -7.163183478948145e-12
+    9.193283329091703e-12
+    2.630895887269698e-11
+ 2.921e+11   
+    2.624043038433537e-11
+    9.212025898154579e-12
+    2.206083340648189e-11
+   -7.150683828660287e-12
+    9.602971766344539e-12
+    2.210916274288338e-11
+    2.885109807795706e-12
+   -7.143313836174894e-12
+    9.197554243263457e-12
+    2.626292927498352e-11
+ 2.926e+11   
+    2.619457457779906e-11
+    9.216152920661534e-12
+    2.202741354926654e-11
+   -7.130853032050088e-12
+    9.585662155998351e-12
+    2.207569916887622e-11
+    2.867875710377991e-12
+    -7.12350496072958e-12
+     9.20176840377847e-12
+    2.621703553942321e-11
+ 2.931e+11   
+    2.614885386486487e-11
+    9.220224222597503e-12
+    2.199409809521228e-11
+   -7.111082743781654e-12
+    9.568380086255678e-12
+    2.204234022140833e-11
+    2.850701104422363e-12
+   -7.103756512029184e-12
+    9.205926547760874e-12
+    2.617127709153783e-11
+ 2.936e+11   
+    2.610326769289813e-11
+     9.22424054368901e-12
+    2.196088592810457e-11
+   -7.091372609954702e-12
+     9.55112557923911e-12
+      2.2009084780256e-11
+    2.833585857400421e-12
+   -7.084068136934672e-12
+    9.210029416749057e-12
+    2.612565337644605e-11
+ 2.941e+11   
+     2.60578155291912e-11
+    9.228202628744051e-12
+    2.192777593264777e-11
+   -7.071722263955948e-12
+    9.533898630258776e-12
+    2.197593172601254e-11
+    2.816529848726389e-12
+   -7.064439469590825e-12
+    9.214077757307415e-12
+    2.608016385914431e-11
+ 2.946e+11   
+    2.601249686124065e-11
+     9.23211122825213e-12
+    2.189476699388011e-11
+   -7.052131326303027e-12
+    9.516699207772707e-12
+    2.194287993950047e-11
+     2.79953296993191e-12
+   -7.044870131270553e-12
+    9.218072321624421e-12
+    2.603480802478126e-11
+ 2.951e+11   
+    2.596731119701811e-11
+    9.235967098970572e-12
+    2.186185799661018e-11
+   -7.032599404492488e-12
+    9.499527253350323e-12
+    2.190992830120402e-11
+    2.782595124830916e-12
+   -7.025359730223147e-12
+    9.222013868096832e-12
+     2.59895853789251e-11
+ 2.956e+11   
+    2.592225806523265e-11
+    9.239771004495457e-12
+    2.182904782487646e-11
+   -7.013126092852281e-12
+    9.482382681641993e-12
+    2.187707569072547e-11
+    2.765716229674498e-12
+   -7.005907861526921e-12
+    9.225903161898995e-12
+     2.59444954478235e-11
+ 2.961e+11   
+    2.587733701558704e-11
+    9.243523715818952e-12
+    2.179633536142799e-11
+    -6.99371097239964e-12
+    9.465265380353449e-12
+     2.18443209862638e-11
+    2.748896213294814e-12
+   -6.986514106946677e-12
+    9.229740975538664e-12
+    2.589953777865607e-11
+ 2.966e+11   
+    2.583254761902439e-11
+    9.247226011871144e-12
+    2.176371948722732e-11
+   -6.974353610703796e-12
+    9.448175210225392e-12
+    2.181166306411282e-11
+    2.732135017239172e-12
+   -6.967178034797673e-12
+    9.233528089396177e-12
+    2.585471193977867e-11
+ 2.971e+11   
+    2.578788946796676e-11
+    9.250878680045669e-12
+    2.173119908097455e-11
+   -6.955053561755436e-12
+    9.431112005021009e-12
+    2.177910079818397e-11
+    2.715432595893679e-12
+   -6.947899199814404e-12
+    9.237265292249436e-12
+    2.581001752095935e-11
+ 2.976e+11   
+    2.574336217654574e-11
+    9.254482516711121e-12
+    2.169877301865216e-11
+   -6.935810365841757e-12
+      9.4140755715181e-12
+    2.174663305954741e-11
+    2.698788916596609e-12
+   -6.928677143025829e-12
+    9.240953381782788e-12
+    2.576545413360479e-11
+ 2.981e+11   
+    2.569896538082227e-11
+    9.258038327705094e-12
+     2.16664401730917e-11
+    -6.91662354942899e-12
+    9.397065689509982e-12
+    2.171425871599668e-11
+    2.682203959740668e-12
+   -6.909511391638468e-12
+    9.244593165080366e-12
+    2.572102141097936e-11
+ 2.986e+11   
+    2.565469873899884e-11
+    9.261546928813442e-12
+    2.163419941355963e-11
+   -6.897492625051352e-12
+    9.380082111811887e-12
+    2.168197663163119e-11
+    2.665677718865415e-12
+   -6.890401458925175e-12
+    9.248185459102549e-12
+    2.567671900841235e-11
+ 2.991e+11   
+    2.561056193162022e-11
+    9.265009146231734e-12
+    2.160204960536463e-11
+   -6.878417091208407e-12
+    9.363124564276412e-12
+    2.164978566646235e-11
+    2.649210200738284e-12
+   -6.871346844122526e-12
+    9.251731091147577e-12
+    2.563254660349839e-11
+ 2.996e+11   
+    2.556655466176534e-11
+    9.268425817011095e-12
+    2.156998960948431e-11
+   -6.859396432269608e-12
+     9.34619274581565e-12
+    2.161768467603702e-11
+    2.632801425425317e-12
+   -6.852347032335529e-12
+    9.255230899294873e-12
+    2.558850389628505e-11
* NOTE: Solution at 1e+08 Hz used as DC point.

.ends
