* BEGIN ANSOFT HEADER
* node 1    trace_p_0_T1
* node 2    trace_n_0_T1
* node 3    trace_p_1_T1
* node 4    trace_n_1_T1
* node 5    trace_p_0_T2
* node 6    trace_n_0_T2
* node 7    trace_p_1_T2
* node 8    trace_n_1_T2
*   Format: HSPICE
*   Topckt: m4lines_HFSS_fws
*     Date: Sat Jun 06 10:16:42 2020
*    Notes: Frequency range: 1e+08 to 7e+10 Hz, 700 points
*         : Maximum number of poles: 10000
*         : S-Matrix fitting error tolerance: 0.001
*         : Causality check tolerance: auto
*         : Passivity enforcement: on (by iterated fitting)
*         : Causality enforcement: off
*         : Fitting method: FastFit
*         : Matrix fitting: By entire matrix (required by FastFit)
*         : Ensure Z-parameter accuracy: on
*         : Relative error control: off
*         : Common ground option: on
*         : Final fitting error: 0.00384938
*         : Final model order: 328
* END ANSOFT HEADER

.subckt m4lines_HFSS_fws 1 2 3 4 5 6 7 8
Vam1 1 n2 dc 0
Rport1 n2 0 50 noise=0
Vam2 2 n4 dc 0
Rport2 n4 0 50 noise=0
Vam3 3 n6 dc 0
Rport3 n6 0 50 noise=0
Vam4 4 n8 dc 0
Rport4 n8 0 50 noise=0
Vam5 5 n10 dc 0
Rport5 n10 0 50 noise=0
Vam6 6 n12 dc 0
Rport6 n12 0 50 noise=0
Vam7 7 n14 dc 0
Rport7 n14 0 50 noise=0
Vam8 8 n16 dc 0
Rport8 n16 0 50 noise=0

Fi1 0 ni1 Vam1 50
Gi1 0 ni1 1 0 1
Rt1 ni1 0 1 noise=0
Fi2 0 ni2 Vam2 50
Gi2 0 ni2 2 0 1
Rt2 ni2 0 1 noise=0
Fi3 0 ni3 Vam3 50
Gi3 0 ni3 3 0 1
Rt3 ni3 0 1 noise=0
Fi4 0 ni4 Vam4 50
Gi4 0 ni4 4 0 1
Rt4 ni4 0 1 noise=0
Fi5 0 ni5 Vam5 50
Gi5 0 ni5 5 0 1
Rt5 ni5 0 1 noise=0
Fi6 0 ni6 Vam6 50
Gi6 0 ni6 6 0 1
Rt6 ni6 0 1 noise=0
Fi7 0 ni7 Vam7 50
Gi7 0 ni7 7 0 1
Rt7 ni7 0 1 noise=0
Fi8 0 ni8 Vam8 50
Gi8 0 ni8 8 0 1
Rt8 ni8 0 1 noise=0

Ca1 ns1 0 1e-12
Ra1 ns1 0 0.0599459941272 noise=0
Ca2 ns2 0 1e-12
Ra2 ns2 0 0.714606679535 noise=0
Ca3 ns3 0 1e-12
Ra3 ns3 0 1.19287160881 noise=0
Ca4 ns4 0 1e-12
Ca5 ns5 0 1e-12
Ra4 ns4 0 26.828727021 noise=0
Ra5 ns5 0 26.828727021 noise=0
Ga4 ns4 0 ns5 0 -0.518048785893
Ga5 ns5 0 ns4 0 0.518048785893
Ca6 ns6 0 1e-12
Ca7 ns7 0 1e-12
Ra6 ns6 0 90.0406412861 noise=0
Ra7 ns7 0 90.0406412861 noise=0
Ga6 ns6 0 ns7 0 -0.487119257249
Ga7 ns7 0 ns6 0 0.487119257249
Ca8 ns8 0 1e-12
Ca9 ns9 0 1e-12
Ra8 ns8 0 29.4872472308 noise=0
Ra9 ns9 0 29.4872472308 noise=0
Ga8 ns8 0 ns9 0 -0.46382169076
Ga9 ns9 0 ns8 0 0.46382169076
Ca10 ns10 0 1e-12
Ca11 ns11 0 1e-12
Ra10 ns10 0 31.4880587202 noise=0
Ra11 ns11 0 31.4880587202 noise=0
Ga10 ns10 0 ns11 0 -0.426117672518
Ga11 ns11 0 ns10 0 0.426117672518
Ca12 ns12 0 1e-12
Ca13 ns13 0 1e-12
Ra12 ns12 0 19.1952084606 noise=0
Ra13 ns13 0 19.1952084606 noise=0
Ga12 ns12 0 ns13 0 -0.398679757461
Ga13 ns13 0 ns12 0 0.398679757461
Ca14 ns14 0 1e-12
Ca15 ns15 0 1e-12
Ra14 ns14 0 38.9735617239 noise=0
Ra15 ns15 0 38.9735617239 noise=0
Ga14 ns14 0 ns15 0 -0.385574664967
Ga15 ns15 0 ns14 0 0.385574664967
Ca16 ns16 0 1e-12
Ca17 ns17 0 1e-12
Ra16 ns16 0 23.3700179636 noise=0
Ra17 ns17 0 23.3700179636 noise=0
Ga16 ns16 0 ns17 0 -0.32363874977
Ga17 ns17 0 ns16 0 0.32363874977
Ca18 ns18 0 1e-12
Ca19 ns19 0 1e-12
Ra18 ns18 0 13.6366308475 noise=0
Ra19 ns19 0 13.6366308475 noise=0
Ga18 ns18 0 ns19 0 -0.2818027486
Ga19 ns19 0 ns18 0 0.2818027486
Ca20 ns20 0 1e-12
Ca21 ns21 0 1e-12
Ra20 ns20 0 36.4720266288 noise=0
Ra21 ns21 0 36.4720266288 noise=0
Ga20 ns20 0 ns21 0 -0.291418716466
Ga21 ns21 0 ns20 0 0.291418716466
Ca22 ns22 0 1e-12
Ca23 ns23 0 1e-12
Ra22 ns22 0 22.570362028 noise=0
Ra23 ns23 0 22.570362028 noise=0
Ga22 ns22 0 ns23 0 -0.219789949348
Ga23 ns23 0 ns22 0 0.219789949348
Ca24 ns24 0 1e-12
Ca25 ns25 0 1e-12
Ra24 ns24 0 35.3564229023 noise=0
Ra25 ns25 0 35.3564229023 noise=0
Ga24 ns24 0 ns25 0 -0.196387080388
Ga25 ns25 0 ns24 0 0.196387080388
Ca26 ns26 0 1e-12
Ca27 ns27 0 1e-12
Ra26 ns26 0 19.3225792178 noise=0
Ra27 ns27 0 19.3225792178 noise=0
Ga26 ns26 0 ns27 0 -0.158984338989
Ga27 ns27 0 ns26 0 0.158984338989
Ca28 ns28 0 1e-12
Ca29 ns29 0 1e-12
Ra28 ns28 0 22.3171225035 noise=0
Ra29 ns29 0 22.3171225035 noise=0
Ga28 ns28 0 ns29 0 -0.112121022154
Ga29 ns29 0 ns28 0 0.112121022154
Ca30 ns30 0 1e-12
Ca31 ns31 0 1e-12
Ra30 ns30 0 35.6994407039 noise=0
Ra31 ns31 0 35.6994407039 noise=0
Ga30 ns30 0 ns31 0 -0.097312790312
Ga31 ns31 0 ns30 0 0.097312790312
Ca32 ns32 0 1e-12
Ca33 ns33 0 1e-12
Ra32 ns32 0 21.0761624353 noise=0
Ra33 ns33 0 21.0761624353 noise=0
Ga32 ns32 0 ns33 0 -0.0785079694625
Ga33 ns33 0 ns32 0 0.0785079694625
Ca34 ns34 0 1e-12
Ca35 ns35 0 1e-12
Ra34 ns34 0 6461.79173097 noise=0
Ra35 ns35 0 6461.79173097 noise=0
Ga34 ns34 0 ns35 0 -0.0625345296116
Ga35 ns35 0 ns34 0 0.0625345296116
Ca36 ns36 0 1e-12
Ca37 ns37 0 1e-12
Ra36 ns36 0 26.8817745081 noise=0
Ra37 ns37 0 26.8817745081 noise=0
Ga36 ns36 0 ns37 0 -0.016065358588
Ga37 ns37 0 ns36 0 0.016065358588
Ca38 ns38 0 1e-12
Ra38 ns38 0 30.8646103733 noise=0
Ca39 ns39 0 1e-12
Ra39 ns39 0 24137.9690629 noise=0
Ca40 ns40 0 1e-12
Ca41 ns41 0 1e-12
Ra40 ns40 0 3536.160082 noise=0
Ra41 ns41 0 3536.160082 noise=0
Ga40 ns40 0 ns41 0 -0.000237869767882
Ga41 ns41 0 ns40 0 0.000237869767882
Ca42 ns42 0 1e-12
Ra42 ns42 0 0.0599459941272 noise=0
Ca43 ns43 0 1e-12
Ra43 ns43 0 0.714606679535 noise=0
Ca44 ns44 0 1e-12
Ra44 ns44 0 1.19287160881 noise=0
Ca45 ns45 0 1e-12
Ca46 ns46 0 1e-12
Ra45 ns45 0 26.828727021 noise=0
Ra46 ns46 0 26.828727021 noise=0
Ga45 ns45 0 ns46 0 -0.518048785893
Ga46 ns46 0 ns45 0 0.518048785893
Ca47 ns47 0 1e-12
Ca48 ns48 0 1e-12
Ra47 ns47 0 90.0406412861 noise=0
Ra48 ns48 0 90.0406412861 noise=0
Ga47 ns47 0 ns48 0 -0.487119257249
Ga48 ns48 0 ns47 0 0.487119257249
Ca49 ns49 0 1e-12
Ca50 ns50 0 1e-12
Ra49 ns49 0 29.4872472308 noise=0
Ra50 ns50 0 29.4872472308 noise=0
Ga49 ns49 0 ns50 0 -0.46382169076
Ga50 ns50 0 ns49 0 0.46382169076
Ca51 ns51 0 1e-12
Ca52 ns52 0 1e-12
Ra51 ns51 0 31.4880587202 noise=0
Ra52 ns52 0 31.4880587202 noise=0
Ga51 ns51 0 ns52 0 -0.426117672518
Ga52 ns52 0 ns51 0 0.426117672518
Ca53 ns53 0 1e-12
Ca54 ns54 0 1e-12
Ra53 ns53 0 19.1952084606 noise=0
Ra54 ns54 0 19.1952084606 noise=0
Ga53 ns53 0 ns54 0 -0.398679757461
Ga54 ns54 0 ns53 0 0.398679757461
Ca55 ns55 0 1e-12
Ca56 ns56 0 1e-12
Ra55 ns55 0 38.9735617239 noise=0
Ra56 ns56 0 38.9735617239 noise=0
Ga55 ns55 0 ns56 0 -0.385574664967
Ga56 ns56 0 ns55 0 0.385574664967
Ca57 ns57 0 1e-12
Ca58 ns58 0 1e-12
Ra57 ns57 0 23.3700179636 noise=0
Ra58 ns58 0 23.3700179636 noise=0
Ga57 ns57 0 ns58 0 -0.32363874977
Ga58 ns58 0 ns57 0 0.32363874977
Ca59 ns59 0 1e-12
Ca60 ns60 0 1e-12
Ra59 ns59 0 13.6366308475 noise=0
Ra60 ns60 0 13.6366308475 noise=0
Ga59 ns59 0 ns60 0 -0.2818027486
Ga60 ns60 0 ns59 0 0.2818027486
Ca61 ns61 0 1e-12
Ca62 ns62 0 1e-12
Ra61 ns61 0 36.4720266288 noise=0
Ra62 ns62 0 36.4720266288 noise=0
Ga61 ns61 0 ns62 0 -0.291418716466
Ga62 ns62 0 ns61 0 0.291418716466
Ca63 ns63 0 1e-12
Ca64 ns64 0 1e-12
Ra63 ns63 0 22.570362028 noise=0
Ra64 ns64 0 22.570362028 noise=0
Ga63 ns63 0 ns64 0 -0.219789949348
Ga64 ns64 0 ns63 0 0.219789949348
Ca65 ns65 0 1e-12
Ca66 ns66 0 1e-12
Ra65 ns65 0 35.3564229023 noise=0
Ra66 ns66 0 35.3564229023 noise=0
Ga65 ns65 0 ns66 0 -0.196387080388
Ga66 ns66 0 ns65 0 0.196387080388
Ca67 ns67 0 1e-12
Ca68 ns68 0 1e-12
Ra67 ns67 0 19.3225792178 noise=0
Ra68 ns68 0 19.3225792178 noise=0
Ga67 ns67 0 ns68 0 -0.158984338989
Ga68 ns68 0 ns67 0 0.158984338989
Ca69 ns69 0 1e-12
Ca70 ns70 0 1e-12
Ra69 ns69 0 22.3171225035 noise=0
Ra70 ns70 0 22.3171225035 noise=0
Ga69 ns69 0 ns70 0 -0.112121022154
Ga70 ns70 0 ns69 0 0.112121022154
Ca71 ns71 0 1e-12
Ca72 ns72 0 1e-12
Ra71 ns71 0 35.6994407039 noise=0
Ra72 ns72 0 35.6994407039 noise=0
Ga71 ns71 0 ns72 0 -0.097312790312
Ga72 ns72 0 ns71 0 0.097312790312
Ca73 ns73 0 1e-12
Ca74 ns74 0 1e-12
Ra73 ns73 0 21.0761624353 noise=0
Ra74 ns74 0 21.0761624353 noise=0
Ga73 ns73 0 ns74 0 -0.0785079694625
Ga74 ns74 0 ns73 0 0.0785079694625
Ca75 ns75 0 1e-12
Ca76 ns76 0 1e-12
Ra75 ns75 0 6461.79173097 noise=0
Ra76 ns76 0 6461.79173097 noise=0
Ga75 ns75 0 ns76 0 -0.0625345296116
Ga76 ns76 0 ns75 0 0.0625345296116
Ca77 ns77 0 1e-12
Ca78 ns78 0 1e-12
Ra77 ns77 0 26.8817745081 noise=0
Ra78 ns78 0 26.8817745081 noise=0
Ga77 ns77 0 ns78 0 -0.016065358588
Ga78 ns78 0 ns77 0 0.016065358588
Ca79 ns79 0 1e-12
Ra79 ns79 0 30.8646103733 noise=0
Ca80 ns80 0 1e-12
Ra80 ns80 0 24137.9690629 noise=0
Ca81 ns81 0 1e-12
Ca82 ns82 0 1e-12
Ra81 ns81 0 3536.160082 noise=0
Ra82 ns82 0 3536.160082 noise=0
Ga81 ns81 0 ns82 0 -0.000237869767882
Ga82 ns82 0 ns81 0 0.000237869767882
Ca83 ns83 0 1e-12
Ra83 ns83 0 0.0599459941272 noise=0
Ca84 ns84 0 1e-12
Ra84 ns84 0 0.714606679535 noise=0
Ca85 ns85 0 1e-12
Ra85 ns85 0 1.19287160881 noise=0
Ca86 ns86 0 1e-12
Ca87 ns87 0 1e-12
Ra86 ns86 0 26.828727021 noise=0
Ra87 ns87 0 26.828727021 noise=0
Ga86 ns86 0 ns87 0 -0.518048785893
Ga87 ns87 0 ns86 0 0.518048785893
Ca88 ns88 0 1e-12
Ca89 ns89 0 1e-12
Ra88 ns88 0 90.0406412861 noise=0
Ra89 ns89 0 90.0406412861 noise=0
Ga88 ns88 0 ns89 0 -0.487119257249
Ga89 ns89 0 ns88 0 0.487119257249
Ca90 ns90 0 1e-12
Ca91 ns91 0 1e-12
Ra90 ns90 0 29.4872472308 noise=0
Ra91 ns91 0 29.4872472308 noise=0
Ga90 ns90 0 ns91 0 -0.46382169076
Ga91 ns91 0 ns90 0 0.46382169076
Ca92 ns92 0 1e-12
Ca93 ns93 0 1e-12
Ra92 ns92 0 31.4880587202 noise=0
Ra93 ns93 0 31.4880587202 noise=0
Ga92 ns92 0 ns93 0 -0.426117672518
Ga93 ns93 0 ns92 0 0.426117672518
Ca94 ns94 0 1e-12
Ca95 ns95 0 1e-12
Ra94 ns94 0 19.1952084606 noise=0
Ra95 ns95 0 19.1952084606 noise=0
Ga94 ns94 0 ns95 0 -0.398679757461
Ga95 ns95 0 ns94 0 0.398679757461
Ca96 ns96 0 1e-12
Ca97 ns97 0 1e-12
Ra96 ns96 0 38.9735617239 noise=0
Ra97 ns97 0 38.9735617239 noise=0
Ga96 ns96 0 ns97 0 -0.385574664967
Ga97 ns97 0 ns96 0 0.385574664967
Ca98 ns98 0 1e-12
Ca99 ns99 0 1e-12
Ra98 ns98 0 23.3700179636 noise=0
Ra99 ns99 0 23.3700179636 noise=0
Ga98 ns98 0 ns99 0 -0.32363874977
Ga99 ns99 0 ns98 0 0.32363874977
Ca100 ns100 0 1e-12
Ca101 ns101 0 1e-12
Ra100 ns100 0 13.6366308475 noise=0
Ra101 ns101 0 13.6366308475 noise=0
Ga100 ns100 0 ns101 0 -0.2818027486
Ga101 ns101 0 ns100 0 0.2818027486
Ca102 ns102 0 1e-12
Ca103 ns103 0 1e-12
Ra102 ns102 0 36.4720266288 noise=0
Ra103 ns103 0 36.4720266288 noise=0
Ga102 ns102 0 ns103 0 -0.291418716466
Ga103 ns103 0 ns102 0 0.291418716466
Ca104 ns104 0 1e-12
Ca105 ns105 0 1e-12
Ra104 ns104 0 22.570362028 noise=0
Ra105 ns105 0 22.570362028 noise=0
Ga104 ns104 0 ns105 0 -0.219789949348
Ga105 ns105 0 ns104 0 0.219789949348
Ca106 ns106 0 1e-12
Ca107 ns107 0 1e-12
Ra106 ns106 0 35.3564229023 noise=0
Ra107 ns107 0 35.3564229023 noise=0
Ga106 ns106 0 ns107 0 -0.196387080388
Ga107 ns107 0 ns106 0 0.196387080388
Ca108 ns108 0 1e-12
Ca109 ns109 0 1e-12
Ra108 ns108 0 19.3225792178 noise=0
Ra109 ns109 0 19.3225792178 noise=0
Ga108 ns108 0 ns109 0 -0.158984338989
Ga109 ns109 0 ns108 0 0.158984338989
Ca110 ns110 0 1e-12
Ca111 ns111 0 1e-12
Ra110 ns110 0 22.3171225035 noise=0
Ra111 ns111 0 22.3171225035 noise=0
Ga110 ns110 0 ns111 0 -0.112121022154
Ga111 ns111 0 ns110 0 0.112121022154
Ca112 ns112 0 1e-12
Ca113 ns113 0 1e-12
Ra112 ns112 0 35.6994407039 noise=0
Ra113 ns113 0 35.6994407039 noise=0
Ga112 ns112 0 ns113 0 -0.097312790312
Ga113 ns113 0 ns112 0 0.097312790312
Ca114 ns114 0 1e-12
Ca115 ns115 0 1e-12
Ra114 ns114 0 21.0761624353 noise=0
Ra115 ns115 0 21.0761624353 noise=0
Ga114 ns114 0 ns115 0 -0.0785079694625
Ga115 ns115 0 ns114 0 0.0785079694625
Ca116 ns116 0 1e-12
Ca117 ns117 0 1e-12
Ra116 ns116 0 6461.79173097 noise=0
Ra117 ns117 0 6461.79173097 noise=0
Ga116 ns116 0 ns117 0 -0.0625345296116
Ga117 ns117 0 ns116 0 0.0625345296116
Ca118 ns118 0 1e-12
Ca119 ns119 0 1e-12
Ra118 ns118 0 26.8817745081 noise=0
Ra119 ns119 0 26.8817745081 noise=0
Ga118 ns118 0 ns119 0 -0.016065358588
Ga119 ns119 0 ns118 0 0.016065358588
Ca120 ns120 0 1e-12
Ra120 ns120 0 30.8646103733 noise=0
Ca121 ns121 0 1e-12
Ra121 ns121 0 24137.9690629 noise=0
Ca122 ns122 0 1e-12
Ca123 ns123 0 1e-12
Ra122 ns122 0 3536.160082 noise=0
Ra123 ns123 0 3536.160082 noise=0
Ga122 ns122 0 ns123 0 -0.000237869767882
Ga123 ns123 0 ns122 0 0.000237869767882
Ca124 ns124 0 1e-12
Ra124 ns124 0 0.0599459941272 noise=0
Ca125 ns125 0 1e-12
Ra125 ns125 0 0.714606679535 noise=0
Ca126 ns126 0 1e-12
Ra126 ns126 0 1.19287160881 noise=0
Ca127 ns127 0 1e-12
Ca128 ns128 0 1e-12
Ra127 ns127 0 26.828727021 noise=0
Ra128 ns128 0 26.828727021 noise=0
Ga127 ns127 0 ns128 0 -0.518048785893
Ga128 ns128 0 ns127 0 0.518048785893
Ca129 ns129 0 1e-12
Ca130 ns130 0 1e-12
Ra129 ns129 0 90.0406412861 noise=0
Ra130 ns130 0 90.0406412861 noise=0
Ga129 ns129 0 ns130 0 -0.487119257249
Ga130 ns130 0 ns129 0 0.487119257249
Ca131 ns131 0 1e-12
Ca132 ns132 0 1e-12
Ra131 ns131 0 29.4872472308 noise=0
Ra132 ns132 0 29.4872472308 noise=0
Ga131 ns131 0 ns132 0 -0.46382169076
Ga132 ns132 0 ns131 0 0.46382169076
Ca133 ns133 0 1e-12
Ca134 ns134 0 1e-12
Ra133 ns133 0 31.4880587202 noise=0
Ra134 ns134 0 31.4880587202 noise=0
Ga133 ns133 0 ns134 0 -0.426117672518
Ga134 ns134 0 ns133 0 0.426117672518
Ca135 ns135 0 1e-12
Ca136 ns136 0 1e-12
Ra135 ns135 0 19.1952084606 noise=0
Ra136 ns136 0 19.1952084606 noise=0
Ga135 ns135 0 ns136 0 -0.398679757461
Ga136 ns136 0 ns135 0 0.398679757461
Ca137 ns137 0 1e-12
Ca138 ns138 0 1e-12
Ra137 ns137 0 38.9735617239 noise=0
Ra138 ns138 0 38.9735617239 noise=0
Ga137 ns137 0 ns138 0 -0.385574664967
Ga138 ns138 0 ns137 0 0.385574664967
Ca139 ns139 0 1e-12
Ca140 ns140 0 1e-12
Ra139 ns139 0 23.3700179636 noise=0
Ra140 ns140 0 23.3700179636 noise=0
Ga139 ns139 0 ns140 0 -0.32363874977
Ga140 ns140 0 ns139 0 0.32363874977
Ca141 ns141 0 1e-12
Ca142 ns142 0 1e-12
Ra141 ns141 0 13.6366308475 noise=0
Ra142 ns142 0 13.6366308475 noise=0
Ga141 ns141 0 ns142 0 -0.2818027486
Ga142 ns142 0 ns141 0 0.2818027486
Ca143 ns143 0 1e-12
Ca144 ns144 0 1e-12
Ra143 ns143 0 36.4720266288 noise=0
Ra144 ns144 0 36.4720266288 noise=0
Ga143 ns143 0 ns144 0 -0.291418716466
Ga144 ns144 0 ns143 0 0.291418716466
Ca145 ns145 0 1e-12
Ca146 ns146 0 1e-12
Ra145 ns145 0 22.570362028 noise=0
Ra146 ns146 0 22.570362028 noise=0
Ga145 ns145 0 ns146 0 -0.219789949348
Ga146 ns146 0 ns145 0 0.219789949348
Ca147 ns147 0 1e-12
Ca148 ns148 0 1e-12
Ra147 ns147 0 35.3564229023 noise=0
Ra148 ns148 0 35.3564229023 noise=0
Ga147 ns147 0 ns148 0 -0.196387080388
Ga148 ns148 0 ns147 0 0.196387080388
Ca149 ns149 0 1e-12
Ca150 ns150 0 1e-12
Ra149 ns149 0 19.3225792178 noise=0
Ra150 ns150 0 19.3225792178 noise=0
Ga149 ns149 0 ns150 0 -0.158984338989
Ga150 ns150 0 ns149 0 0.158984338989
Ca151 ns151 0 1e-12
Ca152 ns152 0 1e-12
Ra151 ns151 0 22.3171225035 noise=0
Ra152 ns152 0 22.3171225035 noise=0
Ga151 ns151 0 ns152 0 -0.112121022154
Ga152 ns152 0 ns151 0 0.112121022154
Ca153 ns153 0 1e-12
Ca154 ns154 0 1e-12
Ra153 ns153 0 35.6994407039 noise=0
Ra154 ns154 0 35.6994407039 noise=0
Ga153 ns153 0 ns154 0 -0.097312790312
Ga154 ns154 0 ns153 0 0.097312790312
Ca155 ns155 0 1e-12
Ca156 ns156 0 1e-12
Ra155 ns155 0 21.0761624353 noise=0
Ra156 ns156 0 21.0761624353 noise=0
Ga155 ns155 0 ns156 0 -0.0785079694625
Ga156 ns156 0 ns155 0 0.0785079694625
Ca157 ns157 0 1e-12
Ca158 ns158 0 1e-12
Ra157 ns157 0 6461.79173097 noise=0
Ra158 ns158 0 6461.79173097 noise=0
Ga157 ns157 0 ns158 0 -0.0625345296116
Ga158 ns158 0 ns157 0 0.0625345296116
Ca159 ns159 0 1e-12
Ca160 ns160 0 1e-12
Ra159 ns159 0 26.8817745081 noise=0
Ra160 ns160 0 26.8817745081 noise=0
Ga159 ns159 0 ns160 0 -0.016065358588
Ga160 ns160 0 ns159 0 0.016065358588
Ca161 ns161 0 1e-12
Ra161 ns161 0 30.8646103733 noise=0
Ca162 ns162 0 1e-12
Ra162 ns162 0 24137.9690629 noise=0
Ca163 ns163 0 1e-12
Ca164 ns164 0 1e-12
Ra163 ns163 0 3536.160082 noise=0
Ra164 ns164 0 3536.160082 noise=0
Ga163 ns163 0 ns164 0 -0.000237869767882
Ga164 ns164 0 ns163 0 0.000237869767882
Ca165 ns165 0 1e-12
Ra165 ns165 0 0.0599459941272 noise=0
Ca166 ns166 0 1e-12
Ra166 ns166 0 0.714606679535 noise=0
Ca167 ns167 0 1e-12
Ra167 ns167 0 1.19287160881 noise=0
Ca168 ns168 0 1e-12
Ca169 ns169 0 1e-12
Ra168 ns168 0 26.828727021 noise=0
Ra169 ns169 0 26.828727021 noise=0
Ga168 ns168 0 ns169 0 -0.518048785893
Ga169 ns169 0 ns168 0 0.518048785893
Ca170 ns170 0 1e-12
Ca171 ns171 0 1e-12
Ra170 ns170 0 90.0406412861 noise=0
Ra171 ns171 0 90.0406412861 noise=0
Ga170 ns170 0 ns171 0 -0.487119257249
Ga171 ns171 0 ns170 0 0.487119257249
Ca172 ns172 0 1e-12
Ca173 ns173 0 1e-12
Ra172 ns172 0 29.4872472308 noise=0
Ra173 ns173 0 29.4872472308 noise=0
Ga172 ns172 0 ns173 0 -0.46382169076
Ga173 ns173 0 ns172 0 0.46382169076
Ca174 ns174 0 1e-12
Ca175 ns175 0 1e-12
Ra174 ns174 0 31.4880587202 noise=0
Ra175 ns175 0 31.4880587202 noise=0
Ga174 ns174 0 ns175 0 -0.426117672518
Ga175 ns175 0 ns174 0 0.426117672518
Ca176 ns176 0 1e-12
Ca177 ns177 0 1e-12
Ra176 ns176 0 19.1952084606 noise=0
Ra177 ns177 0 19.1952084606 noise=0
Ga176 ns176 0 ns177 0 -0.398679757461
Ga177 ns177 0 ns176 0 0.398679757461
Ca178 ns178 0 1e-12
Ca179 ns179 0 1e-12
Ra178 ns178 0 38.9735617239 noise=0
Ra179 ns179 0 38.9735617239 noise=0
Ga178 ns178 0 ns179 0 -0.385574664967
Ga179 ns179 0 ns178 0 0.385574664967
Ca180 ns180 0 1e-12
Ca181 ns181 0 1e-12
Ra180 ns180 0 23.3700179636 noise=0
Ra181 ns181 0 23.3700179636 noise=0
Ga180 ns180 0 ns181 0 -0.32363874977
Ga181 ns181 0 ns180 0 0.32363874977
Ca182 ns182 0 1e-12
Ca183 ns183 0 1e-12
Ra182 ns182 0 13.6366308475 noise=0
Ra183 ns183 0 13.6366308475 noise=0
Ga182 ns182 0 ns183 0 -0.2818027486
Ga183 ns183 0 ns182 0 0.2818027486
Ca184 ns184 0 1e-12
Ca185 ns185 0 1e-12
Ra184 ns184 0 36.4720266288 noise=0
Ra185 ns185 0 36.4720266288 noise=0
Ga184 ns184 0 ns185 0 -0.291418716466
Ga185 ns185 0 ns184 0 0.291418716466
Ca186 ns186 0 1e-12
Ca187 ns187 0 1e-12
Ra186 ns186 0 22.570362028 noise=0
Ra187 ns187 0 22.570362028 noise=0
Ga186 ns186 0 ns187 0 -0.219789949348
Ga187 ns187 0 ns186 0 0.219789949348
Ca188 ns188 0 1e-12
Ca189 ns189 0 1e-12
Ra188 ns188 0 35.3564229023 noise=0
Ra189 ns189 0 35.3564229023 noise=0
Ga188 ns188 0 ns189 0 -0.196387080388
Ga189 ns189 0 ns188 0 0.196387080388
Ca190 ns190 0 1e-12
Ca191 ns191 0 1e-12
Ra190 ns190 0 19.3225792178 noise=0
Ra191 ns191 0 19.3225792178 noise=0
Ga190 ns190 0 ns191 0 -0.158984338989
Ga191 ns191 0 ns190 0 0.158984338989
Ca192 ns192 0 1e-12
Ca193 ns193 0 1e-12
Ra192 ns192 0 22.3171225035 noise=0
Ra193 ns193 0 22.3171225035 noise=0
Ga192 ns192 0 ns193 0 -0.112121022154
Ga193 ns193 0 ns192 0 0.112121022154
Ca194 ns194 0 1e-12
Ca195 ns195 0 1e-12
Ra194 ns194 0 35.6994407039 noise=0
Ra195 ns195 0 35.6994407039 noise=0
Ga194 ns194 0 ns195 0 -0.097312790312
Ga195 ns195 0 ns194 0 0.097312790312
Ca196 ns196 0 1e-12
Ca197 ns197 0 1e-12
Ra196 ns196 0 21.0761624353 noise=0
Ra197 ns197 0 21.0761624353 noise=0
Ga196 ns196 0 ns197 0 -0.0785079694625
Ga197 ns197 0 ns196 0 0.0785079694625
Ca198 ns198 0 1e-12
Ca199 ns199 0 1e-12
Ra198 ns198 0 6461.79173097 noise=0
Ra199 ns199 0 6461.79173097 noise=0
Ga198 ns198 0 ns199 0 -0.0625345296116
Ga199 ns199 0 ns198 0 0.0625345296116
Ca200 ns200 0 1e-12
Ca201 ns201 0 1e-12
Ra200 ns200 0 26.8817745081 noise=0
Ra201 ns201 0 26.8817745081 noise=0
Ga200 ns200 0 ns201 0 -0.016065358588
Ga201 ns201 0 ns200 0 0.016065358588
Ca202 ns202 0 1e-12
Ra202 ns202 0 30.8646103733 noise=0
Ca203 ns203 0 1e-12
Ra203 ns203 0 24137.9690629 noise=0
Ca204 ns204 0 1e-12
Ca205 ns205 0 1e-12
Ra204 ns204 0 3536.160082 noise=0
Ra205 ns205 0 3536.160082 noise=0
Ga204 ns204 0 ns205 0 -0.000237869767882
Ga205 ns205 0 ns204 0 0.000237869767882
Ca206 ns206 0 1e-12
Ra206 ns206 0 0.0599459941272 noise=0
Ca207 ns207 0 1e-12
Ra207 ns207 0 0.714606679535 noise=0
Ca208 ns208 0 1e-12
Ra208 ns208 0 1.19287160881 noise=0
Ca209 ns209 0 1e-12
Ca210 ns210 0 1e-12
Ra209 ns209 0 26.828727021 noise=0
Ra210 ns210 0 26.828727021 noise=0
Ga209 ns209 0 ns210 0 -0.518048785893
Ga210 ns210 0 ns209 0 0.518048785893
Ca211 ns211 0 1e-12
Ca212 ns212 0 1e-12
Ra211 ns211 0 90.0406412861 noise=0
Ra212 ns212 0 90.0406412861 noise=0
Ga211 ns211 0 ns212 0 -0.487119257249
Ga212 ns212 0 ns211 0 0.487119257249
Ca213 ns213 0 1e-12
Ca214 ns214 0 1e-12
Ra213 ns213 0 29.4872472308 noise=0
Ra214 ns214 0 29.4872472308 noise=0
Ga213 ns213 0 ns214 0 -0.46382169076
Ga214 ns214 0 ns213 0 0.46382169076
Ca215 ns215 0 1e-12
Ca216 ns216 0 1e-12
Ra215 ns215 0 31.4880587202 noise=0
Ra216 ns216 0 31.4880587202 noise=0
Ga215 ns215 0 ns216 0 -0.426117672518
Ga216 ns216 0 ns215 0 0.426117672518
Ca217 ns217 0 1e-12
Ca218 ns218 0 1e-12
Ra217 ns217 0 19.1952084606 noise=0
Ra218 ns218 0 19.1952084606 noise=0
Ga217 ns217 0 ns218 0 -0.398679757461
Ga218 ns218 0 ns217 0 0.398679757461
Ca219 ns219 0 1e-12
Ca220 ns220 0 1e-12
Ra219 ns219 0 38.9735617239 noise=0
Ra220 ns220 0 38.9735617239 noise=0
Ga219 ns219 0 ns220 0 -0.385574664967
Ga220 ns220 0 ns219 0 0.385574664967
Ca221 ns221 0 1e-12
Ca222 ns222 0 1e-12
Ra221 ns221 0 23.3700179636 noise=0
Ra222 ns222 0 23.3700179636 noise=0
Ga221 ns221 0 ns222 0 -0.32363874977
Ga222 ns222 0 ns221 0 0.32363874977
Ca223 ns223 0 1e-12
Ca224 ns224 0 1e-12
Ra223 ns223 0 13.6366308475 noise=0
Ra224 ns224 0 13.6366308475 noise=0
Ga223 ns223 0 ns224 0 -0.2818027486
Ga224 ns224 0 ns223 0 0.2818027486
Ca225 ns225 0 1e-12
Ca226 ns226 0 1e-12
Ra225 ns225 0 36.4720266288 noise=0
Ra226 ns226 0 36.4720266288 noise=0
Ga225 ns225 0 ns226 0 -0.291418716466
Ga226 ns226 0 ns225 0 0.291418716466
Ca227 ns227 0 1e-12
Ca228 ns228 0 1e-12
Ra227 ns227 0 22.570362028 noise=0
Ra228 ns228 0 22.570362028 noise=0
Ga227 ns227 0 ns228 0 -0.219789949348
Ga228 ns228 0 ns227 0 0.219789949348
Ca229 ns229 0 1e-12
Ca230 ns230 0 1e-12
Ra229 ns229 0 35.3564229023 noise=0
Ra230 ns230 0 35.3564229023 noise=0
Ga229 ns229 0 ns230 0 -0.196387080388
Ga230 ns230 0 ns229 0 0.196387080388
Ca231 ns231 0 1e-12
Ca232 ns232 0 1e-12
Ra231 ns231 0 19.3225792178 noise=0
Ra232 ns232 0 19.3225792178 noise=0
Ga231 ns231 0 ns232 0 -0.158984338989
Ga232 ns232 0 ns231 0 0.158984338989
Ca233 ns233 0 1e-12
Ca234 ns234 0 1e-12
Ra233 ns233 0 22.3171225035 noise=0
Ra234 ns234 0 22.3171225035 noise=0
Ga233 ns233 0 ns234 0 -0.112121022154
Ga234 ns234 0 ns233 0 0.112121022154
Ca235 ns235 0 1e-12
Ca236 ns236 0 1e-12
Ra235 ns235 0 35.6994407039 noise=0
Ra236 ns236 0 35.6994407039 noise=0
Ga235 ns235 0 ns236 0 -0.097312790312
Ga236 ns236 0 ns235 0 0.097312790312
Ca237 ns237 0 1e-12
Ca238 ns238 0 1e-12
Ra237 ns237 0 21.0761624353 noise=0
Ra238 ns238 0 21.0761624353 noise=0
Ga237 ns237 0 ns238 0 -0.0785079694625
Ga238 ns238 0 ns237 0 0.0785079694625
Ca239 ns239 0 1e-12
Ca240 ns240 0 1e-12
Ra239 ns239 0 6461.79173097 noise=0
Ra240 ns240 0 6461.79173097 noise=0
Ga239 ns239 0 ns240 0 -0.0625345296116
Ga240 ns240 0 ns239 0 0.0625345296116
Ca241 ns241 0 1e-12
Ca242 ns242 0 1e-12
Ra241 ns241 0 26.8817745081 noise=0
Ra242 ns242 0 26.8817745081 noise=0
Ga241 ns241 0 ns242 0 -0.016065358588
Ga242 ns242 0 ns241 0 0.016065358588
Ca243 ns243 0 1e-12
Ra243 ns243 0 30.8646103733 noise=0
Ca244 ns244 0 1e-12
Ra244 ns244 0 24137.9690629 noise=0
Ca245 ns245 0 1e-12
Ca246 ns246 0 1e-12
Ra245 ns245 0 3536.160082 noise=0
Ra246 ns246 0 3536.160082 noise=0
Ga245 ns245 0 ns246 0 -0.000237869767882
Ga246 ns246 0 ns245 0 0.000237869767882
Ca247 ns247 0 1e-12
Ra247 ns247 0 0.0599459941272 noise=0
Ca248 ns248 0 1e-12
Ra248 ns248 0 0.714606679535 noise=0
Ca249 ns249 0 1e-12
Ra249 ns249 0 1.19287160881 noise=0
Ca250 ns250 0 1e-12
Ca251 ns251 0 1e-12
Ra250 ns250 0 26.828727021 noise=0
Ra251 ns251 0 26.828727021 noise=0
Ga250 ns250 0 ns251 0 -0.518048785893
Ga251 ns251 0 ns250 0 0.518048785893
Ca252 ns252 0 1e-12
Ca253 ns253 0 1e-12
Ra252 ns252 0 90.0406412861 noise=0
Ra253 ns253 0 90.0406412861 noise=0
Ga252 ns252 0 ns253 0 -0.487119257249
Ga253 ns253 0 ns252 0 0.487119257249
Ca254 ns254 0 1e-12
Ca255 ns255 0 1e-12
Ra254 ns254 0 29.4872472308 noise=0
Ra255 ns255 0 29.4872472308 noise=0
Ga254 ns254 0 ns255 0 -0.46382169076
Ga255 ns255 0 ns254 0 0.46382169076
Ca256 ns256 0 1e-12
Ca257 ns257 0 1e-12
Ra256 ns256 0 31.4880587202 noise=0
Ra257 ns257 0 31.4880587202 noise=0
Ga256 ns256 0 ns257 0 -0.426117672518
Ga257 ns257 0 ns256 0 0.426117672518
Ca258 ns258 0 1e-12
Ca259 ns259 0 1e-12
Ra258 ns258 0 19.1952084606 noise=0
Ra259 ns259 0 19.1952084606 noise=0
Ga258 ns258 0 ns259 0 -0.398679757461
Ga259 ns259 0 ns258 0 0.398679757461
Ca260 ns260 0 1e-12
Ca261 ns261 0 1e-12
Ra260 ns260 0 38.9735617239 noise=0
Ra261 ns261 0 38.9735617239 noise=0
Ga260 ns260 0 ns261 0 -0.385574664967
Ga261 ns261 0 ns260 0 0.385574664967
Ca262 ns262 0 1e-12
Ca263 ns263 0 1e-12
Ra262 ns262 0 23.3700179636 noise=0
Ra263 ns263 0 23.3700179636 noise=0
Ga262 ns262 0 ns263 0 -0.32363874977
Ga263 ns263 0 ns262 0 0.32363874977
Ca264 ns264 0 1e-12
Ca265 ns265 0 1e-12
Ra264 ns264 0 13.6366308475 noise=0
Ra265 ns265 0 13.6366308475 noise=0
Ga264 ns264 0 ns265 0 -0.2818027486
Ga265 ns265 0 ns264 0 0.2818027486
Ca266 ns266 0 1e-12
Ca267 ns267 0 1e-12
Ra266 ns266 0 36.4720266288 noise=0
Ra267 ns267 0 36.4720266288 noise=0
Ga266 ns266 0 ns267 0 -0.291418716466
Ga267 ns267 0 ns266 0 0.291418716466
Ca268 ns268 0 1e-12
Ca269 ns269 0 1e-12
Ra268 ns268 0 22.570362028 noise=0
Ra269 ns269 0 22.570362028 noise=0
Ga268 ns268 0 ns269 0 -0.219789949348
Ga269 ns269 0 ns268 0 0.219789949348
Ca270 ns270 0 1e-12
Ca271 ns271 0 1e-12
Ra270 ns270 0 35.3564229023 noise=0
Ra271 ns271 0 35.3564229023 noise=0
Ga270 ns270 0 ns271 0 -0.196387080388
Ga271 ns271 0 ns270 0 0.196387080388
Ca272 ns272 0 1e-12
Ca273 ns273 0 1e-12
Ra272 ns272 0 19.3225792178 noise=0
Ra273 ns273 0 19.3225792178 noise=0
Ga272 ns272 0 ns273 0 -0.158984338989
Ga273 ns273 0 ns272 0 0.158984338989
Ca274 ns274 0 1e-12
Ca275 ns275 0 1e-12
Ra274 ns274 0 22.3171225035 noise=0
Ra275 ns275 0 22.3171225035 noise=0
Ga274 ns274 0 ns275 0 -0.112121022154
Ga275 ns275 0 ns274 0 0.112121022154
Ca276 ns276 0 1e-12
Ca277 ns277 0 1e-12
Ra276 ns276 0 35.6994407039 noise=0
Ra277 ns277 0 35.6994407039 noise=0
Ga276 ns276 0 ns277 0 -0.097312790312
Ga277 ns277 0 ns276 0 0.097312790312
Ca278 ns278 0 1e-12
Ca279 ns279 0 1e-12
Ra278 ns278 0 21.0761624353 noise=0
Ra279 ns279 0 21.0761624353 noise=0
Ga278 ns278 0 ns279 0 -0.0785079694625
Ga279 ns279 0 ns278 0 0.0785079694625
Ca280 ns280 0 1e-12
Ca281 ns281 0 1e-12
Ra280 ns280 0 6461.79173097 noise=0
Ra281 ns281 0 6461.79173097 noise=0
Ga280 ns280 0 ns281 0 -0.0625345296116
Ga281 ns281 0 ns280 0 0.0625345296116
Ca282 ns282 0 1e-12
Ca283 ns283 0 1e-12
Ra282 ns282 0 26.8817745081 noise=0
Ra283 ns283 0 26.8817745081 noise=0
Ga282 ns282 0 ns283 0 -0.016065358588
Ga283 ns283 0 ns282 0 0.016065358588
Ca284 ns284 0 1e-12
Ra284 ns284 0 30.8646103733 noise=0
Ca285 ns285 0 1e-12
Ra285 ns285 0 24137.9690629 noise=0
Ca286 ns286 0 1e-12
Ca287 ns287 0 1e-12
Ra286 ns286 0 3536.160082 noise=0
Ra287 ns287 0 3536.160082 noise=0
Ga286 ns286 0 ns287 0 -0.000237869767882
Ga287 ns287 0 ns286 0 0.000237869767882
Ca288 ns288 0 1e-12
Ra288 ns288 0 0.0599459941272 noise=0
Ca289 ns289 0 1e-12
Ra289 ns289 0 0.714606679535 noise=0
Ca290 ns290 0 1e-12
Ra290 ns290 0 1.19287160881 noise=0
Ca291 ns291 0 1e-12
Ca292 ns292 0 1e-12
Ra291 ns291 0 26.828727021 noise=0
Ra292 ns292 0 26.828727021 noise=0
Ga291 ns291 0 ns292 0 -0.518048785893
Ga292 ns292 0 ns291 0 0.518048785893
Ca293 ns293 0 1e-12
Ca294 ns294 0 1e-12
Ra293 ns293 0 90.0406412861 noise=0
Ra294 ns294 0 90.0406412861 noise=0
Ga293 ns293 0 ns294 0 -0.487119257249
Ga294 ns294 0 ns293 0 0.487119257249
Ca295 ns295 0 1e-12
Ca296 ns296 0 1e-12
Ra295 ns295 0 29.4872472308 noise=0
Ra296 ns296 0 29.4872472308 noise=0
Ga295 ns295 0 ns296 0 -0.46382169076
Ga296 ns296 0 ns295 0 0.46382169076
Ca297 ns297 0 1e-12
Ca298 ns298 0 1e-12
Ra297 ns297 0 31.4880587202 noise=0
Ra298 ns298 0 31.4880587202 noise=0
Ga297 ns297 0 ns298 0 -0.426117672518
Ga298 ns298 0 ns297 0 0.426117672518
Ca299 ns299 0 1e-12
Ca300 ns300 0 1e-12
Ra299 ns299 0 19.1952084606 noise=0
Ra300 ns300 0 19.1952084606 noise=0
Ga299 ns299 0 ns300 0 -0.398679757461
Ga300 ns300 0 ns299 0 0.398679757461
Ca301 ns301 0 1e-12
Ca302 ns302 0 1e-12
Ra301 ns301 0 38.9735617239 noise=0
Ra302 ns302 0 38.9735617239 noise=0
Ga301 ns301 0 ns302 0 -0.385574664967
Ga302 ns302 0 ns301 0 0.385574664967
Ca303 ns303 0 1e-12
Ca304 ns304 0 1e-12
Ra303 ns303 0 23.3700179636 noise=0
Ra304 ns304 0 23.3700179636 noise=0
Ga303 ns303 0 ns304 0 -0.32363874977
Ga304 ns304 0 ns303 0 0.32363874977
Ca305 ns305 0 1e-12
Ca306 ns306 0 1e-12
Ra305 ns305 0 13.6366308475 noise=0
Ra306 ns306 0 13.6366308475 noise=0
Ga305 ns305 0 ns306 0 -0.2818027486
Ga306 ns306 0 ns305 0 0.2818027486
Ca307 ns307 0 1e-12
Ca308 ns308 0 1e-12
Ra307 ns307 0 36.4720266288 noise=0
Ra308 ns308 0 36.4720266288 noise=0
Ga307 ns307 0 ns308 0 -0.291418716466
Ga308 ns308 0 ns307 0 0.291418716466
Ca309 ns309 0 1e-12
Ca310 ns310 0 1e-12
Ra309 ns309 0 22.570362028 noise=0
Ra310 ns310 0 22.570362028 noise=0
Ga309 ns309 0 ns310 0 -0.219789949348
Ga310 ns310 0 ns309 0 0.219789949348
Ca311 ns311 0 1e-12
Ca312 ns312 0 1e-12
Ra311 ns311 0 35.3564229023 noise=0
Ra312 ns312 0 35.3564229023 noise=0
Ga311 ns311 0 ns312 0 -0.196387080388
Ga312 ns312 0 ns311 0 0.196387080388
Ca313 ns313 0 1e-12
Ca314 ns314 0 1e-12
Ra313 ns313 0 19.3225792178 noise=0
Ra314 ns314 0 19.3225792178 noise=0
Ga313 ns313 0 ns314 0 -0.158984338989
Ga314 ns314 0 ns313 0 0.158984338989
Ca315 ns315 0 1e-12
Ca316 ns316 0 1e-12
Ra315 ns315 0 22.3171225035 noise=0
Ra316 ns316 0 22.3171225035 noise=0
Ga315 ns315 0 ns316 0 -0.112121022154
Ga316 ns316 0 ns315 0 0.112121022154
Ca317 ns317 0 1e-12
Ca318 ns318 0 1e-12
Ra317 ns317 0 35.6994407039 noise=0
Ra318 ns318 0 35.6994407039 noise=0
Ga317 ns317 0 ns318 0 -0.097312790312
Ga318 ns318 0 ns317 0 0.097312790312
Ca319 ns319 0 1e-12
Ca320 ns320 0 1e-12
Ra319 ns319 0 21.0761624353 noise=0
Ra320 ns320 0 21.0761624353 noise=0
Ga319 ns319 0 ns320 0 -0.0785079694625
Ga320 ns320 0 ns319 0 0.0785079694625
Ca321 ns321 0 1e-12
Ca322 ns322 0 1e-12
Ra321 ns321 0 6461.79173097 noise=0
Ra322 ns322 0 6461.79173097 noise=0
Ga321 ns321 0 ns322 0 -0.0625345296116
Ga322 ns322 0 ns321 0 0.0625345296116
Ca323 ns323 0 1e-12
Ca324 ns324 0 1e-12
Ra323 ns323 0 26.8817745081 noise=0
Ra324 ns324 0 26.8817745081 noise=0
Ga323 ns323 0 ns324 0 -0.016065358588
Ga324 ns324 0 ns323 0 0.016065358588
Ca325 ns325 0 1e-12
Ra325 ns325 0 30.8646103733 noise=0
Ca326 ns326 0 1e-12
Ra326 ns326 0 24137.9690629 noise=0
Ca327 ns327 0 1e-12
Ca328 ns328 0 1e-12
Ra327 ns327 0 3536.160082 noise=0
Ra328 ns328 0 3536.160082 noise=0
Ga327 ns327 0 ns328 0 -0.000237869767882
Ga328 ns328 0 ns327 0 0.000237869767882

Gb1_1 ns1 0 ni1 0 16.6816818131
Gb2_1 ns2 0 ni1 0 1.39937119067
Gb3_1 ns3 0 ni1 0 -0.838313186945
Gb4_1 ns4 0 ni1 0 0.178221203364
Gb5_1 ns5 0 ni1 0 -0.507907632755
Gb6_1 ns6 0 ni1 0 -0.0008419118152
Gb7_1 ns7 0 ni1 0 0.487353275945
Gb8_1 ns8 0 ni1 0 -0.453187972971
Gb9_1 ns9 0 ni1 0 -0.179348461456
Gb10_1 ns10 0 ni1 0 -0.267410962593
Gb11_1 ns11 0 ni1 0 -0.408554727547
Gb12_1 ns12 0 ni1 0 -0.398757728834
Gb13_1 ns13 0 ni1 0 -0.0514996397364
Gb14_1 ns14 0 ni1 0 -0.38110118275
Gb15_1 ns15 0 ni1 0 0.0928824121159
Gb16_1 ns16 0 ni1 0 -0.328038226621
Gb17_1 ns17 0 ni1 0 0.00951467455824
Gb18_1 ns18 0 ni1 0 -0.273688132867
Gb19_1 ns19 0 ni1 0 0.104515066725
Gb20_1 ns20 0 ni1 0 0.021639783359
Gb21_1 ns21 0 ni1 0 0.291962388554
Gb22_1 ns22 0 ni1 0 0.228255995922
Gb23_1 ns23 0 ni1 0 -0.00230804590343
Gb24_1 ns24 0 ni1 0 -0.0353048726126
Gb25_1 ns25 0 ni1 0 -0.195375857914
Gb26_1 ns26 0 ni1 0 0.158298219061
Gb27_1 ns27 0 ni1 0 -0.0538606771897
Gb28_1 ns28 0 ni1 0 -0.125266532438
Gb29_1 ns29 0 ni1 0 0.0119157039555
Gb30_1 ns30 0 ni1 0 0.0397996579039
Gb31_1 ns31 0 ni1 0 0.0939195913421
Gb32_1 ns32 0 ni1 0 0.0237488618908
Gb33_1 ns33 0 ni1 0 -0.092830123943
Gb34_1 ns34 0 ni1 0 0.00194300457983
Gb35_1 ns35 0 ni1 0 -0.0625301041856
Gb36_1 ns36 0 ni1 0 -0.0395543648239
Gb37_1 ns37 0 ni1 0 -0.0106135674783
Gb38_1 ns38 0 ni1 0 0.0323995666203
Gb39_1 ns39 0 ni1 0 4.14285061595e-05
Gb40_1 ns40 0 ni1 0 -3.6782420325e-05
Gb41_1 ns41 0 ni1 0 0.000451936360429
Gb42_2 ns42 0 ni2 0 16.6816818131
Gb43_2 ns43 0 ni2 0 1.39937119067
Gb44_2 ns44 0 ni2 0 -0.838313186945
Gb45_2 ns45 0 ni2 0 0.178221203364
Gb46_2 ns46 0 ni2 0 -0.507907632755
Gb47_2 ns47 0 ni2 0 -0.0008419118152
Gb48_2 ns48 0 ni2 0 0.487353275945
Gb49_2 ns49 0 ni2 0 -0.453187972971
Gb50_2 ns50 0 ni2 0 -0.179348461456
Gb51_2 ns51 0 ni2 0 -0.267410962593
Gb52_2 ns52 0 ni2 0 -0.408554727547
Gb53_2 ns53 0 ni2 0 -0.398757728834
Gb54_2 ns54 0 ni2 0 -0.0514996397364
Gb55_2 ns55 0 ni2 0 -0.38110118275
Gb56_2 ns56 0 ni2 0 0.0928824121159
Gb57_2 ns57 0 ni2 0 -0.328038226621
Gb58_2 ns58 0 ni2 0 0.00951467455824
Gb59_2 ns59 0 ni2 0 -0.273688132867
Gb60_2 ns60 0 ni2 0 0.104515066725
Gb61_2 ns61 0 ni2 0 0.021639783359
Gb62_2 ns62 0 ni2 0 0.291962388554
Gb63_2 ns63 0 ni2 0 0.228255995922
Gb64_2 ns64 0 ni2 0 -0.00230804590343
Gb65_2 ns65 0 ni2 0 -0.0353048726126
Gb66_2 ns66 0 ni2 0 -0.195375857914
Gb67_2 ns67 0 ni2 0 0.158298219061
Gb68_2 ns68 0 ni2 0 -0.0538606771897
Gb69_2 ns69 0 ni2 0 -0.125266532438
Gb70_2 ns70 0 ni2 0 0.0119157039555
Gb71_2 ns71 0 ni2 0 0.0397996579039
Gb72_2 ns72 0 ni2 0 0.0939195913421
Gb73_2 ns73 0 ni2 0 0.0237488618908
Gb74_2 ns74 0 ni2 0 -0.092830123943
Gb75_2 ns75 0 ni2 0 0.00194300457983
Gb76_2 ns76 0 ni2 0 -0.0625301041856
Gb77_2 ns77 0 ni2 0 -0.0395543648239
Gb78_2 ns78 0 ni2 0 -0.0106135674783
Gb79_2 ns79 0 ni2 0 0.0323995666203
Gb80_2 ns80 0 ni2 0 4.14285061595e-05
Gb81_2 ns81 0 ni2 0 -3.6782420325e-05
Gb82_2 ns82 0 ni2 0 0.000451936360429
Gb83_3 ns83 0 ni3 0 16.6816818131
Gb84_3 ns84 0 ni3 0 1.39937119067
Gb85_3 ns85 0 ni3 0 -0.838313186945
Gb86_3 ns86 0 ni3 0 0.178221203364
Gb87_3 ns87 0 ni3 0 -0.507907632755
Gb88_3 ns88 0 ni3 0 -0.0008419118152
Gb89_3 ns89 0 ni3 0 0.487353275945
Gb90_3 ns90 0 ni3 0 -0.453187972971
Gb91_3 ns91 0 ni3 0 -0.179348461456
Gb92_3 ns92 0 ni3 0 -0.267410962593
Gb93_3 ns93 0 ni3 0 -0.408554727547
Gb94_3 ns94 0 ni3 0 -0.398757728834
Gb95_3 ns95 0 ni3 0 -0.0514996397364
Gb96_3 ns96 0 ni3 0 -0.38110118275
Gb97_3 ns97 0 ni3 0 0.0928824121159
Gb98_3 ns98 0 ni3 0 -0.328038226621
Gb99_3 ns99 0 ni3 0 0.00951467455824
Gb100_3 ns100 0 ni3 0 -0.273688132867
Gb101_3 ns101 0 ni3 0 0.104515066725
Gb102_3 ns102 0 ni3 0 0.021639783359
Gb103_3 ns103 0 ni3 0 0.291962388554
Gb104_3 ns104 0 ni3 0 0.228255995922
Gb105_3 ns105 0 ni3 0 -0.00230804590343
Gb106_3 ns106 0 ni3 0 -0.0353048726126
Gb107_3 ns107 0 ni3 0 -0.195375857914
Gb108_3 ns108 0 ni3 0 0.158298219061
Gb109_3 ns109 0 ni3 0 -0.0538606771897
Gb110_3 ns110 0 ni3 0 -0.125266532438
Gb111_3 ns111 0 ni3 0 0.0119157039555
Gb112_3 ns112 0 ni3 0 0.0397996579039
Gb113_3 ns113 0 ni3 0 0.0939195913421
Gb114_3 ns114 0 ni3 0 0.0237488618908
Gb115_3 ns115 0 ni3 0 -0.092830123943
Gb116_3 ns116 0 ni3 0 0.00194300457983
Gb117_3 ns117 0 ni3 0 -0.0625301041856
Gb118_3 ns118 0 ni3 0 -0.0395543648239
Gb119_3 ns119 0 ni3 0 -0.0106135674783
Gb120_3 ns120 0 ni3 0 0.0323995666203
Gb121_3 ns121 0 ni3 0 4.14285061595e-05
Gb122_3 ns122 0 ni3 0 -3.6782420325e-05
Gb123_3 ns123 0 ni3 0 0.000451936360429
Gb124_4 ns124 0 ni4 0 16.6816818131
Gb125_4 ns125 0 ni4 0 1.39937119067
Gb126_4 ns126 0 ni4 0 -0.838313186945
Gb127_4 ns127 0 ni4 0 0.178221203364
Gb128_4 ns128 0 ni4 0 -0.507907632755
Gb129_4 ns129 0 ni4 0 -0.0008419118152
Gb130_4 ns130 0 ni4 0 0.487353275945
Gb131_4 ns131 0 ni4 0 -0.453187972971
Gb132_4 ns132 0 ni4 0 -0.179348461456
Gb133_4 ns133 0 ni4 0 -0.267410962593
Gb134_4 ns134 0 ni4 0 -0.408554727547
Gb135_4 ns135 0 ni4 0 -0.398757728834
Gb136_4 ns136 0 ni4 0 -0.0514996397364
Gb137_4 ns137 0 ni4 0 -0.38110118275
Gb138_4 ns138 0 ni4 0 0.0928824121159
Gb139_4 ns139 0 ni4 0 -0.328038226621
Gb140_4 ns140 0 ni4 0 0.00951467455824
Gb141_4 ns141 0 ni4 0 -0.273688132867
Gb142_4 ns142 0 ni4 0 0.104515066725
Gb143_4 ns143 0 ni4 0 0.021639783359
Gb144_4 ns144 0 ni4 0 0.291962388554
Gb145_4 ns145 0 ni4 0 0.228255995922
Gb146_4 ns146 0 ni4 0 -0.00230804590343
Gb147_4 ns147 0 ni4 0 -0.0353048726126
Gb148_4 ns148 0 ni4 0 -0.195375857914
Gb149_4 ns149 0 ni4 0 0.158298219061
Gb150_4 ns150 0 ni4 0 -0.0538606771897
Gb151_4 ns151 0 ni4 0 -0.125266532438
Gb152_4 ns152 0 ni4 0 0.0119157039555
Gb153_4 ns153 0 ni4 0 0.0397996579039
Gb154_4 ns154 0 ni4 0 0.0939195913421
Gb155_4 ns155 0 ni4 0 0.0237488618908
Gb156_4 ns156 0 ni4 0 -0.092830123943
Gb157_4 ns157 0 ni4 0 0.00194300457983
Gb158_4 ns158 0 ni4 0 -0.0625301041856
Gb159_4 ns159 0 ni4 0 -0.0395543648239
Gb160_4 ns160 0 ni4 0 -0.0106135674783
Gb161_4 ns161 0 ni4 0 0.0323995666203
Gb162_4 ns162 0 ni4 0 4.14285061595e-05
Gb163_4 ns163 0 ni4 0 -3.6782420325e-05
Gb164_4 ns164 0 ni4 0 0.000451936360429
Gb165_5 ns165 0 ni5 0 16.6816818131
Gb166_5 ns166 0 ni5 0 1.39937119067
Gb167_5 ns167 0 ni5 0 -0.838313186945
Gb168_5 ns168 0 ni5 0 0.178221203364
Gb169_5 ns169 0 ni5 0 -0.507907632755
Gb170_5 ns170 0 ni5 0 -0.0008419118152
Gb171_5 ns171 0 ni5 0 0.487353275945
Gb172_5 ns172 0 ni5 0 -0.453187972971
Gb173_5 ns173 0 ni5 0 -0.179348461456
Gb174_5 ns174 0 ni5 0 -0.267410962593
Gb175_5 ns175 0 ni5 0 -0.408554727547
Gb176_5 ns176 0 ni5 0 -0.398757728834
Gb177_5 ns177 0 ni5 0 -0.0514996397364
Gb178_5 ns178 0 ni5 0 -0.38110118275
Gb179_5 ns179 0 ni5 0 0.0928824121159
Gb180_5 ns180 0 ni5 0 -0.328038226621
Gb181_5 ns181 0 ni5 0 0.00951467455824
Gb182_5 ns182 0 ni5 0 -0.273688132867
Gb183_5 ns183 0 ni5 0 0.104515066725
Gb184_5 ns184 0 ni5 0 0.021639783359
Gb185_5 ns185 0 ni5 0 0.291962388554
Gb186_5 ns186 0 ni5 0 0.228255995922
Gb187_5 ns187 0 ni5 0 -0.00230804590343
Gb188_5 ns188 0 ni5 0 -0.0353048726126
Gb189_5 ns189 0 ni5 0 -0.195375857914
Gb190_5 ns190 0 ni5 0 0.158298219061
Gb191_5 ns191 0 ni5 0 -0.0538606771897
Gb192_5 ns192 0 ni5 0 -0.125266532438
Gb193_5 ns193 0 ni5 0 0.0119157039555
Gb194_5 ns194 0 ni5 0 0.0397996579039
Gb195_5 ns195 0 ni5 0 0.0939195913421
Gb196_5 ns196 0 ni5 0 0.0237488618908
Gb197_5 ns197 0 ni5 0 -0.092830123943
Gb198_5 ns198 0 ni5 0 0.00194300457983
Gb199_5 ns199 0 ni5 0 -0.0625301041856
Gb200_5 ns200 0 ni5 0 -0.0395543648239
Gb201_5 ns201 0 ni5 0 -0.0106135674783
Gb202_5 ns202 0 ni5 0 0.0323995666203
Gb203_5 ns203 0 ni5 0 4.14285061595e-05
Gb204_5 ns204 0 ni5 0 -3.6782420325e-05
Gb205_5 ns205 0 ni5 0 0.000451936360429
Gb206_6 ns206 0 ni6 0 16.6816818131
Gb207_6 ns207 0 ni6 0 1.39937119067
Gb208_6 ns208 0 ni6 0 -0.838313186945
Gb209_6 ns209 0 ni6 0 0.178221203364
Gb210_6 ns210 0 ni6 0 -0.507907632755
Gb211_6 ns211 0 ni6 0 -0.0008419118152
Gb212_6 ns212 0 ni6 0 0.487353275945
Gb213_6 ns213 0 ni6 0 -0.453187972971
Gb214_6 ns214 0 ni6 0 -0.179348461456
Gb215_6 ns215 0 ni6 0 -0.267410962593
Gb216_6 ns216 0 ni6 0 -0.408554727547
Gb217_6 ns217 0 ni6 0 -0.398757728834
Gb218_6 ns218 0 ni6 0 -0.0514996397364
Gb219_6 ns219 0 ni6 0 -0.38110118275
Gb220_6 ns220 0 ni6 0 0.0928824121159
Gb221_6 ns221 0 ni6 0 -0.328038226621
Gb222_6 ns222 0 ni6 0 0.00951467455824
Gb223_6 ns223 0 ni6 0 -0.273688132867
Gb224_6 ns224 0 ni6 0 0.104515066725
Gb225_6 ns225 0 ni6 0 0.021639783359
Gb226_6 ns226 0 ni6 0 0.291962388554
Gb227_6 ns227 0 ni6 0 0.228255995922
Gb228_6 ns228 0 ni6 0 -0.00230804590343
Gb229_6 ns229 0 ni6 0 -0.0353048726126
Gb230_6 ns230 0 ni6 0 -0.195375857914
Gb231_6 ns231 0 ni6 0 0.158298219061
Gb232_6 ns232 0 ni6 0 -0.0538606771897
Gb233_6 ns233 0 ni6 0 -0.125266532438
Gb234_6 ns234 0 ni6 0 0.0119157039555
Gb235_6 ns235 0 ni6 0 0.0397996579039
Gb236_6 ns236 0 ni6 0 0.0939195913421
Gb237_6 ns237 0 ni6 0 0.0237488618908
Gb238_6 ns238 0 ni6 0 -0.092830123943
Gb239_6 ns239 0 ni6 0 0.00194300457983
Gb240_6 ns240 0 ni6 0 -0.0625301041856
Gb241_6 ns241 0 ni6 0 -0.0395543648239
Gb242_6 ns242 0 ni6 0 -0.0106135674783
Gb243_6 ns243 0 ni6 0 0.0323995666203
Gb244_6 ns244 0 ni6 0 4.14285061595e-05
Gb245_6 ns245 0 ni6 0 -3.6782420325e-05
Gb246_6 ns246 0 ni6 0 0.000451936360429
Gb247_7 ns247 0 ni7 0 16.6816818131
Gb248_7 ns248 0 ni7 0 1.39937119067
Gb249_7 ns249 0 ni7 0 -0.838313186945
Gb250_7 ns250 0 ni7 0 0.178221203364
Gb251_7 ns251 0 ni7 0 -0.507907632755
Gb252_7 ns252 0 ni7 0 -0.0008419118152
Gb253_7 ns253 0 ni7 0 0.487353275945
Gb254_7 ns254 0 ni7 0 -0.453187972971
Gb255_7 ns255 0 ni7 0 -0.179348461456
Gb256_7 ns256 0 ni7 0 -0.267410962593
Gb257_7 ns257 0 ni7 0 -0.408554727547
Gb258_7 ns258 0 ni7 0 -0.398757728834
Gb259_7 ns259 0 ni7 0 -0.0514996397364
Gb260_7 ns260 0 ni7 0 -0.38110118275
Gb261_7 ns261 0 ni7 0 0.0928824121159
Gb262_7 ns262 0 ni7 0 -0.328038226621
Gb263_7 ns263 0 ni7 0 0.00951467455824
Gb264_7 ns264 0 ni7 0 -0.273688132867
Gb265_7 ns265 0 ni7 0 0.104515066725
Gb266_7 ns266 0 ni7 0 0.021639783359
Gb267_7 ns267 0 ni7 0 0.291962388554
Gb268_7 ns268 0 ni7 0 0.228255995922
Gb269_7 ns269 0 ni7 0 -0.00230804590343
Gb270_7 ns270 0 ni7 0 -0.0353048726126
Gb271_7 ns271 0 ni7 0 -0.195375857914
Gb272_7 ns272 0 ni7 0 0.158298219061
Gb273_7 ns273 0 ni7 0 -0.0538606771897
Gb274_7 ns274 0 ni7 0 -0.125266532438
Gb275_7 ns275 0 ni7 0 0.0119157039555
Gb276_7 ns276 0 ni7 0 0.0397996579039
Gb277_7 ns277 0 ni7 0 0.0939195913421
Gb278_7 ns278 0 ni7 0 0.0237488618908
Gb279_7 ns279 0 ni7 0 -0.092830123943
Gb280_7 ns280 0 ni7 0 0.00194300457983
Gb281_7 ns281 0 ni7 0 -0.0625301041856
Gb282_7 ns282 0 ni7 0 -0.0395543648239
Gb283_7 ns283 0 ni7 0 -0.0106135674783
Gb284_7 ns284 0 ni7 0 0.0323995666203
Gb285_7 ns285 0 ni7 0 4.14285061595e-05
Gb286_7 ns286 0 ni7 0 -3.6782420325e-05
Gb287_7 ns287 0 ni7 0 0.000451936360429
Gb288_8 ns288 0 ni8 0 16.6816818131
Gb289_8 ns289 0 ni8 0 1.39937119067
Gb290_8 ns290 0 ni8 0 -0.838313186945
Gb291_8 ns291 0 ni8 0 0.178221203364
Gb292_8 ns292 0 ni8 0 -0.507907632755
Gb293_8 ns293 0 ni8 0 -0.0008419118152
Gb294_8 ns294 0 ni8 0 0.487353275945
Gb295_8 ns295 0 ni8 0 -0.453187972971
Gb296_8 ns296 0 ni8 0 -0.179348461456
Gb297_8 ns297 0 ni8 0 -0.267410962593
Gb298_8 ns298 0 ni8 0 -0.408554727547
Gb299_8 ns299 0 ni8 0 -0.398757728834
Gb300_8 ns300 0 ni8 0 -0.0514996397364
Gb301_8 ns301 0 ni8 0 -0.38110118275
Gb302_8 ns302 0 ni8 0 0.0928824121159
Gb303_8 ns303 0 ni8 0 -0.328038226621
Gb304_8 ns304 0 ni8 0 0.00951467455824
Gb305_8 ns305 0 ni8 0 -0.273688132867
Gb306_8 ns306 0 ni8 0 0.104515066725
Gb307_8 ns307 0 ni8 0 0.021639783359
Gb308_8 ns308 0 ni8 0 0.291962388554
Gb309_8 ns309 0 ni8 0 0.228255995922
Gb310_8 ns310 0 ni8 0 -0.00230804590343
Gb311_8 ns311 0 ni8 0 -0.0353048726126
Gb312_8 ns312 0 ni8 0 -0.195375857914
Gb313_8 ns313 0 ni8 0 0.158298219061
Gb314_8 ns314 0 ni8 0 -0.0538606771897
Gb315_8 ns315 0 ni8 0 -0.125266532438
Gb316_8 ns316 0 ni8 0 0.0119157039555
Gb317_8 ns317 0 ni8 0 0.0397996579039
Gb318_8 ns318 0 ni8 0 0.0939195913421
Gb319_8 ns319 0 ni8 0 0.0237488618908
Gb320_8 ns320 0 ni8 0 -0.092830123943
Gb321_8 ns321 0 ni8 0 0.00194300457983
Gb322_8 ns322 0 ni8 0 -0.0625301041856
Gb323_8 ns323 0 ni8 0 -0.0395543648239
Gb324_8 ns324 0 ni8 0 -0.0106135674783
Gb325_8 ns325 0 ni8 0 0.0323995666203
Gb326_8 ns326 0 ni8 0 4.14285061595e-05
Gb327_8 ns327 0 ni8 0 -3.6782420325e-05
Gb328_8 ns328 0 ni8 0 0.000451936360429

Gc1_1 0 n2 ns1 0 0.000653604985242
Gc1_2 0 n2 ns2 0 0.000192136107788
Gc1_3 0 n2 ns3 0 0.0161611294191
Gc1_4 0 n2 ns4 0 -3.55966369229e-05
Gc1_5 0 n2 ns5 0 0.00013302302089
Gc1_6 0 n2 ns6 0 1.58608941634e-05
Gc1_7 0 n2 ns7 0 4.25091425612e-05
Gc1_8 0 n2 ns8 0 0.00039843416145
Gc1_9 0 n2 ns9 0 -0.000728123913372
Gc1_10 0 n2 ns10 0 -0.000395609974197
Gc1_11 0 n2 ns11 0 -0.000250300129712
Gc1_12 0 n2 ns12 0 -0.000754179443113
Gc1_13 0 n2 ns13 0 -0.00169504059307
Gc1_14 0 n2 ns14 0 -0.000489541877683
Gc1_15 0 n2 ns15 0 0.000197577886967
Gc1_16 0 n2 ns16 0 -0.00220965986197
Gc1_17 0 n2 ns17 0 0.000662238248014
Gc1_18 0 n2 ns18 0 0.000952047377324
Gc1_19 0 n2 ns19 0 -0.000609152822865
Gc1_20 0 n2 ns20 0 5.61626794087e-05
Gc1_21 0 n2 ns21 0 0.000914544651991
Gc1_22 0 n2 ns22 0 0.00288245828959
Gc1_23 0 n2 ns23 0 -0.000475827166733
Gc1_24 0 n2 ns24 0 -0.000240176113381
Gc1_25 0 n2 ns25 0 -0.00135291465125
Gc1_26 0 n2 ns26 0 -0.000640073975495
Gc1_27 0 n2 ns27 0 -6.62522232183e-06
Gc1_28 0 n2 ns28 0 -0.00433601505131
Gc1_29 0 n2 ns29 0 0.00196034758537
Gc1_30 0 n2 ns30 0 0.000183979615618
Gc1_31 0 n2 ns31 0 0.00198195901661
Gc1_32 0 n2 ns32 0 0.00164284397527
Gc1_33 0 n2 ns33 0 9.71858993858e-05
Gc1_34 0 n2 ns34 0 2.3461920053e-08
Gc1_35 0 n2 ns35 0 -5.11605646961e-08
Gc1_36 0 n2 ns36 0 -0.00352841210908
Gc1_37 0 n2 ns37 0 -0.00225723924961
Gc1_38 0 n2 ns38 0 0.00843224173188
Gc1_39 0 n2 ns39 0 5.53340404641e-05
Gc1_40 0 n2 ns40 0 -4.41434127952e-05
Gc1_41 0 n2 ns41 0 -4.75574509797e-05
Gc1_42 0 n2 ns42 0 0.000509417366594
Gc1_43 0 n2 ns43 0 -4.10114042429e-05
Gc1_44 0 n2 ns44 0 0.0154794270178
Gc1_45 0 n2 ns45 0 -0.000235565806023
Gc1_46 0 n2 ns46 0 -0.000111649582208
Gc1_47 0 n2 ns47 0 1.14325790834e-05
Gc1_48 0 n2 ns48 0 6.00608124347e-05
Gc1_49 0 n2 ns49 0 0.000333801209038
Gc1_50 0 n2 ns50 0 -0.000693306641878
Gc1_51 0 n2 ns51 0 -0.000174227550107
Gc1_52 0 n2 ns52 0 -0.000231472215703
Gc1_53 0 n2 ns53 0 -0.000662232333353
Gc1_54 0 n2 ns54 0 -0.00112175286436
Gc1_55 0 n2 ns55 0 -0.000623431135343
Gc1_56 0 n2 ns56 0 0.000227506340071
Gc1_57 0 n2 ns57 0 -0.00149418649244
Gc1_58 0 n2 ns58 0 0.000190778292277
Gc1_59 0 n2 ns59 0 0.000521494356599
Gc1_60 0 n2 ns60 0 0.000109198022453
Gc1_61 0 n2 ns61 0 6.14167947799e-05
Gc1_62 0 n2 ns62 0 0.00107684530852
Gc1_63 0 n2 ns63 0 0.00206252691465
Gc1_64 0 n2 ns64 0 -0.000164973562382
Gc1_65 0 n2 ns65 0 -0.000289586640367
Gc1_66 0 n2 ns66 0 -0.00156146103104
Gc1_67 0 n2 ns67 0 -0.000375781051817
Gc1_68 0 n2 ns68 0 -0.000225520466349
Gc1_69 0 n2 ns69 0 -0.00345521353081
Gc1_70 0 n2 ns70 0 0.00195550345476
Gc1_71 0 n2 ns71 0 0.000211367146018
Gc1_72 0 n2 ns72 0 0.00222181513603
Gc1_73 0 n2 ns73 0 0.00154061539658
Gc1_74 0 n2 ns74 0 0.000160290569522
Gc1_75 0 n2 ns75 0 -4.46141704512e-09
Gc1_76 0 n2 ns76 0 -2.43776967685e-08
Gc1_77 0 n2 ns77 0 -0.00295990707308
Gc1_78 0 n2 ns78 0 -0.00134045294129
Gc1_79 0 n2 ns79 0 0.00819671610864
Gc1_80 0 n2 ns80 0 2.9342722335e-05
Gc1_81 0 n2 ns81 0 -1.73606003723e-05
Gc1_82 0 n2 ns82 0 -2.95139351393e-05
Gc1_83 0 n2 ns83 0 0.00031091167289
Gc1_84 0 n2 ns84 0 -0.000617407794152
Gc1_85 0 n2 ns85 0 0.00210831519762
Gc1_86 0 n2 ns86 0 -0.000280268285334
Gc1_87 0 n2 ns87 0 -6.88405600277e-05
Gc1_88 0 n2 ns88 0 3.32399573489e-05
Gc1_89 0 n2 ns89 0 1.34257300343e-05
Gc1_90 0 n2 ns90 0 -0.00052181893565
Gc1_91 0 n2 ns91 0 -0.000442014539715
Gc1_92 0 n2 ns92 0 0.000528118579976
Gc1_93 0 n2 ns93 0 5.90663698967e-07
Gc1_94 0 n2 ns94 0 -0.000198443976919
Gc1_95 0 n2 ns95 0 0.00192304822729
Gc1_96 0 n2 ns96 0 -0.000566304014058
Gc1_97 0 n2 ns97 0 0.00012256760803
Gc1_98 0 n2 ns98 0 0.00202026080037
Gc1_99 0 n2 ns99 0 -0.00102483193814
Gc1_100 0 n2 ns100 0 -0.000854051849339
Gc1_101 0 n2 ns101 0 0.00245268348307
Gc1_102 0 n2 ns102 0 3.05914221872e-05
Gc1_103 0 n2 ns103 0 0.000962184330227
Gc1_104 0 n2 ns104 0 -0.00297097634104
Gc1_105 0 n2 ns105 0 0.000379371109319
Gc1_106 0 n2 ns106 0 -0.00028324044423
Gc1_107 0 n2 ns107 0 -0.00130680238245
Gc1_108 0 n2 ns108 0 0.000546654711095
Gc1_109 0 n2 ns109 0 -0.000297402700323
Gc1_110 0 n2 ns110 0 0.00461950741709
Gc1_111 0 n2 ns111 0 -0.0001439513568
Gc1_112 0 n2 ns112 0 -6.79590692418e-06
Gc1_113 0 n2 ns113 0 0.00211122912177
Gc1_114 0 n2 ns114 0 0.000735630706629
Gc1_115 0 n2 ns115 0 -0.00159120806586
Gc1_116 0 n2 ns116 0 -7.68858076876e-08
Gc1_117 0 n2 ns117 0 7.6291707138e-08
Gc1_118 0 n2 ns118 0 0.00365912823775
Gc1_119 0 n2 ns119 0 -0.00129730799691
Gc1_120 0 n2 ns120 0 0.00410036989295
Gc1_121 0 n2 ns121 0 -9.49898222732e-05
Gc1_122 0 n2 ns122 0 7.84699837452e-05
Gc1_123 0 n2 ns123 0 3.67782224181e-05
Gc1_124 0 n2 ns124 0 0.00118894876428
Gc1_125 0 n2 ns125 0 -0.000676916221985
Gc1_126 0 n2 ns126 0 0.0110574898831
Gc1_127 0 n2 ns127 0 -0.000623359645595
Gc1_128 0 n2 ns128 0 -0.000348849163776
Gc1_129 0 n2 ns129 0 3.20295749607e-05
Gc1_130 0 n2 ns130 0 6.15035459955e-05
Gc1_131 0 n2 ns131 0 -2.12540085183e-05
Gc1_132 0 n2 ns132 0 -0.00058198001475
Gc1_133 0 n2 ns133 0 0.00040370252455
Gc1_134 0 n2 ns134 0 -6.63844897679e-05
Gc1_135 0 n2 ns135 0 -0.000944838684617
Gc1_136 0 n2 ns136 0 0.000784345143752
Gc1_137 0 n2 ns137 0 -0.000645758963401
Gc1_138 0 n2 ns138 0 0.000170130812779
Gc1_139 0 n2 ns139 0 0.00111523913078
Gc1_140 0 n2 ns140 0 -0.000433299120747
Gc1_141 0 n2 ns141 0 -0.00171856089915
Gc1_142 0 n2 ns142 0 0.00231266061956
Gc1_143 0 n2 ns143 0 3.09075577578e-05
Gc1_144 0 n2 ns144 0 0.00115021921212
Gc1_145 0 n2 ns145 0 -0.00182175818101
Gc1_146 0 n2 ns146 0 -0.000478204074569
Gc1_147 0 n2 ns147 0 -0.000420842603262
Gc1_148 0 n2 ns148 0 -0.00152062114864
Gc1_149 0 n2 ns149 0 0.00131425885638
Gc1_150 0 n2 ns150 0 -0.000326310967382
Gc1_151 0 n2 ns151 0 0.00250079986343
Gc1_152 0 n2 ns152 0 0.00098150120415
Gc1_153 0 n2 ns153 0 0.000284041659812
Gc1_154 0 n2 ns154 0 0.00237887190633
Gc1_155 0 n2 ns155 0 -0.000964477052103
Gc1_156 0 n2 ns156 0 -0.00199117315295
Gc1_157 0 n2 ns157 0 -4.97420594703e-08
Gc1_158 0 n2 ns158 0 9.21955827619e-08
Gc1_159 0 n2 ns159 0 0.00327616540424
Gc1_160 0 n2 ns160 0 -0.000893711872108
Gc1_161 0 n2 ns161 0 0.00500601606982
Gc1_162 0 n2 ns162 0 -0.000132083028115
Gc1_163 0 n2 ns163 0 0.00011931213272
Gc1_164 0 n2 ns164 0 4.21153676267e-05
Gc1_165 0 n2 ns165 0 -0.000322992498164
Gc1_166 0 n2 ns166 0 0.00121079941865
Gc1_167 0 n2 ns167 0 0.00203083274041
Gc1_168 0 n2 ns168 0 0.000239347633673
Gc1_169 0 n2 ns169 0 -0.000413648364136
Gc1_170 0 n2 ns170 0 -1.87116727315e-05
Gc1_171 0 n2 ns171 0 2.56660642084e-05
Gc1_172 0 n2 ns172 0 0.00065812194839
Gc1_173 0 n2 ns173 0 -0.000710309800897
Gc1_174 0 n2 ns174 0 0.000463646734132
Gc1_175 0 n2 ns175 0 0.000150389752658
Gc1_176 0 n2 ns176 0 2.28895396065e-05
Gc1_177 0 n2 ns177 0 0.00366254488857
Gc1_178 0 n2 ns178 0 0.000598822461919
Gc1_179 0 n2 ns179 0 -0.000235857081027
Gc1_180 0 n2 ns180 0 -0.00205496700146
Gc1_181 0 n2 ns181 0 0.000167887358975
Gc1_182 0 n2 ns182 0 -0.00107283235975
Gc1_183 0 n2 ns183 0 -0.00873147945809
Gc1_184 0 n2 ns184 0 6.78027936751e-05
Gc1_185 0 n2 ns185 0 0.000820861683732
Gc1_186 0 n2 ns186 0 -0.00360753947395
Gc1_187 0 n2 ns187 0 -0.000242586207998
Gc1_188 0 n2 ns188 0 0.000118807667742
Gc1_189 0 n2 ns189 0 0.00148780001584
Gc1_190 0 n2 ns190 0 0.00230778306903
Gc1_191 0 n2 ns191 0 -0.00322170866659
Gc1_192 0 n2 ns192 0 -0.00950201884859
Gc1_193 0 n2 ns193 0 -0.00349161427638
Gc1_194 0 n2 ns194 0 0.000466911470309
Gc1_195 0 n2 ns195 0 0.00323976279313
Gc1_196 0 n2 ns196 0 0.00440658191505
Gc1_197 0 n2 ns197 0 -0.0100823556574
Gc1_198 0 n2 ns198 0 -2.14070143043e-07
Gc1_199 0 n2 ns199 0 3.72242721426e-08
Gc1_200 0 n2 ns200 0 0.00839546283975
Gc1_201 0 n2 ns201 0 0.00649601246276
Gc1_202 0 n2 ns202 0 -0.0112442593235
Gc1_203 0 n2 ns203 0 -0.000171659470034
Gc1_204 0 n2 ns204 0 0.000176355968398
Gc1_205 0 n2 ns205 0 7.82761867979e-05
Gc1_206 0 n2 ns206 0 0.000129489173764
Gc1_207 0 n2 ns207 0 -0.000269648919579
Gc1_208 0 n2 ns208 0 0.00371902788511
Gc1_209 0 n2 ns209 0 -0.000714357936034
Gc1_210 0 n2 ns210 0 -0.00012980463575
Gc1_211 0 n2 ns211 0 8.16105488341e-05
Gc1_212 0 n2 ns212 0 5.70633213323e-05
Gc1_213 0 n2 ns213 0 -0.000744792313413
Gc1_214 0 n2 ns214 0 -0.00133965091802
Gc1_215 0 n2 ns215 0 0.000732360787355
Gc1_216 0 n2 ns216 0 -0.000142450203782
Gc1_217 0 n2 ns217 0 -0.000379192264074
Gc1_218 0 n2 ns218 0 -0.00236207716754
Gc1_219 0 n2 ns219 0 0.000668077300657
Gc1_220 0 n2 ns220 0 -0.000123432273375
Gc1_221 0 n2 ns221 0 -0.00170806728808
Gc1_222 0 n2 ns222 0 0.000644736403657
Gc1_223 0 n2 ns223 0 -0.000792624226082
Gc1_224 0 n2 ns224 0 0.00902109108843
Gc1_225 0 n2 ns225 0 2.99212776946e-05
Gc1_226 0 n2 ns226 0 0.00112254622476
Gc1_227 0 n2 ns227 0 -0.00121377736193
Gc1_228 0 n2 ns228 0 0.000895049429075
Gc1_229 0 n2 ns229 0 0.000331214685896
Gc1_230 0 n2 ns230 0 0.00143144166472
Gc1_231 0 n2 ns231 0 -0.00180690870866
Gc1_232 0 n2 ns232 0 0.00203602157206
Gc1_233 0 n2 ns233 0 2.11484268752e-06
Gc1_234 0 n2 ns234 0 0.00597784861289
Gc1_235 0 n2 ns235 0 2.71194354382e-06
Gc1_236 0 n2 ns236 0 0.00150016479067
Gc1_237 0 n2 ns237 0 -0.00199795512919
Gc1_238 0 n2 ns238 0 0.00588831517404
Gc1_239 0 n2 ns239 0 7.03903895402e-08
Gc1_240 0 n2 ns240 0 5.69689876866e-08
Gc1_241 0 n2 ns241 0 -0.00170578868761
Gc1_242 0 n2 ns242 0 -0.0056954856494
Gc1_243 0 n2 ns243 0 -0.00380621505782
Gc1_244 0 n2 ns244 0 9.79074928358e-06
Gc1_245 0 n2 ns245 0 3.57343931556e-07
Gc1_246 0 n2 ns246 0 -1.96093829331e-05
Gc1_247 0 n2 ns247 0 -0.000164789795134
Gc1_248 0 n2 ns248 0 0.00225479905169
Gc1_249 0 n2 ns249 0 0.0024965882299
Gc1_250 0 n2 ns250 0 0.000255505816644
Gc1_251 0 n2 ns251 0 0.000598839374675
Gc1_252 0 n2 ns252 0 2.87394986455e-05
Gc1_253 0 n2 ns253 0 -9.40368868693e-06
Gc1_254 0 n2 ns254 0 0.000230669085295
Gc1_255 0 n2 ns255 0 -0.000146086581838
Gc1_256 0 n2 ns256 0 -0.000530876068632
Gc1_257 0 n2 ns257 0 -0.000187631378316
Gc1_258 0 n2 ns258 0 -0.00118079987055
Gc1_259 0 n2 ns259 0 -0.000641558812026
Gc1_260 0 n2 ns260 0 0.000693286737067
Gc1_261 0 n2 ns261 0 -0.000122300840187
Gc1_262 0 n2 ns262 0 0.00206095269167
Gc1_263 0 n2 ns263 0 -0.00131207363365
Gc1_264 0 n2 ns264 0 -0.00200806849747
Gc1_265 0 n2 ns265 0 -0.000315648791604
Gc1_266 0 n2 ns266 0 -8.25134113727e-06
Gc1_267 0 n2 ns267 0 0.000936197621045
Gc1_268 0 n2 ns268 0 0.00341868915217
Gc1_269 0 n2 ns269 0 -0.000811476940334
Gc1_270 0 n2 ns270 0 0.00013212213496
Gc1_271 0 n2 ns271 0 0.00131840896138
Gc1_272 0 n2 ns272 0 0.000797156528955
Gc1_273 0 n2 ns273 0 -0.00122822212497
Gc1_274 0 n2 ns274 0 0.00396331299848
Gc1_275 0 n2 ns275 0 0.000327001253976
Gc1_276 0 n2 ns276 0 0.000183650378541
Gc1_277 0 n2 ns277 0 0.00203080972008
Gc1_278 0 n2 ns278 0 0.00030072511871
Gc1_279 0 n2 ns279 0 -0.00132002365855
Gc1_280 0 n2 ns280 0 -4.36399307026e-08
Gc1_281 0 n2 ns281 0 5.67319397418e-08
Gc1_282 0 n2 ns282 0 -0.00321547353649
Gc1_283 0 n2 ns283 0 -0.00239322074869
Gc1_284 0 n2 ns284 0 -0.00152042536271
Gc1_285 0 n2 ns285 0 7.1337956714e-05
Gc1_286 0 n2 ns286 0 -3.68791428127e-05
Gc1_287 0 n2 ns287 0 -5.01194790319e-05
Gc1_288 0 n2 ns288 0 0.000129200501603
Gc1_289 0 n2 ns289 0 0.00143812142506
Gc1_290 0 n2 ns290 0 0.00311200563035
Gc1_291 0 n2 ns291 0 -4.26651064766e-05
Gc1_292 0 n2 ns292 0 0.000608576754077
Gc1_293 0 n2 ns293 0 5.73045104297e-05
Gc1_294 0 n2 ns294 0 -3.06422370402e-06
Gc1_295 0 n2 ns295 0 -0.000278368706478
Gc1_296 0 n2 ns296 0 -0.000249742804885
Gc1_297 0 n2 ns297 0 -0.000259921656958
Gc1_298 0 n2 ns298 0 -0.00029591587534
Gc1_299 0 n2 ns299 0 -0.00142228824628
Gc1_300 0 n2 ns300 0 -0.00118896358902
Gc1_301 0 n2 ns301 0 0.000780977885972
Gc1_302 0 n2 ns302 0 -0.000142897167849
Gc1_303 0 n2 ns303 0 0.00141261260301
Gc1_304 0 n2 ns304 0 -0.00060248863687
Gc1_305 0 n2 ns305 0 -0.000642241279736
Gc1_306 0 n2 ns306 0 0.00211782752024
Gc1_307 0 n2 ns307 0 2.07763608635e-05
Gc1_308 0 n2 ns308 0 0.0010996092254
Gc1_309 0 n2 ns309 0 0.00259324446154
Gc1_310 0 n2 ns310 0 -0.000337708098363
Gc1_311 0 n2 ns311 0 0.000216904090981
Gc1_312 0 n2 ns312 0 0.00151912861142
Gc1_313 0 n2 ns313 0 0.000279864185846
Gc1_314 0 n2 ns314 0 -0.000313665091954
Gc1_315 0 n2 ns315 0 0.0037593064782
Gc1_316 0 n2 ns316 0 0.00186962201902
Gc1_317 0 n2 ns317 0 9.81348974527e-05
Gc1_318 0 n2 ns318 0 0.00212260740484
Gc1_319 0 n2 ns319 0 2.76921910136e-05
Gc1_320 0 n2 ns320 0 0.00069619695359
Gc1_321 0 n2 ns321 0 -2.34484506872e-08
Gc1_322 0 n2 ns322 0 6.80245507091e-08
Gc1_323 0 n2 ns323 0 -0.00338289572517
Gc1_324 0 n2 ns324 0 -0.00298608890181
Gc1_325 0 n2 ns325 0 -0.00267421529966
Gc1_326 0 n2 ns326 0 5.16786442218e-05
Gc1_327 0 n2 ns327 0 -1.84698872915e-05
Gc1_328 0 n2 ns328 0 -4.67016330071e-05
Gd1_1 0 n2 ni1 0 -0.00204503999796
Gd1_2 0 n2 ni2 0 -0.00204737524974
Gd1_3 0 n2 ni3 0 -0.000972172368451
Gd1_4 0 n2 ni4 0 -0.00323933071796
Gd1_5 0 n2 ni5 0 7.49367439409e-05
Gd1_6 0 n2 ni6 0 -0.000656344066583
Gd1_7 0 n2 ni7 0 0.000742357141636
Gd1_8 0 n2 ni8 0 0.000148002286291
Gc2_1 0 n4 ns1 0 0.000509417364437
Gc2_2 0 n4 ns2 0 -4.10114122495e-05
Gc2_3 0 n4 ns3 0 0.0154794270151
Gc2_4 0 n4 ns4 0 -0.00023556580523
Gc2_5 0 n4 ns5 0 -0.000111649579014
Gc2_6 0 n4 ns6 0 1.14325800398e-05
Gc2_7 0 n4 ns7 0 6.00608122008e-05
Gc2_8 0 n4 ns8 0 0.000333801212006
Gc2_9 0 n4 ns9 0 -0.000693306644567
Gc2_10 0 n4 ns10 0 -0.000174227548285
Gc2_11 0 n4 ns11 0 -0.000231472215912
Gc2_12 0 n4 ns12 0 -0.000662232339173
Gc2_13 0 n4 ns13 0 -0.00112175287174
Gc2_14 0 n4 ns14 0 -0.000623431134907
Gc2_15 0 n4 ns15 0 0.000227506340754
Gc2_16 0 n4 ns16 0 -0.0014941864927
Gc2_17 0 n4 ns17 0 0.000190778289638
Gc2_18 0 n4 ns18 0 0.000521494343562
Gc2_19 0 n4 ns19 0 0.000109198025528
Gc2_20 0 n4 ns20 0 6.14167942771e-05
Gc2_21 0 n4 ns21 0 0.00107684530847
Gc2_22 0 n4 ns22 0 0.00206252691819
Gc2_23 0 n4 ns23 0 -0.000164973562246
Gc2_24 0 n4 ns24 0 -0.000289586641328
Gc2_25 0 n4 ns25 0 -0.00156146103152
Gc2_26 0 n4 ns26 0 -0.000375781047878
Gc2_27 0 n4 ns27 0 -0.000225520469882
Gc2_28 0 n4 ns28 0 -0.00345521353148
Gc2_29 0 n4 ns29 0 0.00195550345585
Gc2_30 0 n4 ns30 0 0.000211367144459
Gc2_31 0 n4 ns31 0 0.00222181513682
Gc2_32 0 n4 ns32 0 0.0015406153982
Gc2_33 0 n4 ns33 0 0.000160290561847
Gc2_34 0 n4 ns34 0 -4.46141745935e-09
Gc2_35 0 n4 ns35 0 -2.43776964888e-08
Gc2_36 0 n4 ns36 0 -0.00295990706839
Gc2_37 0 n4 ns37 0 -0.00134045296852
Gc2_38 0 n4 ns38 0 0.00819671612917
Gc2_39 0 n4 ns39 0 2.93427235738e-05
Gc2_40 0 n4 ns40 0 -1.73606037585e-05
Gc2_41 0 n4 ns41 0 -2.9513935581e-05
Gc2_42 0 n4 ns42 0 -0.000248495935087
Gc2_43 0 n4 ns43 0 0.000315913700735
Gc2_44 0 n4 ns44 0 0.011026534282
Gc2_45 0 n4 ns45 0 0.000132265003844
Gc2_46 0 n4 ns46 0 0.000199268110066
Gc2_47 0 n4 ns47 0 3.64751440301e-05
Gc2_48 0 n4 ns48 0 3.29643776283e-05
Gc2_49 0 n4 ns49 0 0.000203574120054
Gc2_50 0 n4 ns50 0 -0.000748898011047
Gc2_51 0 n4 ns51 0 -2.23549390395e-05
Gc2_52 0 n4 ns52 0 -0.00017304118216
Gc2_53 0 n4 ns53 0 -0.000372803682598
Gc2_54 0 n4 ns54 0 -0.00113624109709
Gc2_55 0 n4 ns55 0 -0.000788893201355
Gc2_56 0 n4 ns56 0 0.000281790305379
Gc2_57 0 n4 ns57 0 -0.000980421527287
Gc2_58 0 n4 ns58 0 -1.13457334939e-05
Gc2_59 0 n4 ns59 0 0.000114699123779
Gc2_60 0 n4 ns60 0 -0.000288659377239
Gc2_61 0 n4 ns61 0 7.90671066643e-05
Gc2_62 0 n4 ns62 0 0.00125652666392
Gc2_63 0 n4 ns63 0 0.00134604147589
Gc2_64 0 n4 ns64 0 -8.46314724406e-05
Gc2_65 0 n4 ns65 0 -0.0002758034735
Gc2_66 0 n4 ns66 0 -0.00180421744719
Gc2_67 0 n4 ns67 0 3.70926198308e-05
Gc2_68 0 n4 ns68 0 0.000293344102337
Gc2_69 0 n4 ns69 0 -0.00251295869517
Gc2_70 0 n4 ns70 0 0.00121207722228
Gc2_71 0 n4 ns71 0 0.000244961369471
Gc2_72 0 n4 ns72 0 0.0029167996011
Gc2_73 0 n4 ns73 0 0.000739439893904
Gc2_74 0 n4 ns74 0 -0.000967641159468
Gc2_75 0 n4 ns75 0 -5.49062729853e-08
Gc2_76 0 n4 ns76 0 -1.22505895236e-07
Gc2_77 0 n4 ns77 0 -0.00153803503974
Gc2_78 0 n4 ns78 0 -0.00143307343405
Gc2_79 0 n4 ns79 0 0.00883323900077
Gc2_80 0 n4 ns80 0 8.85835395416e-05
Gc2_81 0 n4 ns81 0 -5.77902102326e-05
Gc2_82 0 n4 ns82 0 -4.5478126664e-05
Gc2_83 0 n4 ns83 0 0.00120082231385
Gc2_84 0 n4 ns84 0 -0.000672266381463
Gc2_85 0 n4 ns85 0 0.0110071498882
Gc2_86 0 n4 ns86 0 -0.000626987869014
Gc2_87 0 n4 ns87 0 -0.000362671547917
Gc2_88 0 n4 ns88 0 2.95357610126e-05
Gc2_89 0 n4 ns89 0 6.14001558011e-05
Gc2_90 0 n4 ns90 0 -2.78461243646e-05
Gc2_91 0 n4 ns91 0 -0.000569945748668
Gc2_92 0 n4 ns92 0 0.000392325643952
Gc2_93 0 n4 ns93 0 -6.35586177674e-05
Gc2_94 0 n4 ns94 0 -0.000915872543139
Gc2_95 0 n4 ns95 0 0.000807216164423
Gc2_96 0 n4 ns96 0 -0.000644933725985
Gc2_97 0 n4 ns97 0 0.000165210660964
Gc2_98 0 n4 ns98 0 0.00112057722853
Gc2_99 0 n4 ns99 0 -0.000412953982667
Gc2_100 0 n4 ns100 0 -0.00168227478152
Gc2_101 0 n4 ns101 0 0.00227949137984
Gc2_102 0 n4 ns102 0 2.88193688839e-05
Gc2_103 0 n4 ns103 0 0.00114430998054
Gc2_104 0 n4 ns104 0 -0.00183249646421
Gc2_105 0 n4 ns105 0 -0.000491925364093
Gc2_106 0 n4 ns106 0 -0.000411746471974
Gc2_107 0 n4 ns107 0 -0.00151364334657
Gc2_108 0 n4 ns108 0 0.00129229854888
Gc2_109 0 n4 ns109 0 -0.000307728429749
Gc2_110 0 n4 ns110 0 0.0025345572764
Gc2_111 0 n4 ns111 0 0.000985415837567
Gc2_112 0 n4 ns112 0 0.000272855985537
Gc2_113 0 n4 ns113 0 0.00237761971851
Gc2_114 0 n4 ns114 0 -0.000928584080853
Gc2_115 0 n4 ns115 0 -0.00197826367811
Gc2_116 0 n4 ns116 0 -4.98398075081e-08
Gc2_117 0 n4 ns117 0 9.01777676549e-08
Gc2_118 0 n4 ns118 0 0.00329828873381
Gc2_119 0 n4 ns119 0 -0.000880741775934
Gc2_120 0 n4 ns120 0 0.00500374263549
Gc2_121 0 n4 ns121 0 -0.000132046681154
Gc2_122 0 n4 ns122 0 0.00012181044622
Gc2_123 0 n4 ns123 0 4.20282947938e-05
Gc2_124 0 n4 ns124 0 0.000671636707144
Gc2_125 0 n4 ns125 0 -0.000321839690563
Gc2_126 0 n4 ns126 0 0.00971084027949
Gc2_127 0 n4 ns127 0 -0.00035540527319
Gc2_128 0 n4 ns128 0 -7.35659618859e-05
Gc2_129 0 n4 ns129 0 2.49026419308e-05
Gc2_130 0 n4 ns130 0 3.88222341397e-05
Gc2_131 0 n4 ns131 0 -0.000189732765334
Gc2_132 0 n4 ns132 0 -0.000800844742877
Gc2_133 0 n4 ns133 0 0.000274833522625
Gc2_134 0 n4 ns134 0 -8.40250401894e-05
Gc2_135 0 n4 ns135 0 -0.000765891827576
Gc2_136 0 n4 ns136 0 0.000922145139069
Gc2_137 0 n4 ns137 0 -0.000762424559896
Gc2_138 0 n4 ns138 0 0.000223423049076
Gc2_139 0 n4 ns139 0 0.00080422625429
Gc2_140 0 n4 ns140 0 -0.00038544313949
Gc2_141 0 n4 ns141 0 -0.00020977064347
Gc2_142 0 n4 ns142 0 0.00215591625586
Gc2_143 0 n4 ns143 0 4.16486505881e-05
Gc2_144 0 n4 ns144 0 0.00129074572478
Gc2_145 0 n4 ns145 0 -0.00140746161631
Gc2_146 0 n4 ns146 0 -0.000128905802284
Gc2_147 0 n4 ns147 0 -0.000319782056858
Gc2_148 0 n4 ns148 0 -0.00174618237992
Gc2_149 0 n4 ns149 0 4.58637529379e-05
Gc2_150 0 n4 ns150 0 -0.00056907046235
Gc2_151 0 n4 ns151 0 0.00218788037101
Gc2_152 0 n4 ns152 0 0.0015377759014
Gc2_153 0 n4 ns153 0 8.59639716377e-05
Gc2_154 0 n4 ns154 0 0.0025792405109
Gc2_155 0 n4 ns155 0 0.00137403887775
Gc2_156 0 n4 ns156 0 -0.000114557140182
Gc2_157 0 n4 ns157 0 -6.49722725287e-09
Gc2_158 0 n4 ns158 0 2.97776962209e-08
Gc2_159 0 n4 ns159 0 0.00149377883045
Gc2_160 0 n4 ns160 0 -0.000183128055622
Gc2_161 0 n4 ns161 0 0.00612151303666
Gc2_162 0 n4 ns162 0 -4.33871914597e-05
Gc2_163 0 n4 ns163 0 2.47057975025e-05
Gc2_164 0 n4 ns164 0 1.8875750893e-05
Gc2_165 0 n4 ns165 0 0.000132934058178
Gc2_166 0 n4 ns166 0 -0.000257149770987
Gc2_167 0 n4 ns167 0 0.00371549143329
Gc2_168 0 n4 ns168 0 -0.000719470011768
Gc2_169 0 n4 ns169 0 -0.000141524833912
Gc2_170 0 n4 ns170 0 8.05254446005e-05
Gc2_171 0 n4 ns171 0 5.75435507903e-05
Gc2_172 0 n4 ns172 0 -0.00074825671214
Gc2_173 0 n4 ns173 0 -0.00132691991945
Gc2_174 0 n4 ns174 0 0.000726677375073
Gc2_175 0 n4 ns175 0 -0.000135228052615
Gc2_176 0 n4 ns176 0 -0.000344217888292
Gc2_177 0 n4 ns177 0 -0.00236548127786
Gc2_178 0 n4 ns178 0 0.00066575292158
Gc2_179 0 n4 ns179 0 -0.000123573553557
Gc2_180 0 n4 ns180 0 -0.00169983824842
Gc2_181 0 n4 ns181 0 0.000644176096002
Gc2_182 0 n4 ns182 0 -0.000798459513047
Gc2_183 0 n4 ns183 0 0.00898286058895
Gc2_184 0 n4 ns184 0 3.17028769115e-05
Gc2_185 0 n4 ns185 0 0.00112134101689
Gc2_186 0 n4 ns186 0 -0.00121178421154
Gc2_187 0 n4 ns187 0 0.000906037633053
Gc2_188 0 n4 ns188 0 0.000331291489705
Gc2_189 0 n4 ns189 0 0.00142696441711
Gc2_190 0 n4 ns190 0 -0.0017969907605
Gc2_191 0 n4 ns191 0 0.00203917426912
Gc2_192 0 n4 ns192 0 -1.56534485863e-05
Gc2_193 0 n4 ns193 0 0.00596420703975
Gc2_194 0 n4 ns194 0 8.0546350538e-06
Gc2_195 0 n4 ns195 0 0.00150076010854
Gc2_196 0 n4 ns196 0 -0.00201222868383
Gc2_197 0 n4 ns197 0 0.00587963329035
Gc2_198 0 n4 ns198 0 6.97571881068e-08
Gc2_199 0 n4 ns199 0 5.65858505129e-08
Gc2_200 0 n4 ns200 0 -0.00169605228984
Gc2_201 0 n4 ns201 0 -0.0057208205976
Gc2_202 0 n4 ns202 0 -0.00378575923694
Gc2_203 0 n4 ns203 0 3.3056972215e-06
Gc2_204 0 n4 ns204 0 -6.96919379609e-07
Gc2_205 0 n4 ns205 0 -1.89231257386e-05
Gc2_206 0 n4 ns206 0 -0.000123587857001
Gc2_207 0 n4 ns207 0 0.00193830282717
Gc2_208 0 n4 ns208 0 0.00398252622921
Gc2_209 0 n4 ns209 0 0.000358815171659
Gc2_210 0 n4 ns210 0 -4.07963646885e-05
Gc2_211 0 n4 ns211 0 -2.41004635069e-05
Gc2_212 0 n4 ns212 0 1.22616443061e-05
Gc2_213 0 n4 ns213 0 0.000665376288964
Gc2_214 0 n4 ns214 0 -0.000394280638338
Gc2_215 0 n4 ns215 0 -1.12847387275e-05
Gc2_216 0 n4 ns216 0 0.000114477614724
Gc2_217 0 n4 ns217 0 -0.000941154289835
Gc2_218 0 n4 ns218 0 0.00341705149756
Gc2_219 0 n4 ns219 0 0.000912896961591
Gc2_220 0 n4 ns220 0 -0.000299117190137
Gc2_221 0 n4 ns221 0 -0.000809481190727
Gc2_222 0 n4 ns222 0 -0.000759467738755
Gc2_223 0 n4 ns223 0 -0.000924355782316
Gc2_224 0 n4 ns224 0 -0.00924034032048
Gc2_225 0 n4 ns225 0 6.47362109427e-05
Gc2_226 0 n4 ns226 0 0.00117877912136
Gc2_227 0 n4 ns227 0 -0.00187943357811
Gc2_228 0 n4 ns228 0 -0.000910123033977
Gc2_229 0 n4 ns229 0 8.8462193507e-05
Gc2_230 0 n4 ns230 0 0.00191192274937
Gc2_231 0 n4 ns231 0 0.00307453564704
Gc2_232 0 n4 ns232 0 -0.00352545963566
Gc2_233 0 n4 ns233 0 -0.00797890164847
Gc2_234 0 n4 ns234 0 -0.00413568241879
Gc2_235 0 n4 ns235 0 0.000514530348373
Gc2_236 0 n4 ns236 0 0.00404920676308
Gc2_237 0 n4 ns237 0 0.0042337774257
Gc2_238 0 n4 ns238 0 -0.0107401261705
Gc2_239 0 n4 ns239 0 -1.99104965628e-07
Gc2_240 0 n4 ns240 0 -2.42524395819e-08
Gc2_241 0 n4 ns241 0 0.006768249448
Gc2_242 0 n4 ns242 0 0.00555048008959
Gc2_243 0 n4 ns243 0 -0.0116614758584
Gc2_244 0 n4 ns244 0 -0.00017898644361
Gc2_245 0 n4 ns245 0 0.000187894609029
Gc2_246 0 n4 ns246 0 7.31872321345e-05
Gc2_247 0 n4 ns247 0 0.000120368782078
Gc2_248 0 n4 ns248 0 0.00141761587563
Gc2_249 0 n4 ns249 0 0.00308861965943
Gc2_250 0 n4 ns250 0 -3.81441477505e-05
Gc2_251 0 n4 ns251 0 0.000625993444554
Gc2_252 0 n4 ns252 0 5.95306144097e-05
Gc2_253 0 n4 ns253 0 -3.72215904003e-06
Gc2_254 0 n4 ns254 0 -0.000271030753118
Gc2_255 0 n4 ns255 0 -0.000259157966057
Gc2_256 0 n4 ns256 0 -0.000249159547621
Gc2_257 0 n4 ns257 0 -0.000298273533832
Gc2_258 0 n4 ns258 0 -0.00144072400925
Gc2_259 0 n4 ns259 0 -0.00121085251519
Gc2_260 0 n4 ns260 0 0.000778751340731
Gc2_261 0 n4 ns261 0 -0.000138389216978
Gc2_262 0 n4 ns262 0 0.00140967166966
Gc2_263 0 n4 ns263 0 -0.000599319344376
Gc2_264 0 n4 ns264 0 -0.000689404866969
Gc2_265 0 n4 ns265 0 0.00211955397194
Gc2_266 0 n4 ns266 0 1.51499485381e-05
Gc2_267 0 n4 ns267 0 0.00109400144693
Gc2_268 0 n4 ns268 0 0.002610025788
Gc2_269 0 n4 ns269 0 -0.000328899166004
Gc2_270 0 n4 ns270 0 0.000205365761812
Gc2_271 0 n4 ns271 0 0.00151413033363
Gc2_272 0 n4 ns272 0 0.000290605444412
Gc2_273 0 n4 ns273 0 -0.000346488635224
Gc2_274 0 n4 ns274 0 0.00377593599183
Gc2_275 0 n4 ns275 0 0.00191056100515
Gc2_276 0 n4 ns276 0 8.0235835078e-05
Gc2_277 0 n4 ns277 0 0.00211760692515
Gc2_278 0 n4 ns278 0 5.08624678301e-05
Gc2_279 0 n4 ns279 0 0.000693789443097
Gc2_280 0 n4 ns280 0 -2.33221462182e-08
Gc2_281 0 n4 ns281 0 6.72235289892e-08
Gc2_282 0 n4 ns282 0 -0.00338153929103
Gc2_283 0 n4 ns283 0 -0.00301873063034
Gc2_284 0 n4 ns284 0 -0.00265158118738
Gc2_285 0 n4 ns285 0 5.78361384284e-05
Gc2_286 0 n4 ns286 0 -2.02627151136e-05
Gc2_287 0 n4 ns287 0 -4.90081615509e-05
Gc2_288 0 n4 ns288 0 -3.90347986794e-05
Gc2_289 0 n4 ns289 0 0.00122820107301
Gc2_290 0 n4 ns290 0 0.00405757659509
Gc2_291 0 n4 ns291 0 -0.000331319104966
Gc2_292 0 n4 ns292 0 0.000199835939404
Gc2_293 0 n4 ns293 0 7.20314699405e-05
Gc2_294 0 n4 ns294 0 4.78487984365e-05
Gc2_295 0 n4 ns295 0 -0.000206780541991
Gc2_296 0 n4 ns296 0 -0.000964601405373
Gc2_297 0 n4 ns297 0 3.27091396576e-05
Gc2_298 0 n4 ns298 0 -0.000281784322818
Gc2_299 0 n4 ns299 0 -0.000603584084769
Gc2_300 0 n4 ns300 0 -0.0012759777352
Gc2_301 0 n4 ns301 0 0.000890196989294
Gc2_302 0 n4 ns302 0 -0.000200270455779
Gc2_303 0 n4 ns303 0 0.000751157897664
Gc2_304 0 n4 ns304 0 -0.000378032696002
Gc2_305 0 n4 ns305 0 -0.00266064982639
Gc2_306 0 n4 ns306 0 0.00359040257277
Gc2_307 0 n4 ns307 0 -1.44229066203e-05
Gc2_308 0 n4 ns308 0 0.00126928959719
Gc2_309 0 n4 ns309 0 0.0021135174451
Gc2_310 0 n4 ns310 0 2.15912543198e-05
Gc2_311 0 n4 ns311 0 0.000206268126809
Gc2_312 0 n4 ns312 0 0.00174681852852
Gc2_313 0 n4 ns313 0 -7.60526987061e-05
Gc2_314 0 n4 ns314 0 -0.000355910953321
Gc2_315 0 n4 ns315 0 0.00282796798101
Gc2_316 0 n4 ns316 0 0.00370740084748
Gc2_317 0 n4 ns317 0 0.000169776049563
Gc2_318 0 n4 ns318 0 0.00221879858178
Gc2_319 0 n4 ns319 0 -0.000886144126939
Gc2_320 0 n4 ns320 0 0.0020780352507
Gc2_321 0 n4 ns321 0 4.12072174582e-09
Gc2_322 0 n4 ns322 0 7.61998085824e-08
Gc2_323 0 n4 ns323 0 -0.00354138121619
Gc2_324 0 n4 ns324 0 -0.00360545538135
Gc2_325 0 n4 ns325 0 -0.00370248519825
Gc2_326 0 n4 ns326 0 3.22615122928e-05
Gc2_327 0 n4 ns327 0 -3.45691091363e-06
Gc2_328 0 n4 ns328 0 -4.03762079518e-05
Gd2_1 0 n4 ni1 0 -0.00204737524993
Gd2_2 0 n4 ni2 0 -0.000505479421988
Gd2_3 0 n4 ni3 0 -0.00323133395129
Gd2_4 0 n4 ni4 0 -0.00201358223983
Gd2_5 0 n4 ni5 0 -0.000649234279772
Gd2_6 0 n4 ni6 0 -0.000135924975429
Gd2_7 0 n4 ni7 0 0.000148706111532
Gd2_8 0 n4 ni8 0 -6.68263993596e-05
Gc3_1 0 n6 ns1 0 0.000310911687899
Gc3_2 0 n6 ns2 0 -0.000617407767406
Gc3_3 0 n6 ns3 0 0.00210831519658
Gc3_4 0 n6 ns4 0 -0.000280268292426
Gc3_5 0 n6 ns5 0 -6.88405764518e-05
Gc3_6 0 n6 ns6 0 3.3239953981e-05
Gc3_7 0 n6 ns7 0 1.34257308653e-05
Gc3_8 0 n6 ns8 0 -0.000521818944506
Gc3_9 0 n6 ns9 0 -0.000442014527029
Gc3_10 0 n6 ns10 0 0.000528118572467
Gc3_11 0 n6 ns11 0 5.90665563413e-07
Gc3_12 0 n6 ns12 0 -0.000198443946721
Gc3_13 0 n6 ns13 0 0.00192304825473
Gc3_14 0 n6 ns14 0 -0.000566304016694
Gc3_15 0 n6 ns15 0 0.000122567605318
Gc3_16 0 n6 ns16 0 0.00202026080356
Gc3_17 0 n6 ns17 0 -0.00102483192939
Gc3_18 0 n6 ns18 0 -0.000854051803251
Gc3_19 0 n6 ns19 0 0.00245268346892
Gc3_20 0 n6 ns20 0 3.05914239039e-05
Gc3_21 0 n6 ns21 0 0.000962184330504
Gc3_22 0 n6 ns22 0 -0.00297097635229
Gc3_23 0 n6 ns23 0 0.000379371110125
Gc3_24 0 n6 ns24 0 -0.000283240441489
Gc3_25 0 n6 ns25 0 -0.0013068023824
Gc3_26 0 n6 ns26 0 0.000546654703808
Gc3_27 0 n6 ns27 0 -0.000297402699456
Gc3_28 0 n6 ns28 0 0.00461950739998
Gc3_29 0 n6 ns29 0 -0.000143951324732
Gc3_30 0 n6 ns30 0 -6.79589454714e-06
Gc3_31 0 n6 ns31 0 0.00211122911201
Gc3_32 0 n6 ns32 0 0.000735630667363
Gc3_33 0 n6 ns33 0 -0.00159120797823
Gc3_34 0 n6 ns34 0 -7.68858091696e-08
Gc3_35 0 n6 ns35 0 7.62916969159e-08
Gc3_36 0 n6 ns36 0 0.00365912822664
Gc3_37 0 n6 ns37 0 -0.00129730774789
Gc3_38 0 n6 ns38 0 0.00410036975743
Gc3_39 0 n6 ns39 0 -9.4989846613e-05
Gc3_40 0 n6 ns40 0 7.84699803462e-05
Gc3_41 0 n6 ns41 0 3.67782252336e-05
Gc3_42 0 n6 ns42 0 0.00120082230502
Gc3_43 0 n6 ns43 0 -0.000672266393221
Gc3_44 0 n6 ns44 0 0.0110071498998
Gc3_45 0 n6 ns45 0 -0.000626987863511
Gc3_46 0 n6 ns46 0 -0.000362671536485
Gc3_47 0 n6 ns47 0 2.95357621462e-05
Gc3_48 0 n6 ns48 0 6.1400156188e-05
Gc3_49 0 n6 ns49 0 -2.78461209382e-05
Gc3_50 0 n6 ns50 0 -0.000569945753631
Gc3_51 0 n6 ns51 0 0.000392325648786
Gc3_52 0 n6 ns52 0 -6.35586166326e-05
Gc3_53 0 n6 ns53 0 -0.000915872558288
Gc3_54 0 n6 ns54 0 0.000807216140168
Gc3_55 0 n6 ns55 0 -0.000644933724948
Gc3_56 0 n6 ns56 0 0.000165210663446
Gc3_57 0 n6 ns57 0 0.0011205772275
Gc3_58 0 n6 ns58 0 -0.000412953991384
Gc3_59 0 n6 ns59 0 -0.00168227482435
Gc3_60 0 n6 ns60 0 0.00227949139312
Gc3_61 0 n6 ns61 0 2.88193669907e-05
Gc3_62 0 n6 ns62 0 0.00114430998004
Gc3_63 0 n6 ns63 0 -0.0018324964529
Gc3_64 0 n6 ns64 0 -0.000491925367295
Gc3_65 0 n6 ns65 0 -0.000411746476074
Gc3_66 0 n6 ns66 0 -0.00151364334553
Gc3_67 0 n6 ns67 0 0.00129229854957
Gc3_68 0 n6 ns68 0 -0.000307728432502
Gc3_69 0 n6 ns69 0 0.00253455728721
Gc3_70 0 n6 ns70 0 0.000985415806304
Gc3_71 0 n6 ns71 0 0.000272855979731
Gc3_72 0 n6 ns72 0 0.00237761973422
Gc3_73 0 n6 ns73 0 -0.00092858408069
Gc3_74 0 n6 ns74 0 -0.00197826374154
Gc3_75 0 n6 ns75 0 -4.98398079008e-08
Gc3_76 0 n6 ns76 0 9.01777729925e-08
Gc3_77 0 n6 ns77 0 0.00329828873602
Gc3_78 0 n6 ns78 0 -0.000880741887456
Gc3_79 0 n6 ns79 0 0.00500374270282
Gc3_80 0 n6 ns80 0 -0.000132046668672
Gc3_81 0 n6 ns81 0 0.000121810446273
Gc3_82 0 n6 ns82 0 4.20282906928e-05
Gc3_83 0 n6 ns83 0 0.000622817735617
Gc3_84 0 n6 ns84 0 0.0003468216456
Gc3_85 0 n6 ns85 0 0.0158488179785
Gc3_86 0 n6 ns86 0 -2.44855724501e-05
Gc3_87 0 n6 ns87 0 0.000118398319894
Gc3_88 0 n6 ns88 0 9.47577534054e-06
Gc3_89 0 n6 ns89 0 4.1017580839e-05
Gc3_90 0 n6 ns90 0 0.000374980821869
Gc3_91 0 n6 ns91 0 -0.000689497583554
Gc3_92 0 n6 ns92 0 -0.000408323102014
Gc3_93 0 n6 ns93 0 -0.000237482062545
Gc3_94 0 n6 ns94 0 -0.000667506981058
Gc3_95 0 n6 ns95 0 -0.00166187550201
Gc3_96 0 n6 ns96 0 -0.000489128435243
Gc3_97 0 n6 ns97 0 0.000191258663054
Gc3_98 0 n6 ns98 0 -0.00219755110943
Gc3_99 0 n6 ns99 0 0.000672397559947
Gc3_100 0 n6 ns100 0 0.00106521144016
Gc3_101 0 n6 ns101 0 -0.000671745141801
Gc3_102 0 n6 ns102 0 5.40910199782e-05
Gc3_103 0 n6 ns103 0 0.0009042352241
Gc3_104 0 n6 ns104 0 0.00285289890823
Gc3_105 0 n6 ns105 0 -0.000462717627875
Gc3_106 0 n6 ns106 0 -0.0002204861447
Gc3_107 0 n6 ns107 0 -0.00134114743243
Gc3_108 0 n6 ns108 0 -0.000708107958391
Gc3_109 0 n6 ns109 0 2.17764798373e-05
Gc3_110 0 n6 ns110 0 -0.0042419988757
Gc3_111 0 n6 ns111 0 0.00194466476079
Gc3_112 0 n6 ns112 0 0.000148294628119
Gc3_113 0 n6 ns113 0 0.00198268924683
Gc3_114 0 n6 ns114 0 0.00175094399968
Gc3_115 0 n6 ns115 0 0.00014080635265
Gc3_116 0 n6 ns116 0 2.20474511245e-08
Gc3_117 0 n6 ns117 0 -5.19212601961e-08
Gc3_118 0 n6 ns118 0 -0.00350008019516
Gc3_119 0 n6 ns119 0 -0.00218540943601
Gc3_120 0 n6 ns120 0 0.00841337577432
Gc3_121 0 n6 ns121 0 6.25986908191e-05
Gc3_122 0 n6 ns122 0 -3.57403029589e-05
Gc3_123 0 n6 ns123 0 -4.94792040011e-05
Gc3_124 0 n6 ns124 0 0.000511082015971
Gc3_125 0 n6 ns125 0 2.60459097861e-05
Gc3_126 0 n6 ns126 0 0.0154176536458
Gc3_127 0 n6 ns127 0 -0.000237142070687
Gc3_128 0 n6 ns128 0 -0.000127244073575
Gc3_129 0 n6 ns129 0 8.04553741206e-06
Gc3_130 0 n6 ns130 0 5.95608255486e-05
Gc3_131 0 n6 ns131 0 0.000328310481782
Gc3_132 0 n6 ns132 0 -0.000671536569042
Gc3_133 0 n6 ns133 0 -0.000183673957917
Gc3_134 0 n6 ns134 0 -0.000223355863493
Gc3_135 0 n6 ns135 0 -0.000621030392938
Gc3_136 0 n6 ns136 0 -0.00111728177183
Gc3_137 0 n6 ns137 0 -0.000622051044025
Gc3_138 0 n6 ns138 0 0.000223059722193
Gc3_139 0 n6 ns139 0 -0.00149122800645
Gc3_140 0 n6 ns140 0 0.000204450854434
Gc3_141 0 n6 ns141 0 0.000550974485488
Gc3_142 0 n6 ns142 0 6.81934240681e-05
Gc3_143 0 n6 ns143 0 5.81525661737e-05
Gc3_144 0 n6 ns144 0 0.00106943623812
Gc3_145 0 n6 ns145 0 0.00205841930736
Gc3_146 0 n6 ns146 0 -0.000170089033529
Gc3_147 0 n6 ns147 0 -0.000279273303972
Gc3_148 0 n6 ns148 0 -0.00155574321076
Gc3_149 0 n6 ns149 0 -0.000384752781555
Gc3_150 0 n6 ns150 0 -0.000213859186646
Gc3_151 0 n6 ns151 0 -0.00344242563413
Gc3_152 0 n6 ns152 0 0.00197289484747
Gc3_153 0 n6 ns153 0 0.000199981301808
Gc3_154 0 n6 ns154 0 0.00221860017269
Gc3_155 0 n6 ns155 0 0.00154522545739
Gc3_156 0 n6 ns156 0 0.000191373689857
Gc3_157 0 n6 ns157 0 -7.60082417947e-09
Gc3_158 0 n6 ns158 0 -2.8317933034e-08
Gc3_159 0 n6 ns159 0 -0.00294465955075
Gc3_160 0 n6 ns160 0 -0.00125670979908
Gc3_161 0 n6 ns161 0 0.00815166706371
Gc3_162 0 n6 ns162 0 2.4472731751e-05
Gc3_163 0 n6 ns163 0 -1.33930383202e-05
Gc3_164 0 n6 ns164 0 -2.80996781838e-05
Gc3_165 0 n6 ns165 0 -0.000166911214883
Gc3_166 0 n6 ns166 0 0.00225027123592
Gc3_167 0 n6 ns167 0 0.00250030242183
Gc3_168 0 n6 ns168 0 0.000256415841454
Gc3_169 0 n6 ns169 0 0.00060152904526
Gc3_170 0 n6 ns170 0 2.89959390936e-05
Gc3_171 0 n6 ns171 0 -9.2244006195e-06
Gc3_172 0 n6 ns172 0 0.000232965964427
Gc3_173 0 n6 ns173 0 -0.000148354462413
Gc3_174 0 n6 ns174 0 -0.000528095958861
Gc3_175 0 n6 ns175 0 -0.000188575028961
Gc3_176 0 n6 ns176 0 -0.00118814310715
Gc3_177 0 n6 ns177 0 -0.000644111809492
Gc3_178 0 n6 ns178 0 0.000693059711843
Gc3_179 0 n6 ns179 0 -0.000122240762253
Gc3_180 0 n6 ns180 0 0.00205913252809
Gc3_181 0 n6 ns181 0 -0.00131126797217
Gc3_182 0 n6 ns182 0 -0.00201614522466
Gc3_183 0 n6 ns183 0 -0.000318179135137
Gc3_184 0 n6 ns184 0 -8.27978616732e-06
Gc3_185 0 n6 ns185 0 0.000934960336034
Gc3_186 0 n6 ns186 0 0.00342219497571
Gc3_187 0 n6 ns187 0 -0.000806628823761
Gc3_188 0 n6 ns188 0 0.000130118722552
Gc3_189 0 n6 ns189 0 0.00131531596526
Gc3_190 0 n6 ns190 0 0.000804840787961
Gc3_191 0 n6 ns191 0 -0.00123634527382
Gc3_192 0 n6 ns192 0 0.00395908494121
Gc3_193 0 n6 ns193 0 0.000337360464878
Gc3_194 0 n6 ns194 0 0.000181403236162
Gc3_195 0 n6 ns195 0 0.00202826099998
Gc3_196 0 n6 ns196 0 0.000301276756349
Gc3_197 0 n6 ns197 0 -0.00132018080944
Gc3_198 0 n6 ns198 0 -4.34154655263e-08
Gc3_199 0 n6 ns199 0 5.71722116413e-08
Gc3_200 0 n6 ns200 0 -0.00321444862015
Gc3_201 0 n6 ns201 0 -0.00240503882459
Gc3_202 0 n6 ns202 0 -0.00151195989564
Gc3_203 0 n6 ns203 0 7.29354649917e-05
Gc3_204 0 n6 ns204 0 -3.63395790626e-05
Gc3_205 0 n6 ns205 0 -5.02559666484e-05
Gc3_206 0 n6 ns206 0 0.000120947908232
Gc3_207 0 n6 ns207 0 0.00141984460315
Gc3_208 0 n6 ns208 0 0.00306340774199
Gc3_209 0 n6 ns209 0 -3.7466019997e-05
Gc3_210 0 n6 ns210 0 0.000623229458563
Gc3_211 0 n6 ns211 0 5.8627222283e-05
Gc3_212 0 n6 ns212 0 -3.69500701307e-06
Gc3_213 0 n6 ns213 0 -0.000275308546505
Gc3_214 0 n6 ns214 0 -0.000256422507209
Gc3_215 0 n6 ns215 0 -0.000252661653207
Gc3_216 0 n6 ns216 0 -0.000298500819321
Gc3_217 0 n6 ns217 0 -0.00142977631652
Gc3_218 0 n6 ns218 0 -0.00120053308458
Gc3_219 0 n6 ns219 0 0.000777804548677
Gc3_220 0 n6 ns220 0 -0.000138856383605
Gc3_221 0 n6 ns221 0 0.0014114589645
Gc3_222 0 n6 ns222 0 -0.000596383799071
Gc3_223 0 n6 ns223 0 -0.000671282342161
Gc3_224 0 n6 ns224 0 0.00211242279142
Gc3_225 0 n6 ns225 0 1.57095753183e-05
Gc3_226 0 n6 ns226 0 0.001094374595
Gc3_227 0 n6 ns227 0 0.00260594385261
Gc3_228 0 n6 ns228 0 -0.000329667617836
Gc3_229 0 n6 ns229 0 0.000206153632373
Gc3_230 0 n6 ns230 0 0.00151603635954
Gc3_231 0 n6 ns231 0 0.000280119206176
Gc3_232 0 n6 ns232 0 -0.000338882994192
Gc3_233 0 n6 ns233 0 0.00378606988822
Gc3_234 0 n6 ns234 0 0.00190296322795
Gc3_235 0 n6 ns235 0 7.97932515163e-05
Gc3_236 0 n6 ns236 0 0.00211858745635
Gc3_237 0 n6 ns237 0 5.95420089525e-05
Gc3_238 0 n6 ns238 0 0.000695606581182
Gc3_239 0 n6 ns239 0 -2.44799803092e-08
Gc3_240 0 n6 ns240 0 6.75831068819e-08
Gc3_241 0 n6 ns241 0 -0.00338132161987
Gc3_242 0 n6 ns242 0 -0.00300610485832
Gc3_243 0 n6 ns243 0 -0.00266091339139
Gc3_244 0 n6 ns244 0 5.70513583392e-05
Gc3_245 0 n6 ns245 0 -2.16848054505e-05
Gc3_246 0 n6 ns246 0 -4.86544341792e-05
Gc3_247 0 n6 ns247 0 -0.000324421345584
Gc3_248 0 n6 ns248 0 0.00118334922662
Gc3_249 0 n6 ns249 0 0.00190977832385
Gc3_250 0 n6 ns250 0 0.000244622141111
Gc3_251 0 n6 ns251 0 -0.000413546465871
Gc3_252 0 n6 ns252 0 -2.02530707159e-05
Gc3_253 0 n6 ns253 0 2.56816640646e-05
Gc3_254 0 n6 ns254 0 0.000651798389401
Gc3_255 0 n6 ns255 0 -0.000703716342385
Gc3_256 0 n6 ns256 0 0.000456184164532
Gc3_257 0 n6 ns257 0 0.000152555134514
Gc3_258 0 n6 ns258 0 3.75099657009e-05
Gc3_259 0 n6 ns259 0 0.00368185821401
Gc3_260 0 n6 ns260 0 0.00059175849675
Gc3_261 0 n6 ns261 0 -0.000233364403769
Gc3_262 0 n6 ns262 0 -0.00205880142326
Gc3_263 0 n6 ns263 0 0.000174107857919
Gc3_264 0 n6 ns264 0 -0.00101899083634
Gc3_265 0 n6 ns265 0 -0.00872636889815
Gc3_266 0 n6 ns266 0 6.3251597381e-05
Gc3_267 0 n6 ns267 0 0.000812915088537
Gc3_268 0 n6 ns268 0 -0.00362540454348
Gc3_269 0 n6 ns269 0 -0.000244979296195
Gc3_270 0 n6 ns270 0 0.000108412629674
Gc3_271 0 n6 ns271 0 0.00148314227644
Gc3_272 0 n6 ns272 0 0.0022740458339
Gc3_273 0 n6 ns273 0 -0.00321242299281
Gc3_274 0 n6 ns274 0 -0.00945958934294
Gc3_275 0 n6 ns275 0 -0.00345308323979
Gc3_276 0 n6 ns276 0 0.000439393336655
Gc3_277 0 n6 ns277 0 0.00323065176491
Gc3_278 0 n6 ns278 0 0.00444676262754
Gc3_279 0 n6 ns279 0 -0.0100174333764
Gc3_280 0 n6 ns280 0 -2.1527097657e-07
Gc3_281 0 n6 ns281 0 3.66329864831e-08
Gc3_282 0 n6 ns282 0 0.00839809988958
Gc3_283 0 n6 ns283 0 0.0065421557599
Gc3_284 0 n6 ns284 0 -0.0112924053477
Gc3_285 0 n6 ns285 0 -0.00016918962574
Gc3_286 0 n6 ns286 0 0.000173093220371
Gc3_287 0 n6 ns287 0 7.85690361575e-05
Gc3_288 0 n6 ns288 0 0.000121286389634
Gc3_289 0 n6 ns289 0 -0.000325115877883
Gc3_290 0 n6 ns290 0 0.00361022284011
Gc3_291 0 n6 ns291 0 -0.000709323501645
Gc3_292 0 n6 ns292 0 -0.000121090531618
Gc3_293 0 n6 ns293 0 8.30519877633e-05
Gc3_294 0 n6 ns294 0 5.67515504533e-05
Gc3_295 0 n6 ns295 0 -0.000742883331771
Gc3_296 0 n6 ns296 0 -0.00133880476727
Gc3_297 0 n6 ns297 0 0.000734752677986
Gc3_298 0 n6 ns298 0 -0.000138596841884
Gc3_299 0 n6 ns299 0 -0.000368478496099
Gc3_300 0 n6 ns300 0 -0.0023773987931
Gc3_301 0 n6 ns301 0 0.000663508639462
Gc3_302 0 n6 ns302 0 -0.00011868787921
Gc3_303 0 n6 ns303 0 -0.00170537641497
Gc3_304 0 n6 ns304 0 0.000645644564635
Gc3_305 0 n6 ns305 0 -0.000828198405349
Gc3_306 0 n6 ns306 0 0.00900347840113
Gc3_307 0 n6 ns307 0 2.57016177928e-05
Gc3_308 0 n6 ns308 0 0.00111487059029
Gc3_309 0 n6 ns309 0 -0.00120183342464
Gc3_310 0 n6 ns310 0 0.000897357900502
Gc3_311 0 n6 ns311 0 0.00031871032977
Gc3_312 0 n6 ns312 0 0.0014265794771
Gc3_313 0 n6 ns313 0 -0.00180708105219
Gc3_314 0 n6 ns314 0 0.00201465869044
Gc3_315 0 n6 ns315 0 -5.06146266076e-06
Gc3_316 0 n6 ns316 0 0.0060181753606
Gc3_317 0 n6 ns317 0 -5.39835575948e-06
Gc3_318 0 n6 ns318 0 0.00149220853054
Gc3_319 0 n6 ns319 0 -0.00201818474574
Gc3_320 0 n6 ns320 0 0.00593758634222
Gc3_321 0 n6 ns321 0 7.218324861e-08
Gc3_322 0 n6 ns322 0 5.68519697512e-08
Gc3_323 0 n6 ns323 0 -0.0017212310191
Gc3_324 0 n6 ns324 0 -0.0055984844277
Gc3_325 0 n6 ns325 0 -0.00387867832314
Gc3_326 0 n6 ns326 0 1.34895797602e-05
Gc3_327 0 n6 ns327 0 -5.70992274257e-06
Gc3_328 0 n6 ns328 0 -2.20135889178e-05
Gd3_1 0 n6 ni1 0 -0.000972172366039
Gd3_2 0 n6 ni2 0 -0.00323133395277
Gd3_3 0 n6 ni3 0 -0.00188647581823
Gd3_4 0 n6 ni4 0 -0.00200310973668
Gd3_5 0 n6 ni5 0 0.000741517560298
Gd3_6 0 n6 ni6 0 0.000154238122533
Gd3_7 0 n6 ni7 0 8.57652214489e-05
Gd3_8 0 n6 ni8 0 -0.000653022950265
Gc4_1 0 n8 ns1 0 0.00118894875336
Gc4_2 0 n8 ns2 0 -0.000676916225506
Gc4_3 0 n8 ns3 0 0.0110574899173
Gc4_4 0 n8 ns4 0 -0.000623359640061
Gc4_5 0 n8 ns5 0 -0.000348849150533
Gc4_6 0 n8 ns6 0 3.20295767788e-05
Gc4_7 0 n8 ns7 0 6.15035459855e-05
Gc4_8 0 n8 ns8 0 -2.12540022456e-05
Gc4_9 0 n8 ns9 0 -0.000581980021629
Gc4_10 0 n8 ns10 0 0.000403702531675
Gc4_11 0 n8 ns11 0 -6.63844884574e-05
Gc4_12 0 n8 ns12 0 -0.000944838708054
Gc4_13 0 n8 ns13 0 0.000784345111546
Gc4_14 0 n8 ns14 0 -0.000645758961471
Gc4_15 0 n8 ns15 0 0.000170130816148
Gc4_16 0 n8 ns16 0 0.00111523912749
Gc4_17 0 n8 ns17 0 -0.000433299131502
Gc4_18 0 n8 ns18 0 -0.00171856094666
Gc4_19 0 n8 ns19 0 0.0023126606395
Gc4_20 0 n8 ns20 0 3.09075555915e-05
Gc4_21 0 n8 ns21 0 0.00115021921206
Gc4_22 0 n8 ns22 0 -0.0018217581713
Gc4_23 0 n8 ns23 0 -0.000478204078206
Gc4_24 0 n8 ns24 0 -0.000420842606176
Gc4_25 0 n8 ns25 0 -0.00152062114668
Gc4_26 0 n8 ns26 0 0.00131425885931
Gc4_27 0 n8 ns27 0 -0.000326310958976
Gc4_28 0 n8 ns28 0 0.00250079986925
Gc4_29 0 n8 ns29 0 0.000981501144642
Gc4_30 0 n8 ns30 0 0.000284041655392
Gc4_31 0 n8 ns31 0 0.00237887192993
Gc4_32 0 n8 ns32 0 -0.000964477057254
Gc4_33 0 n8 ns33 0 -0.0019911732533
Gc4_34 0 n8 ns34 0 -4.9742062343e-08
Gc4_35 0 n8 ns35 0 9.21955919436e-08
Gc4_36 0 n8 ns36 0 0.00327616540576
Gc4_37 0 n8 ns37 0 -0.000893712046492
Gc4_38 0 n8 ns38 0 0.00500601617183
Gc4_39 0 n8 ns39 0 -0.000132083012945
Gc4_40 0 n8 ns40 0 0.000119312133871
Gc4_41 0 n8 ns41 0 4.21153651426e-05
Gc4_42 0 n8 ns42 0 0.000671636723896
Gc4_43 0 n8 ns43 0 -0.000321839657415
Gc4_44 0 n8 ns44 0 0.00971084028064
Gc4_45 0 n8 ns45 0 -0.000355405282424
Gc4_46 0 n8 ns46 0 -7.35659824784e-05
Gc4_47 0 n8 ns47 0 2.4902639054e-05
Gc4_48 0 n8 ns48 0 3.88222338226e-05
Gc4_49 0 n8 ns49 0 -0.000189732774032
Gc4_50 0 n8 ns50 0 -0.000800844730628
Gc4_51 0 n8 ns51 0 0.000274833514475
Gc4_52 0 n8 ns52 0 -8.40250391195e-05
Gc4_53 0 n8 ns53 0 -0.00076589180168
Gc4_54 0 n8 ns54 0 0.00092214517528
Gc4_55 0 n8 ns55 0 -0.00076242456108
Gc4_56 0 n8 ns56 0 0.000223423045858
Gc4_57 0 n8 ns57 0 0.000804226253476
Gc4_58 0 n8 ns58 0 -0.000385443122614
Gc4_59 0 n8 ns59 0 -0.000209770560508
Gc4_60 0 n8 ns60 0 0.0021559162336
Gc4_61 0 n8 ns61 0 4.16486543878e-05
Gc4_62 0 n8 ns62 0 0.00129074572556
Gc4_63 0 n8 ns63 0 -0.00140746164123
Gc4_64 0 n8 ns64 0 -0.000128905797931
Gc4_65 0 n8 ns65 0 -0.00031978204782
Gc4_66 0 n8 ns66 0 -0.00174618237964
Gc4_67 0 n8 ns67 0 4.58637463423e-05
Gc4_68 0 n8 ns68 0 -0.00056907043738
Gc4_69 0 n8 ns69 0 0.0021878803474
Gc4_70 0 n8 ns70 0 0.00153777590791
Gc4_71 0 n8 ns71 0 8.59639878114e-05
Gc4_72 0 n8 ns72 0 0.00257924049568
Gc4_73 0 n8 ns73 0 0.00137403886359
Gc4_74 0 n8 ns74 0 -0.000114557071977
Gc4_75 0 n8 ns75 0 -6.49722977285e-09
Gc4_76 0 n8 ns76 0 2.97776901125e-08
Gc4_77 0 n8 ns77 0 0.00149377882793
Gc4_78 0 n8 ns78 0 -0.000183127913555
Gc4_79 0 n8 ns79 0 0.0061215129511
Gc4_80 0 n8 ns80 0 -4.33872055252e-05
Gc4_81 0 n8 ns81 0 2.47058011547e-05
Gc4_82 0 n8 ns82 0 1.88757541422e-05
Gc4_83 0 n8 ns83 0 0.00051108201962
Gc4_84 0 n8 ns84 0 2.60459130035e-05
Gc4_85 0 n8 ns85 0 0.0154176536344
Gc4_86 0 n8 ns86 0 -0.00023714207219
Gc4_87 0 n8 ns87 0 -0.000127244078721
Gc4_88 0 n8 ns88 0 8.04553588717e-06
Gc4_89 0 n8 ns89 0 5.95608260927e-05
Gc4_90 0 n8 ns90 0 0.000328310476862
Gc4_91 0 n8 ns91 0 -0.000671536563405
Gc4_92 0 n8 ns92 0 -0.000183673961208
Gc4_93 0 n8 ns93 0 -0.000223355862077
Gc4_94 0 n8 ns94 0 -0.000621030379873
Gc4_95 0 n8 ns95 0 -0.00111728176191
Gc4_96 0 n8 ns96 0 -0.000622051045026
Gc4_97 0 n8 ns97 0 0.000223059721304
Gc4_98 0 n8 ns98 0 -0.00149122800518
Gc4_99 0 n8 ns99 0 0.000204450858807
Gc4_100 0 n8 ns100 0 0.000550974507121
Gc4_101 0 n8 ns101 0 6.81934141471e-05
Gc4_102 0 n8 ns102 0 5.81525670574e-05
Gc4_103 0 n8 ns103 0 0.00106943623805
Gc4_104 0 n8 ns104 0 0.00205841930057
Gc4_105 0 n8 ns105 0 -0.000170089032753
Gc4_106 0 n8 ns106 0 -0.000279273301923
Gc4_107 0 n8 ns107 0 -0.00155574321013
Gc4_108 0 n8 ns108 0 -0.000384752789298
Gc4_109 0 n8 ns109 0 -0.000213859177204
Gc4_110 0 n8 ns110 0 -0.00344242562444
Gc4_111 0 n8 ns111 0 0.00197289483767
Gc4_112 0 n8 ns112 0 0.000199981301322
Gc4_113 0 n8 ns113 0 0.00221860017365
Gc4_114 0 n8 ns114 0 0.00154522546965
Gc4_115 0 n8 ns115 0 0.000191373688541
Gc4_116 0 n8 ns116 0 -7.60082504571e-09
Gc4_117 0 n8 ns117 0 -2.83179341953e-08
Gc4_118 0 n8 ns118 0 -0.0029446595374
Gc4_119 0 n8 ns119 0 -0.00125670981526
Gc4_120 0 n8 ns120 0 0.00815166708067
Gc4_121 0 n8 ns121 0 2.44727295537e-05
Gc4_122 0 n8 ns122 0 -1.33930364482e-05
Gc4_123 0 n8 ns123 0 -2.80996788747e-05
Gc4_124 0 n8 ns124 0 -0.000237064260087
Gc4_125 0 n8 ns125 0 0.000350254198921
Gc4_126 0 n8 ns126 0 0.0110781016021
Gc4_127 0 n8 ns127 0 0.000126341252738
Gc4_128 0 n8 ns128 0 0.000190168338928
Gc4_129 0 n8 ns129 0 3.4378312689e-05
Gc4_130 0 n8 ns130 0 3.16607997719e-05
Gc4_131 0 n8 ns131 0 0.000206248018892
Gc4_132 0 n8 ns132 0 -0.0007506090833
Gc4_133 0 n8 ns133 0 -2.55426996219e-05
Gc4_134 0 n8 ns134 0 -0.000174569440609
Gc4_135 0 n8 ns135 0 -0.00038640091249
Gc4_136 0 n8 ns136 0 -0.00112786182533
Gc4_137 0 n8 ns137 0 -0.000786326350457
Gc4_138 0 n8 ns138 0 0.000278865031166
Gc4_139 0 n8 ns139 0 -0.000989072725531
Gc4_140 0 n8 ns140 0 1.86470843787e-07
Gc4_141 0 n8 ns141 0 0.000137484460128
Gc4_142 0 n8 ns142 0 -0.000261321217063
Gc4_143 0 n8 ns143 0 7.73096192588e-05
Gc4_144 0 n8 ns144 0 0.00125577830353
Gc4_145 0 n8 ns145 0 0.00134209183419
Gc4_146 0 n8 ns146 0 -0.000105536174415
Gc4_147 0 n8 ns147 0 -0.000273836698421
Gc4_148 0 n8 ns148 0 -0.00179835980268
Gc4_149 0 n8 ns149 0 9.09278274939e-06
Gc4_150 0 n8 ns150 0 0.000274265593197
Gc4_151 0 n8 ns151 0 -0.0024433185897
Gc4_152 0 n8 ns152 0 0.00126975687625
Gc4_153 0 n8 ns153 0 0.000215931856957
Gc4_154 0 n8 ns154 0 0.00289779124509
Gc4_155 0 n8 ns155 0 0.000826884299992
Gc4_156 0 n8 ns156 0 -0.000941043994351
Gc4_157 0 n8 ns157 0 -4.39987538376e-08
Gc4_158 0 n8 ns158 0 -1.10425852739e-07
Gc4_159 0 n8 ns159 0 -0.00151456198407
Gc4_160 0 n8 ns160 0 -0.00144865658362
Gc4_161 0 n8 ns161 0 0.00884096954382
Gc4_162 0 n8 ns162 0 7.83661883618e-05
Gc4_163 0 n8 ns163 0 -5.52325332421e-05
Gc4_164 0 n8 ns164 0 -4.50717681383e-05
Gc4_165 0 n8 ns165 0 0.000129073015595
Gc4_166 0 n8 ns166 0 0.00141645523799
Gc4_167 0 n8 ns167 0 0.00311287289376
Gc4_168 0 n8 ns168 0 -4.31502771731e-05
Gc4_169 0 n8 ns169 0 0.000612159456529
Gc4_170 0 n8 ns170 0 5.82262908211e-05
Gc4_171 0 n8 ns171 0 -3.08914199957e-06
Gc4_172 0 n8 ns172 0 -0.000274645592877
Gc4_173 0 n8 ns173 0 -0.000252570747624
Gc4_174 0 n8 ns174 0 -0.000256460727935
Gc4_175 0 n8 ns175 0 -0.000296177061116
Gc4_176 0 n8 ns176 0 -0.00143137239016
Gc4_177 0 n8 ns177 0 -0.00119809218779
Gc4_178 0 n8 ns178 0 0.000780778861204
Gc4_179 0 n8 ns179 0 -0.000142207368358
Gc4_180 0 n8 ns180 0 0.00141018840976
Gc4_181 0 n8 ns181 0 -0.000604097708004
Gc4_182 0 n8 ns182 0 -0.00065962835929
Gc4_183 0 n8 ns183 0 0.00212798981143
Gc4_184 0 n8 ns184 0 1.97884506441e-05
Gc4_185 0 n8 ns185 0 0.00109829084526
Gc4_186 0 n8 ns186 0 0.00259709324368
Gc4_187 0 n8 ns187 0 -0.000337979899406
Gc4_188 0 n8 ns188 0 0.000214554901651
Gc4_189 0 n8 ns189 0 0.00151751533948
Gc4_190 0 n8 ns190 0 0.000282669904488
Gc4_191 0 n8 ns191 0 -0.000324800322872
Gc4_192 0 n8 ns192 0 0.0037609198556
Gc4_193 0 n8 ns193 0 0.00188531006715
Gc4_194 0 n8 ns194 0 9.43167389621e-05
Gc4_195 0 n8 ns195 0 0.00211967729628
Gc4_196 0 n8 ns196 0 3.21302792469e-05
Gc4_197 0 n8 ns197 0 0.00070143995301
Gc4_198 0 n8 ns198 0 -2.31218367432e-08
Gc4_199 0 n8 ns199 0 6.84433267611e-08
Gc4_200 0 n8 ns200 0 -0.00337687045367
Gc4_201 0 n8 ns201 0 -0.00299745088388
Gc4_202 0 n8 ns202 0 -0.00266329006808
Gc4_203 0 n8 ns203 0 5.42352492765e-05
Gc4_204 0 n8 ns204 0 -1.67210579632e-05
Gc4_205 0 n8 ns205 0 -4.71736483341e-05
Gc4_206 0 n8 ns206 0 -4.21264438093e-05
Gc4_207 0 n8 ns207 0 0.00124622579437
Gc4_208 0 n8 ns208 0 0.00407799813557
Gc4_209 0 n8 ns209 0 -0.000330812739226
Gc4_210 0 n8 ns210 0 0.000204660697092
Gc4_211 0 n8 ns211 0 7.23805190898e-05
Gc4_212 0 n8 ns212 0 4.68952237992e-05
Gc4_213 0 n8 ns213 0 -0.000204041345023
Gc4_214 0 n8 ns214 0 -0.00096696850206
Gc4_215 0 n8 ns215 0 3.55739968537e-05
Gc4_216 0 n8 ns216 0 -0.000281889469703
Gc4_217 0 n8 ns217 0 -0.000609212426409
Gc4_218 0 n8 ns218 0 -0.00128822937471
Gc4_219 0 n8 ns219 0 0.000890256315592
Gc4_220 0 n8 ns220 0 -0.000198484767072
Gc4_221 0 n8 ns221 0 0.000752281993855
Gc4_222 0 n8 ns222 0 -0.000380875326234
Gc4_223 0 n8 ns223 0 -0.00268074064684
Gc4_224 0 n8 ns224 0 0.00359390730253
Gc4_225 0 n8 ns225 0 -1.59467413408e-05
Gc4_226 0 n8 ns226 0 0.00126913012178
Gc4_227 0 n8 ns227 0 0.00211979390304
Gc4_228 0 n8 ns228 0 2.25911526739e-05
Gc4_229 0 n8 ns229 0 0.000204548170491
Gc4_230 0 n8 ns230 0 0.0017466238491
Gc4_231 0 n8 ns231 0 -6.77781433899e-05
Gc4_232 0 n8 ns232 0 -0.000359136705642
Gc4_233 0 n8 ns233 0 0.00281104568729
Gc4_234 0 n8 ns234 0 0.00370777520941
Gc4_235 0 n8 ns235 0 0.000174675083884
Gc4_236 0 n8 ns236 0 0.00221810100898
Gc4_237 0 n8 ns237 0 -0.000902599595803
Gc4_238 0 n8 ns238 0 0.00207796718514
Gc4_239 0 n8 ns239 0 3.95983836933e-09
Gc4_240 0 n8 ns240 0 7.66605647956e-08
Gc4_241 0 n8 ns241 0 -0.00354740376227
Gc4_242 0 n8 ns242 0 -0.00360204025919
Gc4_243 0 n8 ns243 0 -0.00370562138916
Gc4_244 0 n8 ns244 0 3.4953113228e-05
Gc4_245 0 n8 ns245 0 -3.57372307259e-06
Gc4_246 0 n8 ns246 0 -4.06190464786e-05
Gc4_247 0 n8 ns247 0 0.000121344647971
Gc4_248 0 n8 ns248 0 -0.000325961883094
Gc4_249 0 n8 ns249 0 0.00359742452754
Gc4_250 0 n8 ns250 0 -0.000708945405536
Gc4_251 0 n8 ns251 0 -0.000121411780262
Gc4_252 0 n8 ns252 0 8.30292413242e-05
Gc4_253 0 n8 ns253 0 5.7527700873e-05
Gc4_254 0 n8 ns254 0 -0.000744476642642
Gc4_255 0 n8 ns255 0 -0.00133493948347
Gc4_256 0 n8 ns256 0 0.000733789844695
Gc4_257 0 n8 ns257 0 -0.000136224410206
Gc4_258 0 n8 ns258 0 -0.000359711963098
Gc4_259 0 n8 ns259 0 -0.00238177555209
Gc4_260 0 n8 ns260 0 0.00066286324093
Gc4_261 0 n8 ns261 0 -0.000117838014525
Gc4_262 0 n8 ns262 0 -0.00170325184119
Gc4_263 0 n8 ns263 0 0.000644986545017
Gc4_264 0 n8 ns264 0 -0.000831056432259
Gc4_265 0 n8 ns265 0 0.00899710467423
Gc4_266 0 n8 ns266 0 2.52737816005e-05
Gc4_267 0 n8 ns267 0 0.00111478812059
Gc4_268 0 n8 ns268 0 -0.0012014750705
Gc4_269 0 n8 ns269 0 0.000900661473116
Gc4_270 0 n8 ns270 0 0.000318546828952
Gc4_271 0 n8 ns271 0 0.00142539155153
Gc4_272 0 n8 ns272 0 -0.00180111683314
Gc4_273 0 n8 ns273 0 0.00201394484126
Gc4_274 0 n8 ns274 0 -1.71427684399e-05
Gc4_275 0 n8 ns275 0 0.00602797196564
Gc4_276 0 n8 ns276 0 -1.089463909e-06
Gc4_277 0 n8 ns277 0 0.00148641971301
Gc4_278 0 n8 ns278 0 -0.00202043687441
Gc4_279 0 n8 ns279 0 0.00595636332526
Gc4_280 0 n8 ns280 0 6.9470710593e-08
Gc4_281 0 n8 ns281 0 5.62805767609e-08
Gc4_282 0 n8 ns282 0 -0.00171154845479
Gc4_283 0 n8 ns283 0 -0.00560078744631
Gc4_284 0 n8 ns284 0 -0.00387361141985
Gc4_285 0 n8 ns285 0 1.36841921065e-05
Gc4_286 0 n8 ns286 0 -6.00776963707e-06
Gc4_287 0 n8 ns287 0 -2.2137672939e-05
Gc4_288 0 n8 ns288 0 -0.000123287899883
Gc4_289 0 n8 ns289 0 0.0019210620959
Gc4_290 0 n8 ns290 0 0.00386591022754
Gc4_291 0 n8 ns291 0 0.000360311092183
Gc4_292 0 n8 ns292 0 -4.65304053698e-05
Gc4_293 0 n8 ns293 0 -2.58240941102e-05
Gc4_294 0 n8 ns294 0 1.28825767756e-05
Gc4_295 0 n8 ns295 0 0.000655698641885
Gc4_296 0 n8 ns296 0 -0.000387507592315
Gc4_297 0 n8 ns297 0 -1.36628697013e-05
Gc4_298 0 n8 ns298 0 0.000114932822709
Gc4_299 0 n8 ns299 0 -0.000918842202226
Gc4_300 0 n8 ns300 0 0.00344125534057
Gc4_301 0 n8 ns301 0 0.000910740816851
Gc4_302 0 n8 ns302 0 -0.000299543808355
Gc4_303 0 n8 ns303 0 -0.000812183864768
Gc4_304 0 n8 ns304 0 -0.000740701344855
Gc4_305 0 n8 ns305 0 -0.000872641318431
Gc4_306 0 n8 ns306 0 -0.0092649315276
Gc4_307 0 n8 ns307 0 6.59383207613e-05
Gc4_308 0 n8 ns308 0 0.00117699904677
Gc4_309 0 n8 ns309 0 -0.00189103900896
Gc4_310 0 n8 ns310 0 -0.000902379595139
Gc4_311 0 n8 ns311 0 8.66707659028e-05
Gc4_312 0 n8 ns312 0 0.00191075054617
Gc4_313 0 n8 ns313 0 0.00304938504678
Gc4_314 0 n8 ns314 0 -0.00353907929387
Gc4_315 0 n8 ns315 0 -0.00791964760467
Gc4_316 0 n8 ns316 0 -0.00408517849945
Gc4_317 0 n8 ns317 0 0.000494819851532
Gc4_318 0 n8 ns318 0 0.00403344755383
Gc4_319 0 n8 ns319 0 0.00430921952558
Gc4_320 0 n8 ns320 0 -0.0106919373957
Gc4_321 0 n8 ns321 0 -1.9911159872e-07
Gc4_322 0 n8 ns322 0 -1.6662902663e-08
Gc4_323 0 n8 ns323 0 0.00677979779149
Gc4_324 0 n8 ns324 0 0.0056190282765
Gc4_325 0 n8 ns325 0 -0.0117036921473
Gc4_326 0 n8 ns326 0 -0.000179422020226
Gc4_327 0 n8 ns327 0 0.000188302150097
Gc4_328 0 n8 ns328 0 7.34036547335e-05
Gd4_1 0 n8 ni1 0 -0.00323933071966
Gd4_2 0 n8 ni2 0 -0.00201358223693
Gd4_3 0 n8 ni3 0 -0.00200310973628
Gd4_4 0 n8 ni4 0 -0.000508560646444
Gd4_5 0 n8 ni5 0 0.000139154660234
Gd4_6 0 n8 ni6 0 -6.21146550553e-05
Gd4_7 0 n8 ni7 0 -0.000649725279825
Gd4_8 0 n8 ni8 0 -0.000119260531111
Gc5_1 0 n10 ns1 0 -0.000322992496672
Gc5_2 0 n10 ns2 0 0.00121079940878
Gc5_3 0 n10 ns3 0 0.00203083271785
Gc5_4 0 n10 ns4 0 0.000239347633125
Gc5_5 0 n10 ns5 0 -0.000413648366014
Gc5_6 0 n10 ns6 0 -1.87116733949e-05
Gc5_7 0 n10 ns7 0 2.56660645929e-05
Gc5_8 0 n10 ns8 0 0.000658121946573
Gc5_9 0 n10 ns9 0 -0.000710309798553
Gc5_10 0 n10 ns10 0 0.000463646732997
Gc5_11 0 n10 ns11 0 0.000150389753211
Gc5_12 0 n10 ns12 0 2.28895441532e-05
Gc5_13 0 n10 ns13 0 0.00366254489251
Gc5_14 0 n10 ns14 0 0.000598822461651
Gc5_15 0 n10 ns15 0 -0.000235857081366
Gc5_16 0 n10 ns16 0 -0.00205496700118
Gc5_17 0 n10 ns17 0 0.000167887360801
Gc5_18 0 n10 ns18 0 -0.0010728323505
Gc5_19 0 n10 ns19 0 -0.00873147946016
Gc5_20 0 n10 ns20 0 6.78027940268e-05
Gc5_21 0 n10 ns21 0 0.00082086168373
Gc5_22 0 n10 ns22 0 -0.00360753947577
Gc5_23 0 n10 ns23 0 -0.000242586208815
Gc5_24 0 n10 ns24 0 0.000118807667818
Gc5_25 0 n10 ns25 0 0.00148780001631
Gc5_26 0 n10 ns26 0 0.00230778306253
Gc5_27 0 n10 ns27 0 -0.00322170866839
Gc5_28 0 n10 ns28 0 -0.00950201883598
Gc5_29 0 n10 ns29 0 -0.00349161427077
Gc5_30 0 n10 ns30 0 0.000466911467496
Gc5_31 0 n10 ns31 0 0.0032397627922
Gc5_32 0 n10 ns32 0 0.00440658192551
Gc5_33 0 n10 ns33 0 -0.0100823556489
Gc5_34 0 n10 ns34 0 -2.14070142928e-07
Gc5_35 0 n10 ns35 0 3.72242718744e-08
Gc5_36 0 n10 ns36 0 0.00839546284048
Gc5_37 0 n10 ns37 0 0.00649601247951
Gc5_38 0 n10 ns38 0 -0.0112442593352
Gc5_39 0 n10 ns39 0 -0.000171659471077
Gc5_40 0 n10 ns40 0 0.000176355968619
Gc5_41 0 n10 ns41 0 7.82761874601e-05
Gc5_42 0 n10 ns42 0 0.000132934056899
Gc5_43 0 n10 ns43 0 -0.000257149773705
Gc5_44 0 n10 ns44 0 0.00371549142994
Gc5_45 0 n10 ns45 0 -0.000719470011461
Gc5_46 0 n10 ns46 0 -0.000141524833495
Gc5_47 0 n10 ns47 0 8.0525444626e-05
Gc5_48 0 n10 ns48 0 5.75435505392e-05
Gc5_49 0 n10 ns49 0 -0.000748256712305
Gc5_50 0 n10 ns50 0 -0.00132691991943
Gc5_51 0 n10 ns51 0 0.000726677375263
Gc5_52 0 n10 ns52 0 -0.000135228052002
Gc5_53 0 n10 ns53 0 -0.000344217888005
Gc5_54 0 n10 ns54 0 -0.00236548128053
Gc5_55 0 n10 ns55 0 0.000665752921519
Gc5_56 0 n10 ns56 0 -0.000123573553258
Gc5_57 0 n10 ns57 0 -0.00169983824802
Gc5_58 0 n10 ns58 0 0.000644176094972
Gc5_59 0 n10 ns59 0 -0.000798459518905
Gc5_60 0 n10 ns60 0 0.00898286059012
Gc5_61 0 n10 ns61 0 3.17028766651e-05
Gc5_62 0 n10 ns62 0 0.00112134101667
Gc5_63 0 n10 ns63 0 -0.00121178421006
Gc5_64 0 n10 ns64 0 0.000906037631792
Gc5_65 0 n10 ns65 0 0.000331291489337
Gc5_66 0 n10 ns66 0 0.00142696441725
Gc5_67 0 n10 ns67 0 -0.00179699076009
Gc5_68 0 n10 ns68 0 0.00203917426644
Gc5_69 0 n10 ns69 0 -1.5653449424e-05
Gc5_70 0 n10 ns70 0 0.00596420704353
Gc5_71 0 n10 ns71 0 8.05463472641e-06
Gc5_72 0 n10 ns72 0 0.00150076010786
Gc5_73 0 n10 ns73 0 -0.00201222868688
Gc5_74 0 n10 ns74 0 0.00587963329254
Gc5_75 0 n10 ns75 0 6.97571882663e-08
Gc5_76 0 n10 ns76 0 5.65858505924e-08
Gc5_77 0 n10 ns77 0 -0.00169605229871
Gc5_78 0 n10 ns78 0 -0.00572082057741
Gc5_79 0 n10 ns79 0 -0.0037857592547
Gc5_80 0 n10 ns80 0 3.30569864166e-06
Gc5_81 0 n10 ns81 0 -6.96917937575e-07
Gc5_82 0 n10 ns82 0 -1.89231262395e-05
Gc5_83 0 n10 ns83 0 -0.000166911236891
Gc5_84 0 n10 ns84 0 0.00225027119503
Gc5_85 0 n10 ns85 0 0.00250030242202
Gc5_86 0 n10 ns86 0 0.000256415852394
Gc5_87 0 n10 ns87 0 0.000601529070809
Gc5_88 0 n10 ns88 0 2.89959433545e-05
Gc5_89 0 n10 ns89 0 -9.22440152811e-06
Gc5_90 0 n10 ns90 0 0.000232965975178
Gc5_91 0 n10 ns91 0 -0.000148354481965
Gc5_92 0 n10 ns92 0 -0.000528095950413
Gc5_93 0 n10 ns93 0 -0.000188575033731
Gc5_94 0 n10 ns94 0 -0.00118814313889
Gc5_95 0 n10 ns95 0 -0.000644111839448
Gc5_96 0 n10 ns96 0 0.000693059713603
Gc5_97 0 n10 ns97 0 -0.000122240760072
Gc5_98 0 n10 ns98 0 0.0020591325311
Gc5_99 0 n10 ns99 0 -0.00131126798484
Gc5_100 0 n10 ns100 0 -0.00201614530532
Gc5_101 0 n10 ns101 0 -0.000318179134666
Gc5_102 0 n10 ns102 0 -8.27978876727e-06
Gc5_103 0 n10 ns103 0 0.000934960334052
Gc5_104 0 n10 ns104 0 0.00342219499198
Gc5_105 0 n10 ns105 0 -0.000806628826484
Gc5_106 0 n10 ns106 0 0.000130118720712
Gc5_107 0 n10 ns107 0 0.00131531596721
Gc5_108 0 n10 ns108 0 0.000804840799257
Gc5_109 0 n10 ns109 0 -0.00123634525774
Gc5_110 0 n10 ns110 0 0.00395908496044
Gc5_111 0 n10 ns111 0 0.000337360351978
Gc5_112 0 n10 ns112 0 0.000181403223524
Gc5_113 0 n10 ns113 0 0.00202826105091
Gc5_114 0 n10 ns114 0 0.000301276750324
Gc5_115 0 n10 ns115 0 -0.00132018100296
Gc5_116 0 n10 ns116 0 -4.34154582132e-08
Gc5_117 0 n10 ns117 0 5.71722157563e-08
Gc5_118 0 n10 ns118 0 -0.0032144486359
Gc5_119 0 n10 ns119 0 -0.00240503913425
Gc5_120 0 n10 ns120 0 -0.00151195972703
Gc5_121 0 n10 ns121 0 7.29354904336e-05
Gc5_122 0 n10 ns122 0 -3.63395761703e-05
Gc5_123 0 n10 ns123 0 -5.02559708529e-05
Gc5_124 0 n10 ns124 0 0.0001290730301
Gc5_125 0 n10 ns125 0 0.00141645525246
Gc5_126 0 n10 ns126 0 0.00311287286429
Gc5_127 0 n10 ns127 0 -4.31502861043e-05
Gc5_128 0 n10 ns128 0 0.000612159437615
Gc5_129 0 n10 ns129 0 5.82262888965e-05
Gc5_130 0 n10 ns130 0 -3.08914243137e-06
Gc5_131 0 n10 ns131 0 -0.000274645597111
Gc5_132 0 n10 ns132 0 -0.000252570736705
Gc5_133 0 n10 ns133 0 -0.00025646073279
Gc5_134 0 n10 ns134 0 -0.000296177059388
Gc5_135 0 n10 ns135 0 -0.00143137237421
Gc5_136 0 n10 ns136 0 -0.00119809216591
Gc5_137 0 n10 ns137 0 0.000780778860495
Gc5_138 0 n10 ns138 0 -0.000142207369981
Gc5_139 0 n10 ns139 0 0.00141018840556
Gc5_140 0 n10 ns140 0 -0.000604097700641
Gc5_141 0 n10 ns141 0 -0.000659628303192
Gc5_142 0 n10 ns142 0 0.00212798983214
Gc5_143 0 n10 ns143 0 1.97884518077e-05
Gc5_144 0 n10 ns144 0 0.00109829084714
Gc5_145 0 n10 ns145 0 0.00259709323541
Gc5_146 0 n10 ns146 0 -0.000337979910965
Gc5_147 0 n10 ns147 0 0.000214554899917
Gc5_148 0 n10 ns148 0 0.00151751534304
Gc5_149 0 n10 ns149 0 0.000282669865261
Gc5_150 0 n10 ns150 0 -0.000324800349357
Gc5_151 0 n10 ns151 0 0.00376091989052
Gc5_152 0 n10 ns152 0 0.00188531016649
Gc5_153 0 n10 ns153 0 9.43167340372e-05
Gc5_154 0 n10 ns154 0 0.0021196772536
Gc5_155 0 n10 ns155 0 3.21303382088e-05
Gc5_156 0 n10 ns156 0 0.000701440103913
Gc5_157 0 n10 ns157 0 -2.31218407779e-08
Gc5_158 0 n10 ns158 0 6.84433218562e-08
Gc5_159 0 n10 ns159 0 -0.00337687043633
Gc5_160 0 n10 ns160 0 -0.00299745067638
Gc5_161 0 n10 ns161 0 -0.00266329018727
Gc5_162 0 n10 ns162 0 5.42352343729e-05
Gc5_163 0 n10 ns163 0 -1.67210572071e-05
Gc5_164 0 n10 ns164 0 -4.71736472521e-05
Gc5_165 0 n10 ns165 0 0.000593814951068
Gc5_166 0 n10 ns166 0 0.000380119232448
Gc5_167 0 n10 ns167 0 0.015815244683
Gc5_168 0 n10 ns168 0 -2.43368967048e-05
Gc5_169 0 n10 ns169 0 0.000118493429926
Gc5_170 0 n10 ns170 0 1.0099402119e-05
Gc5_171 0 n10 ns171 0 4.12374908036e-05
Gc5_172 0 n10 ns172 0 0.000379992075518
Gc5_173 0 n10 ns173 0 -0.000689900599877
Gc5_174 0 n10 ns174 0 -0.000406337882737
Gc5_175 0 n10 ns175 0 -0.000231826899362
Gc5_176 0 n10 ns176 0 -0.000674035522729
Gc5_177 0 n10 ns177 0 -0.00167720703208
Gc5_178 0 n10 ns178 0 -0.000495834864986
Gc5_179 0 n10 ns179 0 0.000196774754763
Gc5_180 0 n10 ns180 0 -0.00218335213336
Gc5_181 0 n10 ns181 0 0.000676512343184
Gc5_182 0 n10 ns182 0 0.00104153772084
Gc5_183 0 n10 ns183 0 -0.00067200456148
Gc5_184 0 n10 ns184 0 6.15745161288e-05
Gc5_185 0 n10 ns185 0 0.000911393574616
Gc5_186 0 n10 ns186 0 0.00283151874196
Gc5_187 0 n10 ns187 0 -0.000463035507229
Gc5_188 0 n10 ns188 0 -0.000231569480511
Gc5_189 0 n10 ns189 0 -0.0013447069095
Gc5_190 0 n10 ns190 0 -0.000695903977765
Gc5_191 0 n10 ns191 0 2.84407414933e-05
Gc5_192 0 n10 ns192 0 -0.00422860468662
Gc5_193 0 n10 ns193 0 0.00189834749829
Gc5_194 0 n10 ns194 0 0.00017021823084
Gc5_195 0 n10 ns195 0 0.0019882335804
Gc5_196 0 n10 ns196 0 0.00172910901429
Gc5_197 0 n10 ns197 0 0.000106857541104
Gc5_198 0 n10 ns198 0 2.16027013091e-08
Gc5_199 0 n10 ns199 0 -4.85269232017e-08
Gc5_200 0 n10 ns200 0 -0.00349458238281
Gc5_201 0 n10 ns201 0 -0.0022544854869
Gc5_202 0 n10 ns202 0 0.00842766280008
Gc5_203 0 n10 ns203 0 7.97012799586e-05
Gc5_204 0 n10 ns204 0 -2.983614135e-05
Gc5_205 0 n10 ns205 0 -5.23597367216e-05
Gc5_206 0 n10 ns206 0 0.000495281521284
Gc5_207 0 n10 ns207 0 -0.000204689080058
Gc5_208 0 n10 ns208 0 0.0153852523522
Gc5_209 0 n10 ns209 0 -0.000216882570909
Gc5_210 0 n10 ns210 0 -6.07639011466e-05
Gc5_211 0 n10 ns211 0 1.94627261938e-05
Gc5_212 0 n10 ns212 0 5.89498263858e-05
Gc5_213 0 n10 ns213 0 0.00034139312548
Gc5_214 0 n10 ns214 0 -0.000728090687778
Gc5_215 0 n10 ns215 0 -0.000159383046532
Gc5_216 0 n10 ns216 0 -0.000247302753954
Gc5_217 0 n10 ns217 0 -0.000715210444196
Gc5_218 0 n10 ns218 0 -0.00114180135472
Gc5_219 0 n10 ns219 0 -0.000616402099239
Gc5_220 0 n10 ns220 0 0.000227723916566
Gc5_221 0 n10 ns221 0 -0.0015067726767
Gc5_222 0 n10 ns222 0 0.000157458041127
Gc5_223 0 n10 ns223 0 0.000447971884292
Gc5_224 0 n10 ns224 0 0.00015554427797
Gc5_225 0 n10 ns225 0 5.46298304272e-05
Gc5_226 0 n10 ns226 0 0.00107661706202
Gc5_227 0 n10 ns227 0 0.00210108113258
Gc5_228 0 n10 ns228 0 -0.000157835101192
Gc5_229 0 n10 ns229 0 -0.000297043381923
Gc5_230 0 n10 ns230 0 -0.00156296022472
Gc5_231 0 n10 ns231 0 -0.000355173373648
Gc5_232 0 n10 ns232 0 -0.000248674805423
Gc5_233 0 n10 ns233 0 -0.00352962346973
Gc5_234 0 n10 ns234 0 0.00196380570873
Gc5_235 0 n10 ns235 0 0.000227646090077
Gc5_236 0 n10 ns236 0 0.00221516089013
Gc5_237 0 n10 ns237 0 0.00148122949198
Gc5_238 0 n10 ns238 0 0.000163457169856
Gc5_239 0 n10 ns239 0 -2.41197594749e-09
Gc5_240 0 n10 ns240 0 -2.46462112903e-08
Gc5_241 0 n10 ns241 0 -0.00302121714178
Gc5_242 0 n10 ns242 0 -0.00128694430552
Gc5_243 0 n10 ns243 0 0.00814194497547
Gc5_244 0 n10 ns244 0 4.36514729303e-05
Gc5_245 0 n10 ns245 0 -2.08482352977e-05
Gc5_246 0 n10 ns246 0 -3.10691449195e-05
Gc5_247 0 n10 ns247 0 0.000324362109453
Gc5_248 0 n10 ns248 0 -0.00060665617858
Gc5_249 0 n10 ns249 0 0.00216766102281
Gc5_250 0 n10 ns250 0 -0.000291704305949
Gc5_251 0 n10 ns251 0 -8.40142638813e-05
Gc5_252 0 n10 ns252 0 3.17625564117e-05
Gc5_253 0 n10 ns253 0 1.35643809043e-05
Gc5_254 0 n10 ns254 0 -0.000519359765232
Gc5_255 0 n10 ns255 0 -0.000434917679625
Gc5_256 0 n10 ns256 0 0.000522150705742
Gc5_257 0 n10 ns257 0 5.9387731558e-06
Gc5_258 0 n10 ns258 0 -0.000187188370901
Gc5_259 0 n10 ns259 0 0.00192339120283
Gc5_260 0 n10 ns260 0 -0.000567113931926
Gc5_261 0 n10 ns261 0 0.000121691120549
Gc5_262 0 n10 ns262 0 0.00202275116377
Gc5_263 0 n10 ns263 0 -0.00100884302345
Gc5_264 0 n10 ns264 0 -0.000839408392152
Gc5_265 0 n10 ns265 0 0.00242480890857
Gc5_266 0 n10 ns266 0 3.09405367976e-05
Gc5_267 0 n10 ns267 0 0.000960367992874
Gc5_268 0 n10 ns268 0 -0.00297569701324
Gc5_269 0 n10 ns269 0 0.000375497061495
Gc5_270 0 n10 ns270 0 -0.000278492543444
Gc5_271 0 n10 ns271 0 -0.00130604796225
Gc5_272 0 n10 ns272 0 0.000548430829424
Gc5_273 0 n10 ns273 0 -0.000278576270598
Gc5_274 0 n10 ns274 0 0.00461730548132
Gc5_275 0 n10 ns275 0 -0.000171108608262
Gc5_276 0 n10 ns276 0 -8.79978487622e-06
Gc5_277 0 n10 ns277 0 0.00211938617291
Gc5_278 0 n10 ns278 0 0.000728870812084
Gc5_279 0 n10 ns279 0 -0.00163362506084
Gc5_280 0 n10 ns280 0 -6.98909815683e-08
Gc5_281 0 n10 ns281 0 7.95692991686e-08
Gc5_282 0 n10 ns282 0 0.0036424709915
Gc5_283 0 n10 ns283 0 -0.0012977310869
Gc5_284 0 n10 ns284 0 0.00409855538449
Gc5_285 0 n10 ns285 0 -9.86796006647e-05
Gc5_286 0 n10 ns286 0 7.73304835057e-05
Gc5_287 0 n10 ns287 0 3.66483455664e-05
Gc5_288 0 n10 ns288 0 0.00120623514204
Gc5_289 0 n10 ns289 0 -0.000701146895631
Gc5_290 0 n10 ns290 0 0.011036925741
Gc5_291 0 n10 ns291 0 -0.000632745163888
Gc5_292 0 n10 ns292 0 -0.000362859453148
Gc5_293 0 n10 ns293 0 3.06015025567e-05
Gc5_294 0 n10 ns294 0 6.18126183452e-05
Gc5_295 0 n10 ns295 0 -2.3371889059e-05
Gc5_296 0 n10 ns296 0 -0.0005736784562
Gc5_297 0 n10 ns297 0 0.000396750952063
Gc5_298 0 n10 ns298 0 -6.80616091732e-05
Gc5_299 0 n10 ns299 0 -0.000931945983805
Gc5_300 0 n10 ns300 0 0.000809905746623
Gc5_301 0 n10 ns301 0 -0.000645100691636
Gc5_302 0 n10 ns302 0 0.000166082088785
Gc5_303 0 n10 ns303 0 0.00110724059989
Gc5_304 0 n10 ns304 0 -0.00041560375445
Gc5_305 0 n10 ns305 0 -0.00165175755395
Gc5_306 0 n10 ns306 0 0.00230241894136
Gc5_307 0 n10 ns307 0 3.26728126437e-05
Gc5_308 0 n10 ns308 0 0.00115016415942
Gc5_309 0 n10 ns309 0 -0.00183139608
Gc5_310 0 n10 ns310 0 -0.000487526574934
Gc5_311 0 n10 ns311 0 -0.000416682548475
Gc5_312 0 n10 ns312 0 -0.00151532214369
Gc5_313 0 n10 ns313 0 0.00128474255598
Gc5_314 0 n10 ns314 0 -0.000313138420363
Gc5_315 0 n10 ns315 0 0.00252551350316
Gc5_316 0 n10 ns316 0 0.000991363552516
Gc5_317 0 n10 ns317 0 0.000278903238866
Gc5_318 0 n10 ns318 0 0.00237401749475
Gc5_319 0 n10 ns319 0 -0.000944119680335
Gc5_320 0 n10 ns320 0 -0.00196064299427
Gc5_321 0 n10 ns321 0 -4.70603062739e-08
Gc5_322 0 n10 ns322 0 9.6086558294e-08
Gc5_323 0 n10 ns323 0 0.00326683303185
Gc5_324 0 n10 ns324 0 -0.000783185852075
Gc5_325 0 n10 ns325 0 0.00493174616885
Gc5_326 0 n10 ns326 0 -0.000138234781516
Gc5_327 0 n10 ns327 0 0.00011636055543
Gc5_328 0 n10 ns328 0 4.25857057843e-05
Gd5_1 0 n10 ni1 0 7.49367442558e-05
Gd5_2 0 n10 ni2 0 -0.000649234280069
Gd5_3 0 n10 ni3 0 0.000741517556032
Gd5_4 0 n10 ni4 0 0.000139154663073
Gd5_5 0 n10 ni5 0 -0.00184255616824
Gd5_6 0 n10 ni6 0 -0.00209423907569
Gd5_7 0 n10 ni7 0 -0.000990163718501
Gd5_8 0 n10 ni8 0 -0.00325987892274
Gc6_1 0 n12 ns1 0 0.000129489175019
Gc6_2 0 n12 ns2 0 -0.000269648922389
Gc6_3 0 n12 ns3 0 0.00371902787721
Gc6_4 0 n12 ns4 0 -0.000714357935815
Gc6_5 0 n12 ns5 0 -0.000129804636225
Gc6_6 0 n12 ns6 0 8.16105484995e-05
Gc6_7 0 n12 ns7 0 5.70633215505e-05
Gc6_8 0 n12 ns8 0 -0.000744792315097
Gc6_9 0 n12 ns9 0 -0.00133965091728
Gc6_10 0 n12 ns10 0 0.000732360786287
Gc6_11 0 n12 ns11 0 -0.000142450203608
Gc6_12 0 n12 ns12 0 -0.000379192261636
Gc6_13 0 n12 ns13 0 -0.00236207716482
Gc6_14 0 n12 ns14 0 0.000668077300499
Gc6_15 0 n12 ns15 0 -0.000123432273529
Gc6_16 0 n12 ns16 0 -0.00170806728841
Gc6_17 0 n12 ns17 0 0.000644736404578
Gc6_18 0 n12 ns18 0 -0.000792624219036
Gc6_19 0 n12 ns19 0 0.00902109108902
Gc6_20 0 n12 ns20 0 2.99212778579e-05
Gc6_21 0 n12 ns21 0 0.00112254622498
Gc6_22 0 n12 ns22 0 -0.0012137773644
Gc6_23 0 n12 ns23 0 0.000895049428534
Gc6_24 0 n12 ns24 0 0.000331214686571
Gc6_25 0 n12 ns25 0 0.00143144166507
Gc6_26 0 n12 ns26 0 -0.00180690871172
Gc6_27 0 n12 ns27 0 0.00203602157383
Gc6_28 0 n12 ns28 0 2.114847143e-06
Gc6_29 0 n12 ns29 0 0.00597784861346
Gc6_30 0 n12 ns30 0 2.71194275715e-06
Gc6_31 0 n12 ns31 0 0.00150016479062
Gc6_32 0 n12 ns32 0 -0.0019979551248
Gc6_33 0 n12 ns33 0 0.00588831517778
Gc6_34 0 n12 ns34 0 7.03903896872e-08
Gc6_35 0 n12 ns35 0 5.69689878337e-08
Gc6_36 0 n12 ns36 0 -0.00170578868435
Gc6_37 0 n12 ns37 0 -0.0056954856485
Gc6_38 0 n12 ns38 0 -0.00380621505725
Gc6_39 0 n12 ns39 0 9.79074802349e-06
Gc6_40 0 n12 ns40 0 3.57341931489e-07
Gc6_41 0 n12 ns41 0 -1.96093820168e-05
Gc6_42 0 n12 ns42 0 -0.000123587860593
Gc6_43 0 n12 ns43 0 0.00193830285097
Gc6_44 0 n12 ns44 0 0.00398252628648
Gc6_45 0 n12 ns45 0 0.00035881517251
Gc6_46 0 n12 ns46 0 -4.07963603821e-05
Gc6_47 0 n12 ns47 0 -2.41004626061e-05
Gc6_48 0 n12 ns48 0 1.22616438303e-05
Gc6_49 0 n12 ns49 0 0.000665376292683
Gc6_50 0 n12 ns50 0 -0.000394280642633
Gc6_51 0 n12 ns51 0 -1.12847363992e-05
Gc6_52 0 n12 ns52 0 0.000114477614005
Gc6_53 0 n12 ns53 0 -0.000941154297219
Gc6_54 0 n12 ns54 0 0.00341705148766
Gc6_55 0 n12 ns55 0 0.000912896961929
Gc6_56 0 n12 ns56 0 -0.000299117189324
Gc6_57 0 n12 ns57 0 -0.000809481190016
Gc6_58 0 n12 ns58 0 -0.000759467742538
Gc6_59 0 n12 ns59 0 -0.000924355804593
Gc6_60 0 n12 ns60 0 -0.0092403403253
Gc6_61 0 n12 ns61 0 6.47362103748e-05
Gc6_62 0 n12 ns62 0 0.0011787791211
Gc6_63 0 n12 ns63 0 -0.00187943357477
Gc6_64 0 n12 ns64 0 -0.00091012302846
Gc6_65 0 n12 ns65 0 8.84621943249e-05
Gc6_66 0 n12 ns66 0 0.00191192274769
Gc6_67 0 n12 ns67 0 0.00307453566836
Gc6_68 0 n12 ns68 0 -0.00352545962015
Gc6_69 0 n12 ns69 0 -0.00797890169391
Gc6_70 0 n12 ns70 0 -0.00413568245491
Gc6_71 0 n12 ns71 0 0.000514530360072
Gc6_72 0 n12 ns72 0 0.00404920677089
Gc6_73 0 n12 ns73 0 0.00423377738386
Gc6_74 0 n12 ns74 0 -0.0107401262124
Gc6_75 0 n12 ns75 0 -1.99104965163e-07
Gc6_76 0 n12 ns76 0 -2.42524385996e-08
Gc6_77 0 n12 ns77 0 0.00676824944206
Gc6_78 0 n12 ns78 0 0.00555048003007
Gc6_79 0 n12 ns79 0 -0.0116614758185
Gc6_80 0 n12 ns80 0 -0.000178986442757
Gc6_81 0 n12 ns81 0 0.000187894610478
Gc6_82 0 n12 ns82 0 7.31872304287e-05
Gc6_83 0 n12 ns83 0 0.000120947911102
Gc6_84 0 n12 ns84 0 0.00141984461112
Gc6_85 0 n12 ns85 0 0.00306340773653
Gc6_86 0 n12 ns86 0 -3.74660222597e-05
Gc6_87 0 n12 ns87 0 0.000623229455654
Gc6_88 0 n12 ns88 0 5.86272214832e-05
Gc6_89 0 n12 ns89 0 -3.69500763462e-06
Gc6_90 0 n12 ns90 0 -0.000275308546567
Gc6_91 0 n12 ns91 0 -0.000256422508427
Gc6_92 0 n12 ns92 0 -0.000252661652814
Gc6_93 0 n12 ns93 0 -0.000298500820954
Gc6_94 0 n12 ns94 0 -0.00142977632434
Gc6_95 0 n12 ns95 0 -0.00120053307886
Gc6_96 0 n12 ns96 0 0.000777804549501
Gc6_97 0 n12 ns97 0 -0.000138856383914
Gc6_98 0 n12 ns98 0 0.00141145895975
Gc6_99 0 n12 ns99 0 -0.000596383799998
Gc6_100 0 n12 ns100 0 -0.000671282333253
Gc6_101 0 n12 ns101 0 0.00211242282773
Gc6_102 0 n12 ns102 0 1.57095744471e-05
Gc6_103 0 n12 ns103 0 0.00109437459613
Gc6_104 0 n12 ns104 0 0.00260594385463
Gc6_105 0 n12 ns105 0 -0.000329667634287
Gc6_106 0 n12 ns106 0 0.000206153628218
Gc6_107 0 n12 ns107 0 0.0015160363636
Gc6_108 0 n12 ns108 0 0.000280119168932
Gc6_109 0 n12 ns109 0 -0.000338883024379
Gc6_110 0 n12 ns110 0 0.00378606993495
Gc6_111 0 n12 ns111 0 0.00190296327941
Gc6_112 0 n12 ns112 0 7.97932406304e-05
Gc6_113 0 n12 ns113 0 0.00211858744469
Gc6_114 0 n12 ns114 0 5.95420400541e-05
Gc6_115 0 n12 ns115 0 0.000695606651034
Gc6_116 0 n12 ns116 0 -2.44799807122e-08
Gc6_117 0 n12 ns117 0 6.75831042215e-08
Gc6_118 0 n12 ns118 0 -0.00338132161839
Gc6_119 0 n12 ns119 0 -0.00300610472727
Gc6_120 0 n12 ns120 0 -0.00266091347075
Gc6_121 0 n12 ns121 0 5.70513532958e-05
Gc6_122 0 n12 ns122 0 -2.16848079745e-05
Gc6_123 0 n12 ns123 0 -4.86544349762e-05
Gc6_124 0 n12 ns124 0 -4.21264493587e-05
Gc6_125 0 n12 ns125 0 0.00124622577034
Gc6_126 0 n12 ns126 0 0.00407799811713
Gc6_127 0 n12 ns127 0 -0.000330812734768
Gc6_128 0 n12 ns128 0 0.000204660703836
Gc6_129 0 n12 ns129 0 7.2380520363e-05
Gc6_130 0 n12 ns130 0 4.6895224594e-05
Gc6_131 0 n12 ns131 0 -0.000204041343398
Gc6_132 0 n12 ns132 0 -0.000966968504818
Gc6_133 0 n12 ns133 0 3.55739985402e-05
Gc6_134 0 n12 ns134 0 -0.000281889470201
Gc6_135 0 n12 ns135 0 -0.000609212431353
Gc6_136 0 n12 ns136 0 -0.00128822938175
Gc6_137 0 n12 ns137 0 0.000890256315823
Gc6_138 0 n12 ns138 0 -0.000198484766575
Gc6_139 0 n12 ns139 0 0.000752281994948
Gc6_140 0 n12 ns140 0 -0.000380875328529
Gc6_141 0 n12 ns141 0 -0.00268074065951
Gc6_142 0 n12 ns142 0 0.00359390729721
Gc6_143 0 n12 ns143 0 -1.59467418777e-05
Gc6_144 0 n12 ns144 0 0.00126913012138
Gc6_145 0 n12 ns145 0 0.00211979390226
Gc6_146 0 n12 ns146 0 2.2591155994e-05
Gc6_147 0 n12 ns147 0 0.000204548171007
Gc6_148 0 n12 ns148 0 0.00174662384852
Gc6_149 0 n12 ns149 0 -6.77781407414e-05
Gc6_150 0 n12 ns150 0 -0.000359136691485
Gc6_151 0 n12 ns151 0 0.00281104571156
Gc6_152 0 n12 ns152 0 0.0037077751706
Gc6_153 0 n12 ns153 0 0.000174675068166
Gc6_154 0 n12 ns154 0 0.00221810102207
Gc6_155 0 n12 ns155 0 -0.000902599558008
Gc6_156 0 n12 ns156 0 0.00207796709637
Gc6_157 0 n12 ns157 0 3.9598359273e-09
Gc6_158 0 n12 ns158 0 7.66605704375e-08
Gc6_159 0 n12 ns159 0 -0.00354740374639
Gc6_160 0 n12 ns160 0 -0.00360204044736
Gc6_161 0 n12 ns161 0 -0.00370562126954
Gc6_162 0 n12 ns162 0 3.49531198388e-05
Gc6_163 0 n12 ns163 0 -3.57372052321e-06
Gc6_164 0 n12 ns164 0 -4.06190476565e-05
Gc6_165 0 n12 ns165 0 0.000495281525998
Gc6_166 0 n12 ns166 0 -0.000204689070774
Gc6_167 0 n12 ns167 0 0.0153852523555
Gc6_168 0 n12 ns168 0 -0.000216882572203
Gc6_169 0 n12 ns169 0 -6.07639055084e-05
Gc6_170 0 n12 ns170 0 1.94627249367e-05
Gc6_171 0 n12 ns171 0 5.89498271053e-05
Gc6_172 0 n12 ns172 0 0.000341393121441
Gc6_173 0 n12 ns173 0 -0.000728090683132
Gc6_174 0 n12 ns174 0 -0.000159383049373
Gc6_175 0 n12 ns175 0 -0.00024730275288
Gc6_176 0 n12 ns176 0 -0.00071521043377
Gc6_177 0 n12 ns177 0 -0.00114180134645
Gc6_178 0 n12 ns178 0 -0.000616402100012
Gc6_179 0 n12 ns179 0 0.000227723915903
Gc6_180 0 n12 ns180 0 -0.00150677267583
Gc6_181 0 n12 ns181 0 0.000157458044827
Gc6_182 0 n12 ns182 0 0.000447971901331
Gc6_183 0 n12 ns183 0 0.000155544270063
Gc6_184 0 n12 ns184 0 5.46298311858e-05
Gc6_185 0 n12 ns185 0 0.00107661706192
Gc6_186 0 n12 ns186 0 0.00210108112779
Gc6_187 0 n12 ns187 0 -0.000157835100473
Gc6_188 0 n12 ns188 0 -0.000297043380639
Gc6_189 0 n12 ns189 0 -0.00156296022431
Gc6_190 0 n12 ns190 0 -0.000355173380561
Gc6_191 0 n12 ns191 0 -0.000248674798619
Gc6_192 0 n12 ns192 0 -0.0035296234603
Gc6_193 0 n12 ns193 0 0.00196380569781
Gc6_194 0 n12 ns194 0 0.000227646089537
Gc6_195 0 n12 ns195 0 0.00221516089217
Gc6_196 0 n12 ns196 0 0.0014812295013
Gc6_197 0 n12 ns197 0 0.000163457164095
Gc6_198 0 n12 ns198 0 -2.41197720888e-09
Gc6_199 0 n12 ns199 0 -2.46462118039e-08
Gc6_200 0 n12 ns200 0 -0.00302121713564
Gc6_201 0 n12 ns201 0 -0.00128694431861
Gc6_202 0 n12 ns202 0 0.00814194498623
Gc6_203 0 n12 ns203 0 4.36514697061e-05
Gc6_204 0 n12 ns204 0 -2.08482357413e-05
Gc6_205 0 n12 ns205 0 -3.10691432941e-05
Gc6_206 0 n12 ns206 0 -0.000248061743979
Gc6_207 0 n12 ns207 0 0.000574508320747
Gc6_208 0 n12 ns208 0 0.0109394345032
Gc6_209 0 n12 ns209 0 0.00011313440144
Gc6_210 0 n12 ns210 0 0.000132047954668
Gc6_211 0 n12 ns211 0 2.38801194699e-05
Gc6_212 0 n12 ns212 0 3.34391501625e-05
Gc6_213 0 n12 ns213 0 0.000182240206033
Gc6_214 0 n12 ns214 0 -0.000687289681468
Gc6_215 0 n12 ns215 0 -4.72862993886e-05
Gc6_216 0 n12 ns216 0 -0.000153314770856
Gc6_217 0 n12 ns217 0 -0.000269611333282
Gc6_218 0 n12 ns218 0 -0.00108148009898
Gc6_219 0 n12 ns219 0 -0.000796505408473
Gc6_220 0 n12 ns220 0 0.000274871393398
Gc6_221 0 n12 ns221 0 -0.000971998838248
Gc6_222 0 n12 ns222 0 2.94851595258e-05
Gc6_223 0 n12 ns223 0 0.000295668429573
Gc6_224 0 n12 ns224 0 -0.000323478558784
Gc6_225 0 n12 ns225 0 8.50042647249e-05
Gc6_226 0 n12 ns226 0 0.00125780157946
Gc6_227 0 n12 ns227 0 0.0012853824224
Gc6_228 0 n12 ns228 0 -0.000101561042243
Gc6_229 0 n12 ns229 0 -0.000266838421658
Gc6_230 0 n12 ns230 0 -0.00179214916525
Gc6_231 0 n12 ns231 0 -7.77264794637e-05
Gc6_232 0 n12 ns232 0 0.000301582837911
Gc6_233 0 n12 ns233 0 -0.0022902950266
Gc6_234 0 n12 ns234 0 0.00122707044039
Gc6_235 0 n12 ns235 0 0.000198667827487
Gc6_236 0 n12 ns236 0 0.00291833447563
Gc6_237 0 n12 ns237 0 0.000917876856001
Gc6_238 0 n12 ns238 0 -0.000896267773204
Gc6_239 0 n12 ns239 0 -5.43116247618e-08
Gc6_240 0 n12 ns240 0 -1.20902145373e-07
Gc6_241 0 n12 ns241 0 -0.00151650124501
Gc6_242 0 n12 ns242 0 -0.00128937534882
Gc6_243 0 n12 ns243 0 0.00872445052881
Gc6_244 0 n12 ns244 0 7.05150102776e-05
Gc6_245 0 n12 ns245 0 -5.1005148678e-05
Gc6_246 0 n12 ns246 0 -4.45283096759e-05
Gc6_247 0 n12 ns247 0 0.00121253289374
Gc6_248 0 n12 ns248 0 -0.000689662101094
Gc6_249 0 n12 ns249 0 0.0109394728908
Gc6_250 0 n12 ns250 0 -0.0006333293318
Gc6_251 0 n12 ns251 0 -0.000382151145758
Gc6_252 0 n12 ns252 0 2.6750991093e-05
Gc6_253 0 n12 ns253 0 6.31036366294e-05
Gc6_254 0 n12 ns254 0 -3.60786157554e-05
Gc6_255 0 n12 ns255 0 -0.000555524757844
Gc6_256 0 n12 ns256 0 0.000380665662121
Gc6_257 0 n12 ns257 0 -6.44543007327e-05
Gc6_258 0 n12 ns258 0 -0.00087919692221
Gc6_259 0 n12 ns259 0 0.000849630266216
Gc6_260 0 n12 ns260 0 -0.000647263365503
Gc6_261 0 n12 ns261 0 0.000158480204586
Gc6_262 0 n12 ns262 0 0.00112257812599
Gc6_263 0 n12 ns263 0 -0.000392131666555
Gc6_264 0 n12 ns264 0 -0.00160246994266
Gc6_265 0 n12 ns265 0 0.00223507664274
Gc6_266 0 n12 ns266 0 3.10546072525e-05
Gc6_267 0 n12 ns267 0 0.00114436418797
Gc6_268 0 n12 ns268 0 -0.00185056170905
Gc6_269 0 n12 ns269 0 -0.000488949154909
Gc6_270 0 n12 ns270 0 -0.000404274175596
Gc6_271 0 n12 ns271 0 -0.00151259621893
Gc6_272 0 n12 ns272 0 0.00127252030007
Gc6_273 0 n12 ns273 0 -0.000279632428133
Gc6_274 0 n12 ns274 0 0.00256104415776
Gc6_275 0 n12 ns275 0 0.000966686477443
Gc6_276 0 n12 ns276 0 0.000267621654314
Gc6_277 0 n12 ns277 0 0.00238224840873
Gc6_278 0 n12 ns278 0 -0.000909821171191
Gc6_279 0 n12 ns279 0 -0.00198197356868
Gc6_280 0 n12 ns280 0 -4.79262159019e-08
Gc6_281 0 n12 ns281 0 9.37937347677e-08
Gc6_282 0 n12 ns282 0 0.00329373639474
Gc6_283 0 n12 ns283 0 -0.000810754537099
Gc6_284 0 n12 ns284 0 0.00495834656159
Gc6_285 0 n12 ns285 0 -0.000142957321081
Gc6_286 0 n12 ns286 0 0.000119636693564
Gc6_287 0 n12 ns287 0 4.30569936451e-05
Gc6_288 0 n12 ns288 0 0.00066212958912
Gc6_289 0 n12 ns289 0 -0.000369696464725
Gc6_290 0 n12 ns290 0 0.00972225379514
Gc6_291 0 n12 ns291 0 -0.000348095878004
Gc6_292 0 n12 ns292 0 -4.96526858458e-05
Gc6_293 0 n12 ns293 0 2.90009744621e-05
Gc6_294 0 n12 ns294 0 3.73307773955e-05
Gc6_295 0 n12 ns295 0 -0.000179796544328
Gc6_296 0 n12 ns296 0 -0.000817420213559
Gc6_297 0 n12 ns297 0 0.000285743497911
Gc6_298 0 n12 ns298 0 -8.47263484003e-05
Gc6_299 0 n12 ns299 0 -0.000802924228797
Gc6_300 0 n12 ns300 0 0.000889451931185
Gc6_301 0 n12 ns301 0 -0.000758690771008
Gc6_302 0 n12 ns302 0 0.000225099189711
Gc6_303 0 n12 ns303 0 0.000803868094186
Gc6_304 0 n12 ns304 0 -0.000401908835088
Gc6_305 0 n12 ns305 0 -0.000281879688966
Gc6_306 0 n12 ns306 0 0.0021766814463
Gc6_307 0 n12 ns307 0 3.65721717261e-05
Gc6_308 0 n12 ns308 0 0.00128945198927
Gc6_309 0 n12 ns309 0 -0.00138694510793
Gc6_310 0 n12 ns310 0 -0.000124285585727
Gc6_311 0 n12 ns311 0 -0.000321892538021
Gc6_312 0 n12 ns312 0 -0.00175130119617
Gc6_313 0 n12 ns313 0 8.16695906437e-05
Gc6_314 0 n12 ns314 0 -0.000589309309673
Gc6_315 0 n12 ns315 0 0.00212975008263
Gc6_316 0 n12 ns316 0 0.00155856806869
Gc6_317 0 n12 ns317 0 9.55342150734e-05
Gc6_318 0 n12 ns318 0 0.00257077673645
Gc6_319 0 n12 ns319 0 0.00133664399051
Gc6_320 0 n12 ns320 0 -0.000111140925866
Gc6_321 0 n12 ns321 0 -4.74472647123e-09
Gc6_322 0 n12 ns322 0 2.92726314545e-08
Gc6_323 0 n12 ns323 0 0.0014883062119
Gc6_324 0 n12 ns324 0 -0.000218013240129
Gc6_325 0 n12 ns325 0 0.00614779661239
Gc6_326 0 n12 ns326 0 -3.3877518795e-05
Gc6_327 0 n12 ns327 0 2.56587012835e-05
Gc6_328 0 n12 ns328 0 1.74219769129e-05
Gd6_1 0 n12 ni1 0 -0.000656344066429
Gd6_2 0 n12 ni2 0 -0.000135924976124
Gd6_3 0 n12 ni3 0 0.000154238123033
Gd6_4 0 n12 ni4 0 -6.21146557827e-05
Gd6_5 0 n12 ni5 0 -0.00209423907492
Gd6_6 0 n12 ni6 0 -0.00037423051667
Gd6_7 0 n12 ni7 0 -0.00323273116678
Gd6_8 0 n12 ni8 0 -0.00203460583981
Gc7_1 0 n14 ns1 0 -0.000164789774213
Gc7_2 0 n14 ns2 0 0.00225479908976
Gc7_3 0 n14 ns3 0 0.00249658822831
Gc7_4 0 n14 ns4 0 0.000255505806472
Gc7_5 0 n14 ns5 0 0.000598839350772
Gc7_6 0 n14 ns6 0 2.87394942962e-05
Gc7_7 0 n14 ns7 0 -9.40368767886e-06
Gc7_8 0 n14 ns8 0 0.000230669074535
Gc7_9 0 n14 ns9 0 -0.000146086563074
Gc7_10 0 n14 ns10 0 -0.000530876076723
Gc7_11 0 n14 ns11 0 -0.000187631373707
Gc7_12 0 n14 ns12 0 -0.00118079984034
Gc7_13 0 n14 ns13 0 -0.000641558783504
Gc7_14 0 n14 ns14 0 0.000693286735393
Gc7_15 0 n14 ns15 0 -0.000122300842245
Gc7_16 0 n14 ns16 0 0.00206095268867
Gc7_17 0 n14 ns17 0 -0.00131207362164
Gc7_18 0 n14 ns18 0 -0.00200806842003
Gc7_19 0 n14 ns19 0 -0.000315648791341
Gc7_20 0 n14 ns20 0 -8.25133868237e-06
Gc7_21 0 n14 ns21 0 0.000936197622992
Gc7_22 0 n14 ns22 0 0.00341868913621
Gc7_23 0 n14 ns23 0 -0.000811476938034
Gc7_24 0 n14 ns24 0 0.000132122136811
Gc7_25 0 n14 ns25 0 0.00131840895953
Gc7_26 0 n14 ns26 0 0.000797156516306
Gc7_27 0 n14 ns27 0 -0.00122822213962
Gc7_28 0 n14 ns28 0 0.00396331298329
Gc7_29 0 n14 ns29 0 0.000327001356588
Gc7_30 0 n14 ns30 0 0.000183650390118
Gc7_31 0 n14 ns31 0 0.0020308096742
Gc7_32 0 n14 ns32 0 0.000300725123798
Gc7_33 0 n14 ns33 0 -0.00132002347953
Gc7_34 0 n14 ns34 0 -4.36399376341e-08
Gc7_35 0 n14 ns35 0 5.67319358318e-08
Gc7_36 0 n14 ns36 0 -0.00321547352171
Gc7_37 0 n14 ns37 0 -0.00239322045496
Gc7_38 0 n14 ns38 0 -0.00152042552102
Gc7_39 0 n14 ns39 0 7.13379317053e-05
Gc7_40 0 n14 ns40 0 -3.68791455785e-05
Gc7_41 0 n14 ns41 0 -5.01194754548e-05
Gc7_42 0 n14 ns42 0 0.000120368773815
Gc7_43 0 n14 ns43 0 0.00141761586398
Gc7_44 0 n14 ns44 0 0.00308861967137
Gc7_45 0 n14 ns45 0 -3.81441411517e-05
Gc7_46 0 n14 ns46 0 0.00062599345617
Gc7_47 0 n14 ns47 0 5.95306152388e-05
Gc7_48 0 n14 ns48 0 -3.72215822815e-06
Gc7_49 0 n14 ns49 0 -0.000271030752904
Gc7_50 0 n14 ns50 0 -0.000259157971588
Gc7_51 0 n14 ns51 0 -0.000249159545869
Gc7_52 0 n14 ns52 0 -0.000298273534642
Gc7_53 0 n14 ns53 0 -0.00144072401545
Gc7_54 0 n14 ns54 0 -0.00121085252525
Gc7_55 0 n14 ns55 0 0.000778751340862
Gc7_56 0 n14 ns56 0 -0.000138389216264
Gc7_57 0 n14 ns57 0 0.00140967167252
Gc7_58 0 n14 ns58 0 -0.000599319347625
Gc7_59 0 n14 ns59 0 -0.0006894048937
Gc7_60 0 n14 ns60 0 0.00211955395545
Gc7_61 0 n14 ns61 0 1.51499481024e-05
Gc7_62 0 n14 ns62 0 0.00109400144587
Gc7_63 0 n14 ns63 0 0.00261002578916
Gc7_64 0 n14 ns64 0 -0.000328899157211
Gc7_65 0 n14 ns65 0 0.000205365764117
Gc7_66 0 n14 ns66 0 0.00151413033107
Gc7_67 0 n14 ns67 0 0.000290605468549
Gc7_68 0 n14 ns68 0 -0.000346488611048
Gc7_69 0 n14 ns69 0 0.00377593597089
Gc7_70 0 n14 ns70 0 0.00191056093379
Gc7_71 0 n14 ns71 0 8.0235838068e-05
Gc7_72 0 n14 ns72 0 0.00211760695356
Gc7_73 0 n14 ns73 0 5.0862435586e-05
Gc7_74 0 n14 ns74 0 0.000693789338453
Gc7_75 0 n14 ns75 0 -2.33221446953e-08
Gc7_76 0 n14 ns76 0 6.72235317159e-08
Gc7_77 0 n14 ns77 0 -0.00338153930346
Gc7_78 0 n14 ns78 0 -0.00301873077655
Gc7_79 0 n14 ns79 0 -0.00265158110305
Gc7_80 0 n14 ns80 0 5.7836147229e-05
Gc7_81 0 n14 ns81 0 -2.02627160937e-05
Gc7_82 0 n14 ns82 0 -4.90081618892e-05
Gc7_83 0 n14 ns83 0 -0.000324421346359
Gc7_84 0 n14 ns84 0 0.00118334923666
Gc7_85 0 n14 ns85 0 0.00190977834418
Gc7_86 0 n14 ns86 0 0.000244622141316
Gc7_87 0 n14 ns87 0 -0.00041354646487
Gc7_88 0 n14 ns88 0 -2.02530699206e-05
Gc7_89 0 n14 ns89 0 2.56816635501e-05
Gc7_90 0 n14 ns90 0 0.000651798391208
Gc7_91 0 n14 ns91 0 -0.000703716344799
Gc7_92 0 n14 ns92 0 0.000456184165459
Gc7_93 0 n14 ns93 0 0.000152555133722
Gc7_94 0 n14 ns94 0 3.7509960909e-05
Gc7_95 0 n14 ns95 0 0.00368185821184
Gc7_96 0 n14 ns96 0 0.000591758497084
Gc7_97 0 n14 ns97 0 -0.000233364403572
Gc7_98 0 n14 ns98 0 -0.00205880142396
Gc7_99 0 n14 ns99 0 0.000174107856603
Gc7_100 0 n14 ns100 0 -0.00101899084227
Gc7_101 0 n14 ns101 0 -0.00872636889348
Gc7_102 0 n14 ns102 0 6.32515970403e-05
Gc7_103 0 n14 ns103 0 0.00081291508865
Gc7_104 0 n14 ns104 0 -0.00362540454218
Gc7_105 0 n14 ns105 0 -0.00024497929658
Gc7_106 0 n14 ns106 0 0.000108412629439
Gc7_107 0 n14 ns107 0 0.00148314227629
Gc7_108 0 n14 ns108 0 0.00227404583714
Gc7_109 0 n14 ns109 0 -0.0032124229938
Gc7_110 0 n14 ns110 0 -0.00945958934931
Gc7_111 0 n14 ns111 0 -0.00345308323894
Gc7_112 0 n14 ns112 0 0.000439393337869
Gc7_113 0 n14 ns113 0 0.00323065176437
Gc7_114 0 n14 ns114 0 0.00444676262254
Gc7_115 0 n14 ns115 0 -0.0100174333773
Gc7_116 0 n14 ns116 0 -2.15270976872e-07
Gc7_117 0 n14 ns117 0 3.66329865786e-08
Gc7_118 0 n14 ns118 0 0.00839809988806
Gc7_119 0 n14 ns119 0 0.00654215575589
Gc7_120 0 n14 ns120 0 -0.0112924053454
Gc7_121 0 n14 ns121 0 -0.000169189624488
Gc7_122 0 n14 ns122 0 0.000173093219065
Gc7_123 0 n14 ns123 0 7.85690359958e-05
Gc7_124 0 n14 ns124 0 0.000121344644563
Gc7_125 0 n14 ns125 0 -0.000325961881356
Gc7_126 0 n14 ns126 0 0.00359742454546
Gc7_127 0 n14 ns127 0 -0.000708945403313
Gc7_128 0 n14 ns128 0 -0.000121411774492
Gc7_129 0 n14 ns129 0 8.30292420296e-05
Gc7_130 0 n14 ns130 0 5.75277009093e-05
Gc7_131 0 n14 ns131 0 -0.000744476639593
Gc7_132 0 n14 ns132 0 -0.0013349394887
Gc7_133 0 n14 ns133 0 0.000733789847212
Gc7_134 0 n14 ns134 0 -0.000136224412547
Gc7_135 0 n14 ns135 0 -0.000359711974394
Gc7_136 0 n14 ns136 0 -0.00238177555603
Gc7_137 0 n14 ns137 0 0.000662863241749
Gc7_138 0 n14 ns138 0 -0.000117838014376
Gc7_139 0 n14 ns139 0 -0.00170325184172
Gc7_140 0 n14 ns140 0 0.000644986542995
Gc7_141 0 n14 ns141 0 -0.000831056445457
Gc7_142 0 n14 ns142 0 0.00899710467626
Gc7_143 0 n14 ns143 0 2.52737812013e-05
Gc7_144 0 n14 ns144 0 0.00111478812048
Gc7_145 0 n14 ns145 0 -0.00120147506737
Gc7_146 0 n14 ns146 0 0.000900661474699
Gc7_147 0 n14 ns147 0 0.000318546828185
Gc7_148 0 n14 ns148 0 0.00142539155108
Gc7_149 0 n14 ns149 0 -0.0018011168298
Gc7_150 0 n14 ns150 0 0.0020139448441
Gc7_151 0 n14 ns151 0 -1.71427624552e-05
Gc7_152 0 n14 ns152 0 0.00602797193706
Gc7_153 0 n14 ns153 0 -1.08946895933e-06
Gc7_154 0 n14 ns154 0 0.00148641972662
Gc7_155 0 n14 ns155 0 -0.00202043688293
Gc7_156 0 n14 ns156 0 0.00595636327157
Gc7_157 0 n14 ns157 0 6.94707118822e-08
Gc7_158 0 n14 ns158 0 5.62805782098e-08
Gc7_159 0 n14 ns159 0 -0.00171154846984
Gc7_160 0 n14 ns160 0 -0.00560078748706
Gc7_161 0 n14 ns161 0 -0.00387361140057
Gc7_162 0 n14 ns162 0 1.36841946327e-05
Gc7_163 0 n14 ns163 0 -6.00777093048e-06
Gc7_164 0 n14 ns164 0 -2.21376729585e-05
Gc7_165 0 n14 ns165 0 0.000324362137473
Gc7_166 0 n14 ns166 0 -0.000606656079973
Gc7_167 0 n14 ns167 0 0.0021676611189
Gc7_168 0 n14 ns168 0 -0.000291704321586
Gc7_169 0 n14 ns169 0 -8.40142987774e-05
Gc7_170 0 n14 ns170 0 3.17625516104e-05
Gc7_171 0 n14 ns171 0 1.35643820452e-05
Gc7_172 0 n14 ns172 0 -0.000519359778069
Gc7_173 0 n14 ns173 0 -0.000434917649429
Gc7_174 0 n14 ns174 0 0.000522150692533
Gc7_175 0 n14 ns175 0 5.93878295148e-06
Gc7_176 0 n14 ns176 0 -0.00018718830389
Gc7_177 0 n14 ns177 0 0.00192339123311
Gc7_178 0 n14 ns178 0 -0.000567113937368
Gc7_179 0 n14 ns179 0 0.000121691117493
Gc7_180 0 n14 ns180 0 0.00202275117407
Gc7_181 0 n14 ns181 0 -0.0010088430097
Gc7_182 0 n14 ns182 0 -0.000839408327995
Gc7_183 0 n14 ns183 0 0.00242480884862
Gc7_184 0 n14 ns184 0 3.0940540296e-05
Gc7_185 0 n14 ns185 0 0.000960367992309
Gc7_186 0 n14 ns186 0 -0.00297569703253
Gc7_187 0 n14 ns187 0 0.000375497077652
Gc7_188 0 n14 ns188 0 -0.000278492535277
Gc7_189 0 n14 ns189 0 -0.00130604796512
Gc7_190 0 n14 ns190 0 0.000548430843322
Gc7_191 0 n14 ns191 0 -0.000278576229527
Gc7_192 0 n14 ns192 0 0.0046173054045
Gc7_193 0 n14 ns193 0 -0.000171108652494
Gc7_194 0 n14 ns194 0 -8.79975008652e-06
Gc7_195 0 n14 ns195 0 0.00211938617895
Gc7_196 0 n14 ns196 0 0.00072887070488
Gc7_197 0 n14 ns197 0 -0.00163362502969
Gc7_198 0 n14 ns198 0 -6.98909864829e-08
Gc7_199 0 n14 ns199 0 7.95692848354e-08
Gc7_200 0 n14 ns200 0 0.00364247096763
Gc7_201 0 n14 ns201 0 -0.00129773086077
Gc7_202 0 n14 ns202 0 0.00409855526674
Gc7_203 0 n14 ns203 0 -9.86796288682e-05
Gc7_204 0 n14 ns204 0 7.73304846838e-05
Gc7_205 0 n14 ns205 0 3.66483473045e-05
Gc7_206 0 n14 ns206 0 0.00121253289034
Gc7_207 0 n14 ns207 0 -0.000689662100133
Gc7_208 0 n14 ns208 0 0.0109394729162
Gc7_209 0 n14 ns209 0 -0.000633329329389
Gc7_210 0 n14 ns210 0 -0.000382151141602
Gc7_211 0 n14 ns211 0 2.67509916803e-05
Gc7_212 0 n14 ns212 0 6.31036374983e-05
Gc7_213 0 n14 ns213 0 -3.60786149866e-05
Gc7_214 0 n14 ns214 0 -0.000555524756047
Gc7_215 0 n14 ns215 0 0.000380665663411
Gc7_216 0 n14 ns216 0 -6.44542972484e-05
Gc7_217 0 n14 ns217 0 -0.000879196918108
Gc7_218 0 n14 ns218 0 0.000849630248681
Gc7_219 0 n14 ns219 0 -0.000647263366163
Gc7_220 0 n14 ns220 0 0.000158480206281
Gc7_221 0 n14 ns221 0 0.00112257812954
Gc7_222 0 n14 ns222 0 -0.000392131671173
Gc7_223 0 n14 ns223 0 -0.00160246997297
Gc7_224 0 n14 ns224 0 0.00223507662673
Gc7_225 0 n14 ns225 0 3.10546066302e-05
Gc7_226 0 n14 ns226 0 0.00114436418676
Gc7_227 0 n14 ns227 0 -0.00185056170339
Gc7_228 0 n14 ns228 0 -0.000488949148913
Gc7_229 0 n14 ns229 0 -0.000404274175992
Gc7_230 0 n14 ns230 0 -0.0015125962201
Gc7_231 0 n14 ns231 0 0.00127252031404
Gc7_232 0 n14 ns232 0 -0.000279632409414
Gc7_233 0 n14 ns233 0 0.00256104413606
Gc7_234 0 n14 ns234 0 0.000966686412341
Gc7_235 0 n14 ns235 0 0.000267621660262
Gc7_236 0 n14 ns236 0 0.00238224842807
Gc7_237 0 n14 ns237 0 -0.00090982119831
Gc7_238 0 n14 ns238 0 -0.00198197365466
Gc7_239 0 n14 ns239 0 -4.79262174988e-08
Gc7_240 0 n14 ns240 0 9.37937383707e-08
Gc7_241 0 n14 ns241 0 0.00329373638429
Gc7_242 0 n14 ns242 0 -0.000810754660031
Gc7_243 0 n14 ns243 0 0.00495834663093
Gc7_244 0 n14 ns244 0 -0.000142957313639
Gc7_245 0 n14 ns245 0 0.000119636693665
Gc7_246 0 n14 ns246 0 4.30569944165e-05
Gc7_247 0 n14 ns247 0 0.000598589197397
Gc7_248 0 n14 ns248 0 0.000542528425277
Gc7_249 0 n14 ns249 0 0.0157124693116
Gc7_250 0 n14 ns250 0 -2.78763698294e-05
Gc7_251 0 n14 ns251 0 8.81128514793e-05
Gc7_252 0 n14 ns252 0 2.96664303563e-06
Gc7_253 0 n14 ns253 0 4.04119121599e-05
Gc7_254 0 n14 ns254 0 0.00036112433164
Gc7_255 0 n14 ns255 0 -0.000651629134714
Gc7_256 0 n14 ns256 0 -0.000421925072148
Gc7_257 0 n14 ns257 0 -0.000221742440179
Gc7_258 0 n14 ns258 0 -0.000594362402817
Gc7_259 0 n14 ns259 0 -0.00164018375583
Gc7_260 0 n14 ns260 0 -0.000495472539511
Gc7_261 0 n14 ns261 0 0.000189038759372
Gc7_262 0 n14 ns262 0 -0.00218266557713
Gc7_263 0 n14 ns263 0 0.000691195906456
Gc7_264 0 n14 ns264 0 0.00115763509461
Gc7_265 0 n14 ns265 0 -0.000712623595424
Gc7_266 0 n14 ns266 0 5.81679494369e-05
Gc7_267 0 n14 ns267 0 0.000903633147994
Gc7_268 0 n14 ns268 0 0.00281275706506
Gc7_269 0 n14 ns269 0 -0.000461694273737
Gc7_270 0 n14 ns270 0 -0.000214550648703
Gc7_271 0 n14 ns271 0 -0.00133439577086
Gc7_272 0 n14 ns272 0 -0.0007684281554
Gc7_273 0 n14 ns273 0 4.05938246194e-05
Gc7_274 0 n14 ns274 0 -0.00412847401404
Gc7_275 0 n14 ns275 0 0.00191269431991
Gc7_276 0 n14 ns276 0 0.000131572839941
Gc7_277 0 n14 ns277 0 0.00198746821501
Gc7_278 0 n14 ns278 0 0.00184561555086
Gc7_279 0 n14 ns279 0 0.000163408899531
Gc7_280 0 n14 ns280 0 2.01794742121e-08
Gc7_281 0 n14 ns281 0 -4.97863994823e-08
Gc7_282 0 n14 ns282 0 -0.00347241035743
Gc7_283 0 n14 ns283 0 -0.00217948893272
Gc7_284 0 n14 ns284 0 0.0084054932548
Gc7_285 0 n14 ns285 0 6.43751747221e-05
Gc7_286 0 n14 ns286 0 -2.60697068899e-05
Gc7_287 0 n14 ns287 0 -5.1365335824e-05
Gc7_288 0 n14 ns288 0 0.000488806637333
Gc7_289 0 n14 ns289 0 -0.000121707611509
Gc7_290 0 n14 ns290 0 0.015317450714
Gc7_291 0 n14 ns291 0 -0.000217332661
Gc7_292 0 n14 ns292 0 -7.85933951057e-05
Gc7_293 0 n14 ns293 0 1.59813684049e-05
Gc7_294 0 n14 ns294 0 5.85903484073e-05
Gc7_295 0 n14 ns295 0 0.000338221237277
Gc7_296 0 n14 ns296 0 -0.000706994183079
Gc7_297 0 n14 ns297 0 -0.000167284208654
Gc7_298 0 n14 ns298 0 -0.000238337637349
Gc7_299 0 n14 ns299 0 -0.000678757203719
Gc7_300 0 n14 ns300 0 -0.00114138345187
Gc7_301 0 n14 ns301 0 -0.000615916180093
Gc7_302 0 n14 ns302 0 0.000224048269453
Gc7_303 0 n14 ns303 0 -0.00150197786711
Gc7_304 0 n14 ns304 0 0.000171852887982
Gc7_305 0 n14 ns305 0 0.000471733576548
Gc7_306 0 n14 ns306 0 0.000113592272498
Gc7_307 0 n14 ns307 0 5.17569338131e-05
Gc7_308 0 n14 ns308 0 0.00106988747082
Gc7_309 0 n14 ns309 0 0.00209471941082
Gc7_310 0 n14 ns310 0 -0.000163089218329
Gc7_311 0 n14 ns311 0 -0.000286382530906
Gc7_312 0 n14 ns312 0 -0.00155838061283
Gc7_313 0 n14 ns313 0 -0.000359361894428
Gc7_314 0 n14 ns314 0 -0.000236634379074
Gc7_315 0 n14 ns315 0 -0.00351601104325
Gc7_316 0 n14 ns316 0 0.00198367381193
Gc7_317 0 n14 ns317 0 0.000215104915465
Gc7_318 0 n14 ns318 0 0.00221112500189
Gc7_319 0 n14 ns319 0 0.00149095173986
Gc7_320 0 n14 ns320 0 0.000190979029339
Gc7_321 0 n14 ns321 0 -6.03049585401e-09
Gc7_322 0 n14 ns322 0 -2.81688239442e-08
Gc7_323 0 n14 ns323 0 -0.00300201769444
Gc7_324 0 n14 ns324 0 -0.00122235469562
Gc7_325 0 n14 ns325 0 0.0081106290634
Gc7_326 0 n14 ns326 0 3.96227595649e-05
Gc7_327 0 n14 ns327 0 -1.63064337427e-05
Gc7_328 0 n14 ns328 0 -2.98308191037e-05
Gd7_1 0 n14 ni1 0 0.000742357145657
Gd7_2 0 n14 ni2 0 0.000148706109866
Gd7_3 0 n14 ni3 0 8.5765221287e-05
Gd7_4 0 n14 ni4 0 -0.000649725280204
Gd7_5 0 n14 ni5 0 -0.000990163714005
Gd7_6 0 n14 ni6 0 -0.00323273116709
Gd7_7 0 n14 ni7 0 -0.00175453838447
Gd7_8 0 n14 ni8 0 -0.0020359667903
Gc8_1 0 n16 ns1 0 0.000129200492722
Gc8_2 0 n16 ns2 0 0.00143812142092
Gc8_3 0 n16 ns3 0 0.00311200566457
Gc8_4 0 n16 ns4 0 -4.26651022879e-05
Gc8_5 0 n16 ns5 0 0.000608576763813
Gc8_6 0 n16 ns6 0 5.73045125268e-05
Gc8_7 0 n16 ns7 0 -3.06422370313e-06
Gc8_8 0 n16 ns8 0 -0.000278368701934
Gc8_9 0 n16 ns9 0 -0.000249742809764
Gc8_10 0 n16 ns10 0 -0.000259921654222
Gc8_11 0 n16 ns11 0 -0.000295915875073
Gc8_12 0 n16 ns12 0 -0.00142228824903
Gc8_13 0 n16 ns13 0 -0.00118896360546
Gc8_14 0 n16 ns14 0 0.00078097788579
Gc8_15 0 n16 ns15 0 -0.000142897166768
Gc8_16 0 n16 ns16 0 0.00141261260893
Gc8_17 0 n16 ns17 0 -0.000602488639772
Gc8_18 0 n16 ns18 0 -0.000642241316229
Gc8_19 0 n16 ns19 0 0.00211782747929
Gc8_20 0 n16 ns20 0 2.07763610639e-05
Gc8_21 0 n16 ns21 0 0.00109960922353
Gc8_22 0 n16 ns22 0 0.00259324446524
Gc8_23 0 n16 ns23 0 -0.000337708078212
Gc8_24 0 n16 ns24 0 0.000216904095182
Gc8_25 0 n16 ns25 0 0.00151912860617
Gc8_26 0 n16 ns26 0 0.000279864239956
Gc8_27 0 n16 ns27 0 -0.000313665055588
Gc8_28 0 n16 ns28 0 0.0037593064145
Gc8_29 0 n16 ns29 0 0.00186962193254
Gc8_30 0 n16 ns30 0 9.81349109998e-05
Gc8_31 0 n16 ns31 0 0.0021226074323
Gc8_32 0 n16 ns32 0 2.76921307526e-05
Gc8_33 0 n16 ns33 0 0.000696196828794
Gc8_34 0 n16 ns34 0 -2.34484482692e-08
Gc8_35 0 n16 ns35 0 6.80245549808e-08
Gc8_36 0 n16 ns36 0 -0.00338289573071
Gc8_37 0 n16 ns37 0 -0.00298608910805
Gc8_38 0 n16 ns38 0 -0.00267421517599
Gc8_39 0 n16 ns39 0 5.16786547521e-05
Gc8_40 0 n16 ns40 0 -1.84698842705e-05
Gc8_41 0 n16 ns41 0 -4.67016325596e-05
Gc8_42 0 n16 ns42 0 -3.90347921127e-05
Gc8_43 0 n16 ns43 0 0.00122820110248
Gc8_44 0 n16 ns44 0 0.00405757662049
Gc8_45 0 n16 ns45 0 -0.000331319110322
Gc8_46 0 n16 ns46 0 0.000199835931002
Gc8_47 0 n16 ns47 0 7.20314688268e-05
Gc8_48 0 n16 ns48 0 4.78487974435e-05
Gc8_49 0 n16 ns49 0 -0.000206780543342
Gc8_50 0 n16 ns50 0 -0.000964601402025
Gc8_51 0 n16 ns51 0 3.27091376306e-05
Gc8_52 0 n16 ns52 0 -0.000281784322233
Gc8_53 0 n16 ns53 0 -0.000603584078124
Gc8_54 0 n16 ns54 0 -0.00127597772681
Gc8_55 0 n16 ns55 0 0.000890196988939
Gc8_56 0 n16 ns56 0 -0.00020027045641
Gc8_57 0 n16 ns57 0 0.000751157896736
Gc8_58 0 n16 ns58 0 -0.000378032692889
Gc8_59 0 n16 ns59 0 -0.00266064981004
Gc8_60 0 n16 ns60 0 0.00359040257482
Gc8_61 0 n16 ns61 0 -1.44229058465e-05
Gc8_62 0 n16 ns62 0 0.00126928959761
Gc8_63 0 n16 ns63 0 0.00211351744437
Gc8_64 0 n16 ns64 0 2.15912527364e-05
Gc8_65 0 n16 ns65 0 0.000206268127114
Gc8_66 0 n16 ns66 0 0.00174681852872
Gc8_67 0 n16 ns67 0 -7.60526970294e-05
Gc8_68 0 n16 ns68 0 -0.000355910963093
Gc8_69 0 n16 ns69 0 0.0028279679434
Gc8_70 0 n16 ns70 0 0.00370740088411
Gc8_71 0 n16 ns71 0 0.000169776070582
Gc8_72 0 n16 ns72 0 0.00221879856751
Gc8_73 0 n16 ns73 0 -0.000886144176239
Gc8_74 0 n16 ns74 0 0.00207803534601
Gc8_75 0 n16 ns75 0 4.1207240788e-09
Gc8_76 0 n16 ns76 0 7.61998023784e-08
Gc8_77 0 n16 ns77 0 -0.00354138123239
Gc8_78 0 n16 ns78 0 -0.00360545518404
Gc8_79 0 n16 ns79 0 -0.00370248532381
Gc8_80 0 n16 ns80 0 3.22615051287e-05
Gc8_81 0 n16 ns81 0 -3.456913642e-06
Gc8_82 0 n16 ns82 0 -4.03762060161e-05
Gc8_83 0 n16 ns83 0 0.000121286392708
Gc8_84 0 n16 ns84 0 -0.000325115880156
Gc8_85 0 n16 ns85 0 0.00361022282299
Gc8_86 0 n16 ns86 0 -0.000709323503895
Gc8_87 0 n16 ns87 0 -0.000121090536664
Gc8_88 0 n16 ns88 0 8.30519871877e-05
Gc8_89 0 n16 ns89 0 5.67515506652e-05
Gc8_90 0 n16 ns90 0 -0.000742883333356
Gc8_91 0 n16 ns91 0 -0.00133880476237
Gc8_92 0 n16 ns92 0 0.000734752676517
Gc8_93 0 n16 ns93 0 -0.00013859683999
Gc8_94 0 n16 ns94 0 -0.000368478487855
Gc8_95 0 n16 ns95 0 -0.00237739879019
Gc8_96 0 n16 ns96 0 0.00066350863894
Gc8_97 0 n16 ns97 0 -0.000118687879394
Gc8_98 0 n16 ns98 0 -0.00170537641468
Gc8_99 0 n16 ns99 0 0.000645644566496
Gc8_100 0 n16 ns100 0 -0.000828198394233
Gc8_101 0 n16 ns101 0 0.00900347839935
Gc8_102 0 n16 ns102 0 2.57016181956e-05
Gc8_103 0 n16 ns103 0 0.00111487059041
Gc8_104 0 n16 ns104 0 -0.00120183342605
Gc8_105 0 n16 ns105 0 0.000897357899241
Gc8_106 0 n16 ns106 0 0.000318710329749
Gc8_107 0 n16 ns107 0 0.00142657947752
Gc8_108 0 n16 ns108 0 -0.00180708105584
Gc8_109 0 n16 ns109 0 0.0020146586857
Gc8_110 0 n16 ns110 0 -5.0614671563e-06
Gc8_111 0 n16 ns111 0 0.0060181753889
Gc8_112 0 n16 ns112 0 -5.39835127984e-06
Gc8_113 0 n16 ns113 0 0.00149220851767
Gc8_114 0 n16 ns114 0 -0.00201818473726
Gc8_115 0 n16 ns115 0 0.00593758639381
Gc8_116 0 n16 ns116 0 7.21832478937e-08
Gc8_117 0 n16 ns117 0 5.68519688171e-08
Gc8_118 0 n16 ns118 0 -0.00172123100108
Gc8_119 0 n16 ns119 0 -0.00559848439106
Gc8_120 0 n16 ns120 0 -0.00387867833708
Gc8_121 0 n16 ns121 0 1.34895776389e-05
Gc8_122 0 n16 ns122 0 -5.7099212978e-06
Gc8_123 0 n16 ns123 0 -2.2013589657e-05
Gc8_124 0 n16 ns124 0 -0.000123287896978
Gc8_125 0 n16 ns125 0 0.00192106207098
Gc8_126 0 n16 ns126 0 0.0038659101706
Gc8_127 0 n16 ns127 0 0.000360311091882
Gc8_128 0 n16 ns128 0 -4.65304088619e-05
Gc8_129 0 n16 ns129 0 -2.58240952217e-05
Gc8_130 0 n16 ns130 0 1.28825774688e-05
Gc8_131 0 n16 ns131 0 0.000655698637605
Gc8_132 0 n16 ns132 0 -0.000387507587757
Gc8_133 0 n16 ns133 0 -1.36628721664e-05
Gc8_134 0 n16 ns134 0 0.000114932823678
Gc8_135 0 n16 ns135 0 -0.000918842193587
Gc8_136 0 n16 ns136 0 0.00344125534981
Gc8_137 0 n16 ns137 0 0.000910740816363
Gc8_138 0 n16 ns138 0 -0.000299543809142
Gc8_139 0 n16 ns139 0 -0.00081218386473
Gc8_140 0 n16 ns140 0 -0.000740701341117
Gc8_141 0 n16 ns141 0 -0.000872641298128
Gc8_142 0 n16 ns142 0 -0.00926493152717
Gc8_143 0 n16 ns143 0 6.59383213829e-05
Gc8_144 0 n16 ns144 0 0.00117699904685
Gc8_145 0 n16 ns145 0 -0.00189103901226
Gc8_146 0 n16 ns146 0 -0.000902379599053
Gc8_147 0 n16 ns147 0 8.66707654315e-05
Gc8_148 0 n16 ns148 0 0.00191075054754
Gc8_149 0 n16 ns149 0 0.00304938502866
Gc8_150 0 n16 ns150 0 -0.00353907930482
Gc8_151 0 n16 ns151 0 -0.00791964756614
Gc8_152 0 n16 ns152 0 -0.00408517847298
Gc8_153 0 n16 ns153 0 0.000494819841808
Gc8_154 0 n16 ns154 0 0.00403344754835
Gc8_155 0 n16 ns155 0 0.00430921956087
Gc8_156 0 n16 ns156 0 -0.0106919373642
Gc8_157 0 n16 ns157 0 -1.99111599014e-07
Gc8_158 0 n16 ns158 0 -1.66629034345e-08
Gc8_159 0 n16 ns159 0 0.00677979779801
Gc8_160 0 n16 ns160 0 0.00561902832113
Gc8_161 0 n16 ns161 0 -0.0117036921764
Gc8_162 0 n16 ns162 0 -0.000179422021423
Gc8_163 0 n16 ns163 0 0.000188302149884
Gc8_164 0 n16 ns164 0 7.34036559034e-05
Gc8_165 0 n16 ns165 0 0.00120623512833
Gc8_166 0 n16 ns166 0 -0.000701146913438
Gc8_167 0 n16 ns167 0 0.0110369257601
Gc8_168 0 n16 ns168 0 -0.000632745156639
Gc8_169 0 n16 ns169 0 -0.000362859435817
Gc8_170 0 n16 ns170 0 3.06015047543e-05
Gc8_171 0 n16 ns171 0 6.18126186158e-05
Gc8_172 0 n16 ns172 0 -2.33718816659e-05
Gc8_173 0 n16 ns173 0 -0.000573678465587
Gc8_174 0 n16 ns174 0 0.000396750960111
Gc8_175 0 n16 ns175 0 -6.80616080693e-05
Gc8_176 0 n16 ns176 0 -0.000931946011315
Gc8_177 0 n16 ns177 0 0.000809905707676
Gc8_178 0 n16 ns178 0 -0.000645100689635
Gc8_179 0 n16 ns179 0 0.000166082093062
Gc8_180 0 n16 ns180 0 0.00110724059572
Gc8_181 0 n16 ns181 0 -0.000415603768283
Gc8_182 0 n16 ns182 0 -0.00165175761237
Gc8_183 0 n16 ns183 0 0.00230241896974
Gc8_184 0 n16 ns184 0 3.26728097477e-05
Gc8_185 0 n16 ns185 0 0.00115016415955
Gc8_186 0 n16 ns186 0 -0.00183139606771
Gc8_187 0 n16 ns187 0 -0.000487526581443
Gc8_188 0 n16 ns188 0 -0.00041668255263
Gc8_189 0 n16 ns189 0 -0.0015153221409
Gc8_190 0 n16 ns190 0 0.00128474255547
Gc8_191 0 n16 ns191 0 -0.000313138416003
Gc8_192 0 n16 ns192 0 0.00252551352219
Gc8_193 0 n16 ns193 0 0.000991363493121
Gc8_194 0 n16 ns194 0 0.00027890322939
Gc8_195 0 n16 ns195 0 0.00237401752166
Gc8_196 0 n16 ns196 0 -0.000944119675588
Gc8_197 0 n16 ns197 0 -0.00196064310516
Gc8_198 0 n16 ns198 0 -4.70603070273e-08
Gc8_199 0 n16 ns199 0 9.60865683451e-08
Gc8_200 0 n16 ns200 0 0.00326683303911
Gc8_201 0 n16 ns201 0 -0.000783186052384
Gc8_202 0 n16 ns202 0 0.00493174628985
Gc8_203 0 n16 ns203 0 -0.000138234768639
Gc8_204 0 n16 ns204 0 0.000116360558207
Gc8_205 0 n16 ns205 0 4.25857047551e-05
Gc8_206 0 n16 ns206 0 0.000662129585673
Gc8_207 0 n16 ns207 0 -0.000369696478081
Gc8_208 0 n16 ns208 0 0.0097222537687
Gc8_209 0 n16 ns209 0 -0.000348095876792
Gc8_210 0 n16 ns210 0 -4.96526805405e-05
Gc8_211 0 n16 ns211 0 2.900097469e-05
Gc8_212 0 n16 ns212 0 3.73307760683e-05
Gc8_213 0 n16 ns213 0 -0.000179796542278
Gc8_214 0 n16 ns214 0 -0.000817420222906
Gc8_215 0 n16 ns215 0 0.000285743500178
Gc8_216 0 n16 ns216 0 -8.47263532499e-05
Gc8_217 0 n16 ns217 0 -0.000802924249545
Gc8_218 0 n16 ns218 0 0.000889451935992
Gc8_219 0 n16 ns219 0 -0.000758690769129
Gc8_220 0 n16 ns220 0 0.000225099189414
Gc8_221 0 n16 ns221 0 0.000803868087317
Gc8_222 0 n16 ns222 0 -0.000401908836134
Gc8_223 0 n16 ns223 0 -0.000281879679259
Gc8_224 0 n16 ns224 0 0.00217668148183
Gc8_225 0 n16 ns225 0 3.65721710915e-05
Gc8_226 0 n16 ns226 0 0.00128945199091
Gc8_227 0 n16 ns227 0 -0.00138694510942
Gc8_228 0 n16 ns228 0 -0.00012428559767
Gc8_229 0 n16 ns229 0 -0.000321892539492
Gc8_230 0 n16 ns230 0 -0.00175130119228
Gc8_231 0 n16 ns231 0 8.16695705633e-05
Gc8_232 0 n16 ns232 0 -0.000589309326038
Gc8_233 0 n16 ns233 0 0.00212975011276
Gc8_234 0 n16 ns234 0 0.00155856811034
Gc8_235 0 n16 ns235 0 9.55342063148e-05
Gc8_236 0 n16 ns236 0 0.00257077672737
Gc8_237 0 n16 ns237 0 0.00133664401823
Gc8_238 0 n16 ns238 0 -0.000111140876988
Gc8_239 0 n16 ns239 0 -4.74472647789e-09
Gc8_240 0 n16 ns240 0 2.92726298004e-08
Gc8_241 0 n16 ns241 0 0.00148830622455
Gc8_242 0 n16 ns242 0 -0.000218013176027
Gc8_243 0 n16 ns243 0 0.00614779658209
Gc8_244 0 n16 ns244 0 -3.38775194513e-05
Gc8_245 0 n16 ns245 0 2.56586959099e-05
Gc8_246 0 n16 ns246 0 1.74219738972e-05
Gc8_247 0 n16 ns247 0 0.000488806639915
Gc8_248 0 n16 ns248 0 -0.000121707612644
Gc8_249 0 n16 ns249 0 0.0153174507029
Gc8_250 0 n16 ns250 0 -0.000217332663822
Gc8_251 0 n16 ns251 0 -7.859340068e-05
Gc8_252 0 n16 ns252 0 1.59813686044e-05
Gc8_253 0 n16 ns253 0 5.85903479358e-05
Gc8_254 0 n16 ns254 0 0.00033822123697
Gc8_255 0 n16 ns255 0 -0.000706994179481
Gc8_256 0 n16 ns256 0 -0.000167284210302
Gc8_257 0 n16 ns257 0 -0.000238337635933
Gc8_258 0 n16 ns258 0 -0.000678757194408
Gc8_259 0 n16 ns259 0 -0.00114138344817
Gc8_260 0 n16 ns260 0 -0.000615916180777
Gc8_261 0 n16 ns261 0 0.000224048269081
Gc8_262 0 n16 ns262 0 -0.00150197786586
Gc8_263 0 n16 ns263 0 0.000171852890424
Gc8_264 0 n16 ns264 0 0.000471733589674
Gc8_265 0 n16 ns265 0 0.00011359226387
Gc8_266 0 n16 ns266 0 5.17569343385e-05
Gc8_267 0 n16 ns267 0 0.00106988747077
Gc8_268 0 n16 ns268 0 0.00209471940558
Gc8_269 0 n16 ns269 0 -0.000163089217068
Gc8_270 0 n16 ns270 0 -0.000286382529022
Gc8_271 0 n16 ns271 0 -0.00155838061251
Gc8_272 0 n16 ns272 0 -0.000359361898118
Gc8_273 0 n16 ns273 0 -0.000236634368391
Gc8_274 0 n16 ns274 0 -0.00351601104443
Gc8_275 0 n16 ns275 0 0.00198367379537
Gc8_276 0 n16 ns276 0 0.000215104918693
Gc8_277 0 n16 ns277 0 0.0022111250039
Gc8_278 0 n16 ns278 0 0.00149095173978
Gc8_279 0 n16 ns279 0 0.000190979022823
Gc8_280 0 n16 ns280 0 -6.03049667139e-09
Gc8_281 0 n16 ns281 0 -2.81688244429e-08
Gc8_282 0 n16 ns282 0 -0.00300201768687
Gc8_283 0 n16 ns283 0 -0.00122235471103
Gc8_284 0 n16 ns284 0 0.00811062907708
Gc8_285 0 n16 ns285 0 3.96227592679e-05
Gc8_286 0 n16 ns286 0 -1.63064348841e-05
Gc8_287 0 n16 ns287 0 -2.98308186104e-05
Gc8_288 0 n16 ns288 0 -0.000241957910758
Gc8_289 0 n16 ns289 0 0.000548523262111
Gc8_290 0 n16 ns290 0 0.0109615595421
Gc8_291 0 n16 ns291 0 0.000114025946576
Gc8_292 0 n16 ns292 0 0.000143975705159
Gc8_293 0 n16 ns293 0 2.55532398714e-05
Gc8_294 0 n16 ns294 0 3.18629475332e-05
Gc8_295 0 n16 ns295 0 0.000188719360747
Gc8_296 0 n16 ns296 0 -0.000706914148037
Gc8_297 0 n16 ns297 0 -4.51142008695e-05
Gc8_298 0 n16 ns298 0 -0.000160719513019
Gc8_299 0 n16 ns299 0 -0.000313222184088
Gc8_300 0 n16 ns300 0 -0.00107992318559
Gc8_301 0 n16 ns301 0 -0.000792786141141
Gc8_302 0 n16 ns302 0 0.000274228048978
Gc8_303 0 n16 ns303 0 -0.000983863269934
Gc8_304 0 n16 ns304 0 3.31285646803e-05
Gc8_305 0 n16 ns305 0 0.000286638095679
Gc8_306 0 n16 ns306 0 -0.000265559608915
Gc8_307 0 n16 ns307 0 8.3222522373e-05
Gc8_308 0 n16 ns308 0 0.00125775507331
Gc8_309 0 n16 ns309 0 0.00129117260479
Gc8_310 0 n16 ns310 0 -0.000126084837226
Gc8_311 0 n16 ns311 0 -0.000268697925147
Gc8_312 0 n16 ns312 0 -0.00178609040732
Gc8_313 0 n16 ns313 0 -8.33947560889e-05
Gc8_314 0 n16 ns314 0 0.000259058580985
Gc8_315 0 n16 ns315 0 -0.00229863058632
Gc8_316 0 n16 ns316 0 0.00135512088881
Gc8_317 0 n16 ns317 0 0.000200249091015
Gc8_318 0 n16 ns318 0 0.00286979844732
Gc8_319 0 n16 ns319 0 0.000947420921859
Gc8_320 0 n16 ns320 0 -0.000737236996886
Gc8_321 0 n16 ns321 0 -4.48292434693e-08
Gc8_322 0 n16 ns322 0 -1.10084906017e-07
Gc8_323 0 n16 ns323 0 -0.00148554190749
Gc8_324 0 n16 ns324 0 -0.00116550741197
Gc8_325 0 n16 ns325 0 0.00865060068263
Gc8_326 0 n16 ns326 0 7.53222285982e-05
Gc8_327 0 n16 ns327 0 -4.689984228e-05
Gc8_328 0 n16 ns328 0 -4.60318354747e-05
Gd8_1 0 n16 ni1 0 0.000148002284693
Gd8_2 0 n16 ni2 0 -6.68263984249e-05
Gd8_3 0 n16 ni3 0 -0.000653022949879
Gd8_4 0 n16 ni4 0 -0.000119260530555
Gd8_5 0 n16 ni5 0 -0.00325987892481
Gd8_6 0 n16 ni6 0 -0.00203460584088
Gd8_7 0 n16 ni7 0 -0.00203596678986
Gd8_8 0 n16 ni8 0 -0.000395144808391
.ends m4lines_HFSS_fws
