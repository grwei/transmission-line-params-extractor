* BEGIN ANSOFT HEADER
* node 1    1:trace_p_0_T1_A
* node 2    1:trace_n_0_T1_A
* node 3    1:trace_n_1_T1_A
* node 4    1:trace_p_1_T1_A
* node 5    Ground_A
* node 6    1:trace_p_0_T1_B
* node 7    1:trace_n_0_T1_B
* node 8    1:trace_n_1_T1_B
* node 9    1:trace_p_1_T1_B
* node 10   Ground_B
*  Project: 4lines
*   Design: 2-diff-pairs
*   Length: 5
*   Format: HSPICE
*  Creator: Ansoft HFSS
*     Date: Wed Jun 03 22:25:27 2020
* END ANSOFT HEADER

.subckt ckt_m4lines_HFSS_W 1 2 3 4 inref 5 6 7 8 outref length=5.08M

.model m4lines_HFSS_W_1 W MODELTYPE=table N=4 RMODEL=r_m4lines_HFSS_W_1
+ LMODEL=l_m4lines_HFSS_W_1 GMODEL=g_m4lines_HFSS_W_1 CMODEL=c_m4lines_HFSS_W_1

* Example usage:
W1 1 2 3 4 inref 5 6 7 8 outref N=4 L=length TABLEMODEL=m4lines_HFSS_W_1

.model r_m4lines_HFSS_W_1 sp N=4 SPACING=nonuniform VALTYPE=real
+ INTERPOLATION=spline
+ DATA = 700
+ 0           
+        6.906563104539061
+       0.6824161915317021
+        7.004584896377449
+       0.2837910405679777
+       0.9085696485041762
+        7.004887839056049
+       0.1145299239677343
+       0.2838404372629029
+       0.6766741287148066
+        6.856349044729821
+ 2e+08       
+        10.30113018179325
+        1.016369991615166
+        10.42632538041021
+       0.4018314087202817
+        1.334554596554753
+        10.41166364888455
+       0.1591891771844975
+       0.4037052692906891
+       0.9956869977619988
+        10.18231608077756
+ 3e+08       
+        12.64693105855384
+        1.143445082924333
+        12.80083132398006
+       0.4676939192679698
+         1.61106569253252
+         12.7762878231201
+       0.1753503940366344
+       0.4722341824890993
+        1.128844953370267
+        12.46352802132555
+ 4e+08       
+        14.63939197932881
+        1.258953351911071
+        14.82210135968447
+       0.5156127722746302
+        1.846192710895932
+          14.787841859159
+        0.181877090736275
+         0.52253867378994
+        1.249142618813348
+        14.39228693024461
+ 5e+08       
+        16.47200157222983
+        1.384934013041704
+        16.67790545488358
+       0.5602022126706039
+         2.06378850362835
+        16.63424818619715
+       0.1888717287836398
+       0.5693786520762407
+        1.377373107058749
+         16.1634982631831
+ 6e+08       
+        18.17011827891403
+        1.505648952327599
+        18.39373979737844
+       0.6034369240157705
+        2.264998191080702
+        18.34147658651015
+       0.1975974737755371
+       0.6147865607558634
+        1.498931333523312
+        17.80301996088844
+ 7e+08       
+        19.73880326064288
+        1.612446501113803
+        19.97721181134416
+       0.6444640535755874
+        2.449893571943583
+        19.91722839205754
+       0.2069202905547622
+       0.6578909896267338
+         1.60593246301257
+        19.31551094799766
+ 8e+08       
+        21.19426812974825
+        1.706646351512395
+        21.44648842603627
+       0.6826178836295976
+        2.620744225052114
+        21.37958398469257
+        0.215746200272815
+       0.6980109576400029
+        1.700104153249248
+        20.71677202728548
+ 9e+08       
+        22.56356240548607
+        1.795012715869257
+        22.82888586693532
+       0.7179645651863509
+        2.781310092291281
+        22.75579286350476
+       0.2235815349106163
+       0.7352228720687354
+        1.788452779992685
+        22.03380519838202
+ 1e+09       
+         23.8787626072638
+        1.885970198019283
+        24.15519908538059
+       0.7511468146685966
+         2.93583252969783
+        24.07668354204158
+       0.2304596376260809
+       0.7701990279719761
+        1.879579575967833
+        23.29895651296864
+ 1.1e+09     
+        25.23439621010591
+        1.953162989074464
+        25.40345676362819
+       0.6593952729784762
+        3.148419621962343
+         25.3161644270457
+       0.1461949917291049
+       0.6817102154408293
+        1.945272982535724
+        24.58812206945865
+ 1.2e+09     
+        26.46320012231223
+         2.02063262456289
+        26.52069742130246
+       0.5469368294826072
+        3.343671707458796
+        26.42528229185394
+      0.04862027002646629
+       0.5728135520858197
+         2.01145038260318
+        25.75327161632415
+ 1.3e+09     
+        27.58402771207589
+        2.088827533567694
+        27.54102337932396
+       0.4165514416650284
+         3.52381049901621
+        27.43818470785323
+     -0.06079701305075014
+       0.4462646860096726
+        2.078588998106512
+        26.81368916092968
+ 1.4e+09     
+        28.61624070571794
+        2.158152179055198
+        28.49205550505558
+       0.2712847251276949
+        3.690963973019537
+        28.38250013861808
+      -0.1803518493948287
+       0.3050782898185129
+        2.147100649617516
+        27.78892959902038
+ 1.5e+09     
+        29.57799063756573
+        2.228915191430468
+        29.39545077521032
+       0.1143696146813646
+        3.847015400556654
+        29.27986878256016
+      -0.3081714503715181
+       0.1524497328883166
+        2.217283710879249
+        28.69715789096771
+ 1.6e+09     
+        30.48533575901105
+         2.30130041959475
+        30.26771852544634
+     -0.05082360867929564
+        3.993573113791732
+        30.14676802371403
+      -0.4422685868574739
+    -0.008294854025377552
+        2.289298680834283
+        29.55431662562588
+ 1.7e+09     
+        31.35189918105111
+        2.375359832175536
+        31.12108935549303
+       -0.220824370874063
+        4.131994239483678
+        30.99538778192991
+      -0.5805828775022301
+      -0.1737355589058064
+        2.363165507904725
+        30.37382640655958
+ 1.8e+09     
+        32.18885545861282
+        2.451023078794199
+        31.96432736370161
+      -0.3920955000229395
+        4.263427821359292
+        31.83444729901646
+      -0.7210138125970227
+      -0.3403922114131879
+        2.438777035716231
+        31.16660625765551
+ 1.9e+09     
+        33.00510089456017
+        2.528117570375593
+        32.80344410963028
+      -0.5610695746838341
+        4.388860161391539
+        32.66991230350523
+      -0.8614485909170186
+      -0.5047603611920921
+        2.515922241345403
+        31.94127001602118
+ 2e+09       
+        33.80751369524279
+        2.606393606121469
+        33.64230485301013
+      -0.7241916713465375
+        4.509154407381867
+        33.50560345123922
+       -0.999787139501255
+      -0.6633533438789048
+        2.594313765874542
+        32.70440586118993
+ 2.1e+09     
+        34.60124573833206
+        2.685550343167307
+        34.48313199445361
+      -0.8779706353607907
+        4.625081204118231
+        34.34370120284491
+       -1.133966040680134
+      -0.8127524471172156
+        2.673615596315901
+        33.46088186354036
+ 2.2e+09     
+        35.39001164040534
+        2.765259735361215
+         35.3269163744954
+       -1.019039642511279
+        4.737339702947222
+        35.18515796543529
+       -1.261982512496776
+      -0.9496658529693009
+         2.75346813185731
+        34.21414433573324
+ 2.3e+09     
+        36.17635637239407
+        2.845186728976064
+        36.17374873534568
+       -1.144225525170154
+        4.846569513089414
+        36.03002993535437
+       -1.381919066278972
+       -1.070995781000009
+        2.833509041746479
+        34.96649123242305
+ 2.4e+09     
+        36.96189250444421
+        2.925004927692871
+        37.02308345176027
+        -1.25062502845818
+        4.953354866427934
+         36.8777408567727
+       -1.491968987447172
+       -1.173912008882052
+        2.913389241194899
+        35.71931254145159
+ 2.5e+09     
+        37.74750418522496
+        3.004407632571453
+        37.87394567126356
+       -1.335684853205919
+        5.058222653704513
+        37.72728892863883
+       -1.590462350787365
+       -1.255928716397642
+        2.992783989461196
+          36.473295485976
+ 2.6e+09     
+        38.53351850155399
+         3.08311465557189
+        38.72509177590008
+       -1.397281124408313
+        5.161636212456091
+        38.57740685278258
+       -1.675891899736072
+       -1.314980467318209
+        3.071399586978406
+        37.22859575427067
+ 2.7e+09     
+        39.31984681273151
+        3.160875630119862
+        39.57513181559552
+       -1.433792943493563
+        5.263986856331318
+        39.42668374477483
+       -1.746937812441757
+       -1.349492246964928
+        3.148976452460623
+        37.98497779218613
+ 2.8e+09     
+        40.10609959439464
+        3.237470725409665
+        40.42262136063299
+       -1.444164116870594
+        5.365585136117939
+        40.27365641849038
+       -1.802490174354668
+       -1.358437972514315
+        3.225289525147481
+        38.74192802156916
+ 2.9e+09     
+        40.89167863596374
+        3.312709731900933
+        41.26612910828744
+       -1.427947171098186
+        5.466653699851197
+        41.11687643459521
+        -1.84166790658272
+        -1.34138194104701
+        3.300146982762012
+        39.49874506551137
+ 3e+09       
+        41.67585035541597
+        3.386430439471702
+        42.10428555993581
+       -1.385324483905359
+        5.567323357548169
+        41.95495827493593
+       -1.863832980811929
+       -1.298498380740017
+        3.373388209084733
+        40.25461090964913
+ 3.1e+09     
+        42.45780368090296
+        3.458497093472171
+        42.93581715495404
+       -1.317102803005441
+        5.667633554239472
+         42.7866130634611
+       -1.868598986810249
+        -1.23056564003772
+        3.444881803119109
+        41.00864656219305
+ 3.2e+09     
+        43.23669550433806
+        3.528799508594032
+         43.7595694023579
+       -1.224679490643998
+        5.767537934838863
+        43.61067139579429
+       -1.855833485053278
+       -1.138933492036627
+        3.514524215365588
+        41.75995529512773
+ 3.3e+09     
+        44.01168621057353
+         3.59725317332586
+        44.57452179115793
+       -1.109981294193038
+        5.866915092933232
+        44.42609806546056
+       -1.825654027824317
+       -1.025464335818596
+        3.582239351937065
+        42.50765602482033
+ 3.4e+09     
+        44.78196728164778
+        3.663800421055237
+        45.37979659166803
+      -0.9753789773522212
+        5.965583999684664
+        45.23200079225182
+       -1.778418201571806
+      -0.8924514441676257
+        3.647979234813808
+        43.25090887283485
+ 3.5e+09     
+        45.54678251042557
+        3.728412511017551
+        46.17466309121643
+        -0.82358338858228
+        6.063323083968034
+        46.02763447772607
+       -1.714708458869945
+      -0.7425195034248713
+        3.711725578089788
+        43.98893447489696
+ 3.6e+09     
+        46.30544396165354
+        3.791092282546663
+        46.95853834662977
+      -0.6575301631230126
+        6.159891549045332
+        46.81240204360293
+       -1.635312805832286
+      -0.5785142126239258
+        3.773491963270625
+        44.72102820429551
+ 3.7e+09     
+        47.05734350864434
+        3.851876939280309
+        47.73098518555846
+      -0.4802610259606301
+        6.255051311590887
+        47.58585255496042
+       -1.541202548573005
+      -0.4033884459439694
+        3.833326190328933
+        45.44657016074333
+ 3.8e+09     
+        47.80196055536629
+        3.910840493192913
+          48.491707944954
+       -0.294809508378398
+         6.34858795180259
+        48.34767708742416
+       -1.433508270168335
+      -0.2200923611148129
+        3.891312352010152
+        46.16503155047057
+ 3.9e+09     
+        48.53886641963123
+        3.968095445163181
+        49.24054628551657
+      -0.1040978920580746
+        6.440329251528217
+         49.0977026530875
+       -1.313495030425659
+      -0.0314739279808478
+        3.947572220825245
+        46.87597794089004
+ 4e+09       
+        49.26772578715676
+        4.023793381855205
+        49.97746734691398
+       0.0891494351182244
+        6.530160226059773
+        49.83588443342689
+       -1.182537503966494
+       0.1598051520346946
+         4.00226563479839
+        47.57906979805205
+ 4.1e+09     
+        49.98829562712768
+         4.07812430409034
+        50.70255648748267
+       0.2824729995019888
+        6.618033963392385
+        50.56229655490868
+       -1.042095461210265
+        0.351334999400374
+        4.055589696629013
+        48.27406068698603
+ 4.2e+09     
+        50.70042196538204
+        4.131314644574092
+        51.41600686143131
+       0.4737244396323648
+        6.703978008191916
+        51.27712166017943
+      -0.8936897151151582
+       0.5410033346830772
+        4.107776737546093
+        48.96079351293947
+ 4.3e+09     
+        51.40403492232471
+        4.183624061279523
+        52.11810810666439
+       0.6610924811194593
+        6.788096411210989
+        51.98063955404108
+      -0.7388784543509379
+       0.7270219348495548
+        4.159091121025503
+        49.63919518711285
+ 4.4e+09     
+        52.09914242544348
+        4.235341192077501
+        52.80923443287153
+       0.8431106949397799
+        6.870567869819677
+        52.67321522385314
+      -0.5792337900234559
+       0.9079355686109936
+        4.209825058193634
+        50.30927010041344
+ 4.5e+09     
+        52.78582299338279
+        4.286778619091918
+        53.48983240381461
+        1.018649978949857
+         6.95164059249044
+        53.35528653993624
+      -0.4163183631772143
+        1.082616122675828
+        4.260293668875963
+        50.97109277545249
+ 4.6e+09     
+        53.46421795820315
+        4.338267317609341
+        54.16040869669686
+         1.18689916374194
+        7.031624628185568
+        54.02735193016781
+      -0.2516619773819797
+        1.250245100742717
+        4.310829549394542
+        51.62480003827157
+ 4.7e+09     
+        54.13452344723491
+        4.390150859233423
+        54.82151809595067
+         1.34733719734475
+        7.110882422679433
+        54.68995829570875
+     -0.08673840230708407
+        1.410287760825369
+        4.361777104969342
+        52.27058300905453
+ 4.8e+09     
+        54.79698239090284
+        4.442779610508947
+        55.47375194226283
+        1.499700108192199
+        7.189818317786447
+        55.34368939582529
+      0.07705730018598445
+         1.56246194363732
+          4.4134868785468
+        52.90867915970404
+ 4.9e+09     
+        55.45187676390717
+         4.49650512546706
+        56.11772721471809
+        1.643945492103074
+        7.268867618719126
+        55.98915488413235
+       0.2384303869855979
+        1.706704236479956
+        4.466310067702525
+        53.53936463103001
+ 5e+09       
+        56.09952020972347
+        4.551674881889117
+        56.75407637911045
+        1.780216718252641
+        7.348485740476222
+        56.62698013124619
+       0.3962063035116419
+        1.843135608561677
+         4.52059337498957
+        54.16294694843417
+ 5.1e+09     
+        56.74025114674738
+        4.608627463232895
+        57.38343809242001
+        1.908808483122076
+        7.429137823553472
+        57.25779692370116
+       0.5493480711506598
+        1.972028122965897
+        4.576674291274063
+        54.77975822642067
+ 5.2e+09     
+        57.37442641128784
+        4.667688245782703
+        58.00644881491762
+        2.030134818035732
+        7.511289094920525
+        57.88223508886706
+       0.6969704734299453
+        2.093773833809825
+        4.634876870766169
+        55.39014891161275
+ 5.3e+09     
+        58.00241545918104
+        4.729165616231512
+        58.62373534873527
+        2.144700209599714
+         7.59539614991247
+        58.50091506197121
+       0.8383504269113118
+        2.208856548987831
+        4.695508023201953
+         55.9944820824002
+ 5.4e+09     
+        58.62459512395108
+        4.793347719441153
+        59.23590829570482
+        2.253074138003138
+        7.681899248261838
+        59.11444138470807
+       0.9729330964027905
+        2.317826795191567
+        4.758854323870316
+        56.59312830082704
+ 5.5e+09     
+        59.24134491410202
+        4.860499719081026
+        59.84355640753864
+        2.355869076016511
+        7.771215653724818
+        59.72339710501554
+        1.100333534495925
+        2.421280064458819
+        4.825179325509017
+        57.18646099791028
+ 5.6e+09     
+        59.85304282373424
+        4.930861543958017
+        60.44724178747165
+        2.453721812525617
+        7.863734000432979
+        60.32833903371738
+        1.220333866574083
+        2.519838242845152
+         4.89472134634806
+        57.77485236574953
+ 5.7e+09     
+        60.46006162736956
+        5.004646088431924
+        61.04749589334734
+        2.547277854382907
+        7.959809637859202
+        60.92979380487113
+        1.332876278121296
+         2.61413400928693
+        4.967691704144528
+        58.35866972683655
+ 5.8e+09     
+        61.06276562989861
+        5.082037834641732
+           61.64481628691
+        2.637178603536839
+        8.059760887299255
+        61.52825468180288
+        1.438052268519506
+        2.704797931765427
+        5.044273365263104
+        58.93827235119232
+ 5.9e+09     
+        61.66150784440074
+        5.163191865779935
+        62.23966407179014
+        2.724050987730438
+        8.163866133186897
+        62.12417904897848
+        1.536088797444306
+        2.792447964404713
+         5.12461997920817
+        59.51400869390536
+ 6e+09       
+         62.2566275730743
+        5.248233242101479
+        62.83246196258457
+         2.80849922955024
+        8.272361669783024
+        62.71798653017948
+        1.627332056440023
+        2.877681050730939
+        5.208855271277552
+        60.08621402817482
+ 6.1e+09     
+        62.84844836879067
+        5.337256713851726
+        63.42359292877376
+        2.891098459930848
+        8.385440225614468
+        63.31005767523818
+          1.7122296464214
+        2.961066555079492
+        5.297072768330548
+        60.65520845128823
+ 6.2e+09     
+        63.43727635646332
+        5.430326747305504
+        64.01339935953422
+        2.972389910765693
+        8.503250092730568
+        63.90073316025664
+        1.791311935203386
+         3.04314126866899
+        5.389335834513971
+        61.22129524266624
+ 6.3e+09     
+        64.02339889427012
+        5.527477841385385
+        64.60218269830716
+        3.052877451880484
+        8.625894794053407
+        64.49031344939998
+        1.865173315968903
+        3.124405764074452
+        5.485677994924254
+        61.78475955398833
+ 6.4e+09     
+        64.60708355486344
+        5.628715112859169
+        65.19020349903387
+        3.133025267125158
+        8.753433228859265
+        65.07905886969348
+        1.934453999099894
+         3.20532189860561
+        5.586103525614651
+        62.34586741157024
+ 6.5e+09     
+        65.18857740620162
+        5.734015128027647
+        65.77768185903815
+        3.213256491130001
+        8.885880243091631
+        65.66719005357949
+        1.999822858399566
+        3.286311291707227
+        5.690588288167354
+        62.90486501069999
+ 6.6e+09     
+        65.76810657076047
+        5.843326958310633
+        66.36479818650191
+         3.29395265167414
+        9.023207577347909
+        66.25488870719124
+        2.061961730425951
+        3.367754623281609
+        5.799080786492144
+        63.46197828084793
+ 6.7e+09     
+        66.34587604091162
+        5.956573436445303
+        66.95169426327817
+        3.375453782724173
+         9.16534515077935
+        66.84229866526819
+        2.121551442896806
+        3.449991618735401
+        5.911503422762128
+        64.01741269974198
+ 6.8e+09     
+        66.92206972733892
+        6.073652589335466
+        67.53847456636944
+        3.458059090356322
+        9.312182643699282
+        67.42952719639486
+        2.179259733174163
+        3.533321602849558
+         6.02775392868927
+         64.5713533334612
+ 6.9e+09     
+        67.49685071671759
+        6.194439223084251
+        68.12520781379371
+        3.542028068482243
+         9.46357134540313
+        68.01664652475307
+        2.235731116469437
+        3.618004518711144
+        6.147706947811631
+        65.12396507911257
+ 7e+09       
+        68.07036171456087
+        6.318786635528872
+        68.71192870271911
+        3.627581974060839
+        9.619326236617484
+        68.60369553685125
+        2.291578679042134
+        3.704262320342204
+        6.271215744233668
+        65.67539308639957
+ 7.1e+09     
+        68.64272564922702
+        6.446528431728077
+        69.29863980977339
+         3.71490558272468
+        9.779228278217611
+        69.19068164380326
+        2.347377705600044
+        3.792280658706304
+        6.398114013382971
+        66.22576333452828
+ 7.2e+09     
+        69.21404641354935
+        6.577480418341556
+        69.88531362527564
+        3.804149155791216
+        9.943026879476404
+        69.77758277162167
+        2.403661002038801
+        3.882210790724437
+        6.528217770828435
+        66.77518334141219
+ 7.3e+09     
+        69.78440972138773
+        6.711442553677697
+        70.47189469487788
+        3.895430558721928
+        10.11044252027321
+        70.36434945379135
+        2.460915743084835
+        3.974171650019243
+        6.661327296041604
+        67.32374298301268
+ 7.4e+09     
+        70.35388405753692
+        6.848200931319363
+        71.05830184373873
+        3.988837479351773
+        10.28116950248563
+        70.95090700204095
+        2.519581657111241
+        4.068252026409978
+         6.79722910910783
+         67.8715154018078
+ 7.5e+09     
+        70.92252170080896
+        6.987529776620136
+        71.64443045992537
+        4.084429701760936
+        10.45487880634927
+        71.53715773282438
+         2.58005035482102
+        4.164512808811732
+        6.935697959780478
+        68.41855798479571
+ 7.6e+09     
+        71.49035980165159
+        7.129193436921554
+        72.23015481524921
+        4.182241398505878
+        10.63122102796545
+        72.12298322852945
+        2.642665612020356
+        4.262989253139562
+        7.076498809828461
+        68.96491339297573
+ 7.7e+09     
+        72.05742149731019
+        7.272948348040332
+        72.81533040323229
+        4.282283410140281
+        10.80982937447416
+        72.70824661391704
+        2.707724426875765
+        4.363693243134266
+        7.219388791315939
+        69.51061062591683
+ 7.8e+09     
+        72.62371704924809
+         7.41854496132487
+        73.39979627535543
+        4.384545486510778
+        10.99032269374268
+        73.29279482971519
+        2.775478686693892
+        4.466615517701296
+         7.36411912521177
+        70.05566610670252
+ 7.9e+09     
+        73.18924498921301
+        7.565729617368286
+        73.98337735818751
+        4.488998469259622
+         11.1723085158145
+        73.87646088672322
+        2.846137296547624
+         4.57172784339952
+        7.510436986502843
+        70.60008477422232
+ 8e+09       
+        73.75399326199809
+        7.714246354230073
+        74.56588673543737
+        4.595596399308209
+        11.35538608385582
+        74.45906608516275
+        2.919868640547862
+        4.678985115166403
+        7.658087303749084
+        71.14386117140393
+ 8.1e+09     
+        74.31794035451091
+        7.863838639737295
+        75.14712788038878
+        4.704278536878035
+        11.53914935296835
+         75.0404221854031
+        2.996803265107634
+        4.788327372235653
+        7.806814482731127
+        71.68698051952923
+ 8.2e+09     
+        74.88105640224697
+         8.01425101908549
+        75.72689682560873
+         4.81497128484467
+        11.72318993601625
+        75.62033351755051
+        3.077036691369254
+        4.899681719539435
+        7.956364045488229
+        72.22941977022829
+ 8.3e+09     
+        75.44330426563657
+        8.165230670524519
+        76.30498425822618
+        4.927590008985948
+        11.90709997656074
+        76.19859901874426
+        3.160632280528591
+        5.012964147713809
+        8.106484177597096
+        72.77114862808797
+ 8.4e+09     
+        76.00464056999732
+        8.316528863380109
+         76.8811775304676
+        5.042040751002745
+        12.09047493010791
+        76.77501418832784
+         3.24762409077713
+        5.128081247218457
+         8.25692717800689
+        73.31213053803111
+ 8.5e+09     
+        76.56501670397159
+        8.467902314024597
+        77.45526257650975
+        5.158221832111155
+        12.27291623614379
+        77.34937295238029
+        3.338019677829982
+        5.244931814061527
+        8.407450807099796
+        73.85232363274359
+ 8.6e+09     
+        77.12437977235852
+        8.619114436669205
+        78.02702572804822
+         5.27602534658484
+        12.45403386484758
+        77.92146943035615
+         3.43180280249099
+        5.363408346251457
+        8.557819529896708
+        74.39168163640731
+ 8.7e+09     
+        77.68267350018496
+        8.769936486999127
+        78.59625542229159
+        5.395338545907473
+        12.63344872392152
+        78.49109959783368
+        3.528936018479454
+        5.483398431414656
+        8.707805652471258
+        74.93015472189202
+ 8.8e+09     
+        78.23983908567416
+        8.920148597722875
+        79.16274379734683
+        5.516045115213791
+        12.81079491263147
+         79.0580628405677
+        3.629363121916956
+        5.604786027092562
+        8.857190350678501
+        75.46769031934687
+ 8.9e+09     
+        78.79581600050452
+        9.069540706045554
+        79.72628817117675
+        5.638026344502647
+        12.98572181189125
+        79.62216339618797
+        3.733011450592613
+        5.727452636044832
+        9.005764591234634
+        76.00423387480332
+ 9e+09       
+        79.35054273639791
+        9.217913373930834
+        80.28669240146702
+        5.761162197731713
+        13.15789600102755
+        80.18321168099015
+        3.839794026561771
+        5.851278379562588
+        9.153329946034258
+        76.53972955802729
+ 9.1e+09     
+        79.90395749761467
+        9.365078502759864
+        80.84376812483124
+        5.885332283369802
+        13.32700299369518
+        80.74102550029616
+        3.949611539937878
+        5.976142972270436
+        9.299699301327687
+        77.07412091935501
+ 9.2e+09     
+        80.45599883945025
+          9.5108599446681
+        81.39733587480764
+        6.010416730333379
+        13.49274878725419
+        81.29543114183765
+        4.062354175089631
+        6.101926602275222
+        9.444697464048357
+        77.60735149571788
+ 9.3e+09     
+        81.00660625321798
+        9.655094013413571
+        81.94722607905587
+        6.136296973484192
+        13.65486122174987
+        81.84626435252413
+        4.177903282988984
+        6.228510720772228
+        9.588161668146215
+        78.13936536642808
+ 9.4e+09     
+        81.55572069858347
+        9.797629898134426
+        82.49327993703548
+        6.262856453019245
+        13.81309114641801
+        82.39337119978596
+        4.296132905320679
+        6.355778745412136
+        9.729941984286103
+         78.6701076596423
+ 9.5e+09     
+        82.10328508440983
+        9.938329983777493
+        83.03535018025374
+        6.389981232193721
+         13.9672133933645
+         82.9366088194503
+        4.416911157271768
+        6.483616681826128
+        9.869901636682739
+        79.19952501067833
+ 9.6e+09     
+        82.64924469953644
+        10.07707008233487
+        83.57330171787937
+        6.517560537853092
+        14.11702755970774
+        83.47584605279143
+         4.54010147678441
+         6.61191366777215
+        10.00791723120293
+        79.72756597359975
+ 9.7e+09     
+        83.19354759512345
+        10.21373957931698
+        84.10701217117315
+         6.64548722826687
+        14.26235860101994
+        84.01096397601174
+        4.665563748562646
+         6.74056244437292
+        10.14387889914845
+        80.25418138766837
+ 9.8e+09     
+        83.73614492036984
+        10.34824150011937
+        84.63637230072899
+        6.773658192704313
+         14.4030572403298
+        84.54185632593909
+         4.79315531135112
+        6.869459758888739
+        10.27769036136089
+        80.77932470041311
+ 9.9e+09     
+        84.27699121355737
+        10.48049250111602
+        85.16128633101846
+        6.901974687161552
+        14.53900019826523
+        85.06842982620633
+        4.922731857020121
+        6.998506703420581
+        10.40926891746241
+        81.30295224918703
+ 1e+10       
+        84.81604465047202
+        10.61042279043266
+        85.68167217712174
+        7.030342610544302
+        14.67009025108539
+        85.59060441854601
+        5.054148229843528
+        7.127608993862992
+        10.53854536516506
+         81.8250235031658
+ 1.01e+10    
+        85.35326725234566
+        10.73797598342876
+        86.19746157886698
+        7.158672725537701
+        14.79625612439672
+        86.10831340418054
+        5.187259134089564
+        7.256677193323336
+        10.66546385465629
+        82.34550126782048
+ 1.02e+10    
+        85.88862505550701
+        10.86310889795184
+        86.70860014786366
+        7.286880828259504
+        14.91745223124517
+        86.62150350052161
+         5.32191975769913
+        7.385626884135728
+        10.78998168309922
+         82.8643518539243
+ 1.03e+10    
+         86.4220882449783
+        10.98579129441547
+        87.21504733309898
+        7.414887870701227
+        15.03365826403806
+        87.13013481860192
+        5.457986319420447
+        7.514378792458704
+        10.91206903427745
+        83.38154521318189
+ 1.04e+10    
+        86.95363125425386
+        11.10600556571707
+        87.71677631091119
+         7.54262003980212
+        15.14487865036899
+        87.63418076678191
+        5.595316546331411
+        7.642858869328222
+        11.03170866837303
+        83.89705504258433
+ 1.05e+10    
+        87.48323283351054
+        11.22374638193162
+        88.21377380521461
+        7.670008796887885
+        15.25114188330321
+        88.13362788636145
+        5.733770088230568
+        7.770998331900492
+         11.1488955667927
+         84.4108588595616
+ 1.06e+10    
+        88.01087608846734
+        11.33902029462217
+         88.7060398438813
+        7.796990881047355
+         15.3524997370367
+        88.62847562474627
+        5.873208874916378
+        7.898733668472889
+        11.26363653685765
+        84.92293805001117
+ 1.07e+10    
+        88.53654849209954
+        11.45184530548019
+        89.19358745714867
+        7.923508279887803
+         15.4490263790696
+        89.11873605180351
+        6.013497421927616
+        8.026006610731017
+        11.37594978104534
+        85.43327789121879
+ 1.08e+10    
+        89.06024187135628
+        11.56225040386386
+        89.67644232385568
+        8.049508170941731
+        15.54081739014938
+        89.60443352497606
+        6.154503089875818
+        8.152764076512073
+        11.48586443533013
+        85.94186755166612
+ 1.09e+10    
+        89.58195237098867
+        11.67027507763877
+        90.15464237119184
+        8.174942836869025
+        15.62798870324347
+        90.08560430862846
+        6.296096302085266
+        8.278958086231714
+        11.59342008100327
+        86.44870006965562
+ 1.1e+10     
+        90.10168039653584
+         11.7759688015479
+         90.6282373335066
+        8.299769557416949
+         15.7106754727051
+        90.56229615296365
+        6.438150724852967
+        8.404545655959659
+        11.69866623418024
+        86.95377231263296
+ 1.11e+10    
+        90.61943053844513
+        11.87939050714636
+        91.09728827554507
+        8.423950480976792
+        15.78903088461334
+        91.03456783768848
+        6.580543414269663
+        8.529488669974171
+        11.80166181700838
+         87.4570849190174
+ 1.12e+10    
+        91.13521147924244
+        11.98060803813748
+        91.56186708527669
+        8.547452478390394
+        15.86322491900223
+        91.50248868542324
+         6.72315493318991
+        8.653753735484244
+        11.90247461439461
+        87.95864222428499
+ 1.13e+10    
+        91.64903588558229
+        12.07969759474111
+        92.02205594127129
+        8.670246981537023
+        15.93344307435853
+        91.96613804964146
+        6.865869441613684
+        8.777312022030882
+        12.00118071986352
+        88.45845217297889
+ 1.14e+10    
+         92.1609202869307
+        12.17674317050935
+        92.47794675932353
+        8.792309809048344
+         15.9998850643708
+        92.42560478170496
+        7.008574763439726
+        8.900139087949359
+        12.09786397394799
+        88.95652621824253
+ 1.15e+10    
+        92.67088494255933
+        12.27183598479485
+        92.92964062279191
+        8.913620981374427
+        16.06276349646276
+          92.880986681328
+        7.151162432271456
+        9.022214696103376
+        12.19261539829944
+        89.45287921039944
+ 1.16e+10    
+        93.17895369843198
+        12.36507391385568
+        93.37724720085151
+        9.034164527257277
+        16.12230254115374
+        93.33238993454674
+        7.293527718702199
+        9.143522620971034
+        12.28553262849018
+        89.94752927602194
+ 1.17e+10    
+        93.68515383549588
+        12.45656092337193
+        93.82088415858796
+        9.153928283538562
+        16.17873660076073
+        93.77992854303798
+        7.435569641270814
+        9.264050449000592
+        12.37671934826615
+        90.44049768885266
+ 1.18e+10    
+        94.18951591078678
+        12.54640650492549
+        94.26067656260329
+        9.272903690067091
+        16.23230898540188
+        94.22372374835209
+        7.577190963063095
+        9.383789374023003
+        12.46628472779598
+        90.93180873386851
+ 1.19e+10    
+        94.69207359269011
+        12.63472511879323
+        94.69675628551583
+        9.391085581351572
+        16.28327060369078
+         94.6639034543812
+        7.718298175740737
+        9.502733989357653
+         12.5543428682504
+        91.42148956569351
+ 1.2e+10     
+        95.19286349160136
+        12.72163564519117
+        95.12926141248461
+        9.508471976460774
+        16.33187867492331
+        95.10060165112813
+          7.8588014726023
+        9.620882078131306
+        12.64101225484334
+        91.90957006248948
+ 1.21e+10    
+        95.69192498714895
+         12.8072608459064
+        95.55833565260367
+        9.625063868540286
+        16.37839546896592
+        95.53395784257451
+        7.998614712114265
+        9.738234403174053
+        12.72641522026359
+        92.39608267638661
+ 1.22e+10    
+        96.18930005307075
+        12.89172683806041
+        95.98412775776617
+        9.740865015198644
+        16.42308707946232
+        95.96411648120528
+        8.137655373209785
+          9.8547944977519
+         12.8106774202304
+        92.88106228142708
+ 1.23e+10    
+        96.68503308073805
+        12.97516258155446
+        96.40679095133382
+        9.855881730883739
+        16.46622223538624
+        96.39122641150236
+         8.27584450351276
+        9.970568458266111
+        12.89392732272154
+        93.36454601993276
+ 1.24e+10    
+         97.1791707022543
+        13.05769938156813
+        96.82648236869917
+        9.970122682264252
+        16.50807115538428
+        96.81544032447425
+         8.41310666152976
+        10.08556473992691
+        12.97629571223558
+        93.84657314813776
+ 1.25e+10    
+        97.67176161397933
+        13.13947040730819
+        97.24336251159733
+        10.08359868751695
+        16.54890444879107
+        97.23691422506943
+        8.549369853739673
+        10.19979395631106
+        13.05791521028296
+        94.32718488184537
+ 1.26e+10    
+        98.16285640125054
+        13.22061022803556
+        97.65759471778905
+        10.19632252030877
+        16.58899206663911
+         97.6558069140923
+        8.684565467412311
+        10.31326868359342
+        13.13891981312963
+        94.80642424282564
+ 1.27e+10    
+        98.65250736500883
+        13.30125436724366
+         98.0693446475194
+        10.30830871917496
+        16.62860230545796
+        98.07227948603085
+        8.818628199900694
+        10.42600327015558
+        13.21944444766191
+        95.28433590657995
+ 1.28e+10    
+        99.14076835096149
+         13.3815388757089
+        98.47877978795357
+        10.41957340288724
+        16.66800086614279
+        98.48649484400983
+        8.951495985066565
+        10.53801365217049
+        13.29962454609149
+         95.7609660520598
+ 1.29e+10    
+        99.62769458185923
+        13.46159992399386
+        98.88606897658902
+        10.53013409232746
+        16.70744996968339
+        98.89861723288747
+        9.083109917429592
+        10.64931717566529
+        13.37959564007972
+        96.23636221385732
+ 1.3e+10     
+        100.1133424933896
+        13.54157341485129
+        99.29138194446882
+        10.64000953928674
+        16.74720753108156
+        99.30881179133105
+        9.213414174563628
+        10.75993242550873
+        13.45949297472516
+        96.71057313733257
+ 1.31e+10    
+         100.597769574148
+        13.62159461585197
+        99.69488887983421
+        10.74921956254239
+        16.78752639234686
+        99.71724412355182
+         9.34235593820341
+        10.86987906165248
+        13.53945114273852
+         97.1836486370897
+ 1.32e+10    
+        101.0810342100701
+        13.70179781244528
+        100.0967600127103
+        10.85778489148657
+        16.82865361504938
+        100.1240798912057
+        9.469885314472901
+        10.97917766291147
+        13.61960373901139
+        97.65563945916607
+ 1.33e+10    
+        101.5631955336756
+          13.782315981552
+        100.4971652207575
+        10.96572701750849
+         16.8708298325269
+        100.5294844258353
+        9.595955253597509
+        11.08784957848809
+        13.70008303567838
+        98.12659714724768
+ 1.34e+10    
+        102.0443132784151
+        13.86328048569141
+        100.8962736565887
+        11.07306805327513
+        16.91428866148836
+        100.9336223620789
+         9.72052146941969
+        11.19591678737982
+        13.78101967767395
+        98.59657391318461
+ 1.35e+10    
+        102.5244476383607
+        13.94482078755308
+        101.2942533966273
+        11.17983059999697
+        16.95925617242906
+        101.3366572917622
+        9.843542358996862
+        11.30340176575865
+        13.86254239869378
+        99.06562251203258
+ 1.36e+10    
+        103.0036591334499
+        14.02706418483953
+        101.6912711114605
+        11.28603762270463
+        17.00595041797692
+        101.7387514388642
+        9.964978922528216
+        11.41032736234976
+        13.94477775738817
+        99.53379612181406
+ 1.37e+10    
+         103.482008480442
+        14.11013556513218
+        102.0874917575457
+        11.39171233352247
+        17.05458101801848
+        102.1400653552475
+        10.08479468382289
+        11.51671668179793
+        14.02784989353838
+        100.0011482281516
+ 1.38e+10    
+        103.9595564697041
+        14.19415718046236
+        102.4830782900262
+        11.49687808287897
+        17.10534880020981
+        102.5407576369545
+        10.20295561149436
+        11.62259297595136
+         14.1118803038994
+        100.4677325138927
+ 1.39e+10    
+        104.4363638479274
+        14.27924844120871
+         102.878191396331
+        11.60155825854459
+        17.15844549426505
+        102.9409846607783
+        10.31943004104145
+        11.72797954297037
+         14.1969876373301
+        100.9336027538169
+ 1.4e+10     
+        104.9124912068174
+        14.36552572888744
+        103.2729892501619
+        11.70577619237259
+        17.21405347822497
+        103.3409003407494
+        10.43418859795171
+        11.83289963411813
+        14.28328750877824
+        101.3988127144836
+ 1.41e+10    
+         105.387998877794
+        14.45310222735386
+        103.6676272853955
+        11.80955507456032
+        17.27234557474259
+        103.7406559041092
+        10.54720412194442
+        11.93737636806592
+        14.37089233163854
+        101.8634160592533
+ 1.42e+10    
+        105.8629468326932
+         14.5420877718899
+        104.0622579893859
+        11.91291787524942
+        17.33348489528912
+        104.1403996862852
+        10.65845159245012
+        12.04143265251998
+        14.45991116796054
+        102.3274662584914
+ 1.43e+10    
+        106.3373945904463
+        14.63258871561832
+        104.4570307150844
+        12.01588727323068
+        17.39762473006038
+        104.5402769443294
+        10.76790805540932
+        12.14509111294767
+        14.55044959594596
+        102.7910165049408
+ 1.44e+10    
+        106.8114011296904
+        14.72470781265046
+        104.8520915113707
+        12.11848559152631
+        17.46490848127772
+        104.9404296882441
+        10.87555255145583
+        12.24837402816063
+        14.64260959414417
+        103.2541196342267
+ 1.45e+10    
+        107.2850248072367
+        14.81854411735121
+        105.2475829709446
+        12.22073473958363
+        17.53546963750053
+        105.3409965295789
+        10.98136604554029
+        12.35130327250394
+        14.73648944173078
+         103.716828050447
+ 1.46e+10    
+        107.7583232823084
+        14.91419289908153
+        105.6436440950949
+        12.32265616181145
+        17.60943178651456
+        105.7421125466566
+        11.08533135803431
+        12.45390026437045
+        14.83218363422793
+        104.1791936567688
+ 1.47e+10    
+        108.2313534464493
+        15.01174557176519
+        106.0404101746583
+        12.42427079217774
+        17.68690866433202
+        106.1439091657575
+        11.18743309734846
+        12.55618592076723
+        14.92978281401633
+        104.6412677909569
+ 1.48e+10    
+        108.7041713589767
+        15.11128963761036
+        106.4380126864424
+        12.52559901457406
+        17.76800423781528
+        106.5465140575857
+        11.28765759408633
+        12.65818061763606
+        15.02937371496975
+        105.1031011657332
+ 1.49e+10    
+        109.1768321878532
+        15.21290864431301
+        106.8365792043958
+        12.62666062865156
+        17.85281281844033
+        106.9500510483116
+        11.38599283674882
+         12.7599041556333
+        15.13103912053741
+        105.5647438138542
+ 1.5e+10     
+         109.649390155826
+        15.31668215505922
+        107.2362333247876
+        12.72747482082991
+          17.941419204731
+        107.3546400444969
+        11.48242840899683
+         12.8613757310664
+        15.23485783459709
+         106.026245037793
+ 1.51e+10    
+        110.1218984916962
+        15.42268573064917
+        107.6370946046705
+        12.82806014017211
+        18.03389885091817
+         107.760396971187
+        11.57695542847359
+        12.96261391168953
+        15.34090466439499
+        106.4876533638972
+ 1.52e+10    
+        110.5944093865378
+        15.53099092305822
+        108.0392785128906
+        12.92843447882231
+          18.130318059423
+        108.1674337224708
+        11.66956648718134
+         13.0636366170503
+        15.44925041489722
+        106.9490165008833
+ 1.53e+10    
+        111.0669739547132
+        15.64166527976392
+        108.4428963929234
+         13.0286150567136
+        18.23073419481069
+        108.5758581238046
+        11.76025559340439
+         13.1644611030888
+        15.55996189387452
+        107.4103813025311
+ 1.54e+10    
+        111.5396421995111
+        15.75477235817033
+        108.8480554368229
+         13.1286184102431
+        18.33519591692408
+        108.9857739054074
+        11.84901811516484
+        13.26510395069653
+        15.67310192705747
+        107.8717937344275
+ 1.55e+10    
+        112.0124629832219
+        15.87037174946989
+        109.2548586695768
+        13.22846038462238
+        18.44374343097361
+        109.3972806860475
+        11.93585072519412
+        13.36558105793945
+        15.78872938270094
+        108.3332988446119
+ 1.56e+10    
+        112.4854840014754
+        15.98851911129769
+        109.6634049431845
+        13.32815612962406
+        18.55640875243758
+        109.8104739665452
+        12.02075134740058
+        13.46590763566186
+        15.90689920491331
+         108.794940737967
+ 1.57e+10    
+        112.9587517616598
+        16.10926620854299
+        110.0737889397838
+        13.42772009843773
+          18.673215984709
+        110.2254451323463
+        12.10371910481032
+        13.56609820619417
+        16.02766245511723
+        109.2567625542019
+ 1.58e+10    
+        113.4323115652357
+        16.23266096170184
+        110.4861011831801
+        13.52716604937699
+        18.79418160751446
+        110.6422814645236
+         12.1847542689571
+        13.66616660489514
+         16.1510663610246
+        109.7188064492638
+ 1.59e+10    
+        113.9062074937595
+         16.3587475021656
+        110.9004280581383
+        13.62650705016715
+        18.91931477422018
+        111.0610661585941
+        12.26385821069468
+        13.76612598426779
+        16.27715437252306
+         110.181113580032
+ 1.6e+10     
+        114.3804823984333
+        16.48756623386286
+        111.3168518368349
+        13.72575548456806
+        19.04861761623732
+        111.4818783505502
+        12.34103335240293
+        13.86598882040003
+        16.40596622389102
+        110.6437240921208
+ 1.61e+10    
+        114.8551778930019
+        16.61915390068845
+        111.7354507118826
+        13.82492306109431
+        19.18208555283769
+        111.9047931495372
+        12.41628312156004
+        13.96576692148821
+        16.53753800177502
+        111.1066771106468
+ 1.62e+10    
+        115.3303343498109
+        16.75354365917223
+        112.1562988353616
+        13.92402082359745
+        19.31970760478719
+        112.3298816766152
+        12.48961190564922
+        14.06547143821888
+        16.67190221838516
+        111.5700107337994
+ 1.63e+10    
+        115.8059908988478
+         16.8907651558618
+        112.5794663633219
+        14.02305916349435
+        19.46146671030755
+        112.7572111090859
+        12.56102500836991
+        14.16511287578583
+        16.80908788938013
+        112.0337620290596
+ 1.64e+10    
+        116.2821854295933
+        17.03084460891345
+        113.0050195052416
+        14.12204783344181
+        19.60734004197595
+        113.1868447298714
+        12.63052860712311
+        14.26470110734008
+        16.94912061593995
+        112.4979670319151
+ 1.65e+10    
+        116.7589545955049
+        17.17380489340679
+        113.4330205779541
+        14.22099596224814
+        19.75729932327097
+        113.6188419814659
+        12.69812971173703
+        14.36424538867346
+        17.09202267053975
+        112.9626607469252
+ 1.66e+10    
+        117.2363338209696
+        17.31966562992026
+        113.8635280635785
+         14.3199120708524
+        19.91131114357568
+        114.0532585240051
+          12.763836124405
+        14.46375437395976
+        17.23781308596454
+        113.4278771509867
+ 1.67e+10    
+        117.7143573105514
+         17.4684432759247
+        114.2965966710193
+        14.41880408918825
+        20.06933727053944
+        114.4901462970139
+        12.82765640080034
+        14.56323613237099
+        17.38650774712177
+        113.8936491986568
+ 1.68e+10    
+        118.1930580603855
+        17.62015121957721
+         114.732277400615
+        14.51767937377753
+        20.23133495880303
+        114.9295535844292
+         12.8895998123398
+        14.66269816541829
+        17.53811948523395
+        114.3600088293947
+ 1.69e+10    
+         118.672467871546
+        17.77479987551422
+        115.1706176115553
+        14.61654472590032
+        20.39725725417596
+        115.3715250825085
+        12.94967630956331
+         14.7621474248619
+        17.69265817401336
+        114.8269869765893
+ 1.7e+10     
+        119.1526173652516
+        17.93239678226923
+        115.6116610916968
+        14.71540641020617
+        20.56705329245213
+        115.8161019702598
+        13.00789648659898
+        14.86159033105497
+        17.85013082744076
+        115.2946135782312
+ 1.71e+10    
+        119.6335359997518
+        18.09294670095803
+         116.055448129438
+        14.81427017363437
+        20.74066859213035
+         116.263321982061
+        13.06427154668374
+        14.96103279159007
+        18.01054169879621
+        115.7629175891161
+ 1.72e+10    
+        120.1152520887552
+         18.2564517148969
+        116.5020155873361
+        14.91314126452873
+        20.91804534039425
+        116.7132194821404
+        13.11881326870987
+        15.06048022013569
+        18.17389238060402
+        116.2319269944426
+ 1.73e+10    
+        120.5977928212621
+        18.42291132983895
+        116.9513969771724
+        15.01202445183903
+        21.09912267178172
+        117.1658255406317
+        13.17153397476824
+        15.15993755535384
+        18.34018190518106
+        116.7016688246927
+ 1.74e+10    
+         121.081184282673
+         18.5923225745363
+        117.4036225361888
+        15.11092404430991
+        21.28383693905365
+        117.6211680109252
+        13.22244649865912
+          15.259409279799
+        18.50940684549266
+        117.1721691716817
+ 1.75e+10    
+        121.5654514770419
+        18.76468010135034
+        117.8587193042474
+        15.20984390956907
+        21.47212197584072
+        118.0792716080598
+        13.27156415534375
+        15.35889943871521
+        18.68156141604339
+        117.6434532056595
+ 1.76e+10    
+        122.0506183503554
+        18.93997628665705
+        118.3167112016781
+        15.30878749303709
+          21.663909350716
+        118.5401579879239
+        13.31890071130863
+        15.45841165864727
+        18.85663757354759
+        118.1155451933694
+ 1.77e+10    
+        122.5367078147263
+        19.11820133081016
+        118.7776191076022
+        15.40775783658773
+        21.85912861240833
+        119.0038458270464
+        13.36447035581706
+         15.5579491658002
+        19.03462511714185
+        118.5884685169511
+ 1.78e+10    
+        123.0237417733824
+        19.29934335744282
+        119.2414609385414
+        15.50675759689061
+        22.05770752592425
+        119.4703509027799
+        13.40828767302098
+        15.65751480408146
+        19.21551178792356
+        119.0622456936037
+ 1.79e+10    
+        123.5117411463548
+        19.48338851190585
+        119.7082517271272
+        15.60578906338892
+        22.25957229941104
+        119.9396861737005
+        13.45036761490906
+        15.75711105277065
+        19.39928336761263
+        119.5368983959073
+ 1.8e+10     
+        124.0007258967565
+        19.67032105865942
+        120.1780037007603
+         15.7048541758601
+        22.46464780163941
+         120.411861860048
+        13.49072547506735
+        15.85674004377246
+        19.58592377615173
+        120.0124474727195
+ 1.81e+10    
+        124.4907150575672
+        19.86012347744736
+          120.65072636007
+        15.80395454151682
+        22.67285777003545
+        120.8868855240711
+        13.52937686322762
+        15.95640357841149
+        19.77541516807984
+        120.4889129705658
+ 1.82e+10    
+        124.9817267588226
+        20.05277655810323
+        121.1264265570489
+        15.90309145161376
+          22.884125009234
+        121.3647621501297
+        13.56633768058148
+        16.05610314372529
+         19.9677380275217
+        120.9663141554422
+ 1.83e+10    
+        125.4737782551335
+        20.24825949384824
+         121.605108572742
+        16.00226589753608
+        23.09837158017017
+        121.8454942244416
+        13.60162409583941
+        16.15583992824614
+        20.16287126165891
+        121.4446695349567
+ 1.84e+10    
+        125.9668859534491
+        20.44654997295725
+        122.0867741943982
+        16.10147858633907
+        23.31551897975818
+        122.3290818143675
+        13.63525252201124
+         16.2556148372262
+        20.36079229255772
+        121.9239968807383
+ 1.85e+10    
+        126.4610654409881
+        20.64762426868155
+        122.5714227919858
+        16.20072995572403
+        23.53548831124294
+        122.8155226471237
+        13.66723959389029
+        16.35542850730697
+        20.56147714724153
+        122.4043132510527
+ 1.86e+10    
+        126.9563315132722
+        20.85145732733128
+        123.0590513939996
+        16.30002018843579
+        23.75820044534031
+        123.3048121878562
+        13.69760214621878
+        16.45528132060472
+        20.76490054591164
+        122.8856350135513
+ 1.87e+10    
+        127.4526982021926
+        21.05802285443226
+        123.5496547624972
+        16.39934922607235
+        23.98357617230963
+        123.7969437169909
+        13.72635719251793
+         16.5551734182139
+        20.97103598823142
+        123.3679778681098
+ 1.88e+10    
+        127.9501788040449
+        21.26729339887905
+        124.0432254672955
+        16.49871678230094
+         24.2115363451229
+        124.2919084067952
+        13.75352190456272
+        16.65510471311593
+        21.17985583759669
+        123.8513568696885
+ 1.89e+10    
+        128.4487859074785
+        21.47924043502561
+         124.539753959295
+        16.59812235547844
+        24.44200201392141
+        124.7896953971012
+        13.77911359248493
+        16.75507490249806
+        21.39133140333167
+        124.3357864511718
+ 1.9e+10     
+         128.948531421306
+         21.6938344426569
+        125.0392286428832
+        16.69756524067669
+        24.67489455196392
+        125.2902918701371
+        13.80314968548573
+         16.8550834794737
+        21.60543302075566
+        124.8212804461352
+ 1.91e+10    
+        129.4494266021223
+        21.91104498479819
+        125.5416359473913
+        16.79704454111534
+        24.91013577329119
+        125.7936831244325
+        13.82564771314357
+        16.95512974422162
+        21.82213012907687
+        125.3078521114994
+ 1.92e+10    
+        129.9514820816844
+        22.13084078332793
+         126.046960397578
+        16.89655917901355
+        25.14764804234163
+        126.2998526477602
+        13.84662528729985
+        17.05521281453984
+        22.04139134707872
+        125.7955141500231
+ 1.93e+10    
+        130.4547078940161
+        22.35318979236759
+        126.5551846831275
+        16.99610790586328
+         25.3873543757659
+        126.8087821890915
+        13.86610008450843
+        17.15533163583134
+        22.26318454657213
+        126.2842787326105
+ 1.94e+10    
+        130.9591135021913
+        22.57805926942816
+         127.066289727143
+        17.09568931213688
+          25.629178536696
+        127.3204518295422
+        13.88408982903284
+        17.25548499052478
+        22.48747692359367
+        126.7741575203798
+ 1.95e+10    
+        131.4647078247637
+        22.80541584430341
+        127.5802547536378
+        17.19530183644633
+         25.8730451217355
+        127.8348400522966
+        13.90061227637904
+        17.35567150695246
+        22.71423506734152
+        127.2651616864807
+ 1.96e+10    
+        131.9714992618132
+        23.03522558570736
+        128.0970573540226
+        17.29494377415903
+        26.11887964093608
+        128.3519238114965
+         13.9156851973486
+        17.45588966769231
+        22.94342502683886
+         127.757301937616
+ 1.97e+10    
+        132.4794957205702
+        23.26745406565135
+         128.616673552583
+        17.39461328549493
+        26.36660859103667
+        128.8716786000863
+         13.9293263625998
+         17.5561378173926
+        23.17501237533178
+        128.2505885352502
+ 1.98e+10    
+        132.9887046406025
+        23.50206642157413
+         129.139077870966
+        17.49430840311236
+        26.61615952223865
+         129.394078516621
+        13.94155352770399
+        17.65641417009803
+        23.40896227242522
+        128.7450313164758
+ 1.99e+10    
+         133.499133018534
+        23.73902741623506
+        129.6642433916776
+        17.59402703920934
+        26.86746109879386
+         129.919096331023
+        13.95238441868548
+          17.756716816091
+        23.64523952396942
+        129.2406397145211
+ 2e+10       
+        134.0107874322737
+        23.97830149538735
+        130.1921418206098
+        17.69376699214952
+         27.1204431536809
+        130.4467035493045
+        13.96183671803232
+        17.85704372826964
+        23.88380863971616
+        129.7374227788733
+ 2.01e+10    
+        134.5236740647376
+        24.21985284325295
+        130.7227435486058
+        17.79352595263741
+        27.37503673764291
+        130.9768704772511
+        13.96992805116766
+        17.95739276807862
+          24.124633888763
+        130.2353891950048
+ 2.02e+10    
+        135.0377987270514
+        24.46364543582681
+        131.2560177120892
+        17.89330150945818
+        27.63117416286092
+        131.5095662830834
+           13.97667597337
+        18.05776169101711
+        24.36767935281406
+        130.7345473036868
+ 2.03e+10    
+        135.5531668812108
+        24.70964309203737
+         131.791932252768
+        17.99309115480385
+        27.88878904152707
+        132.0447590590915
+        13.98209795713241
+        18.15814815173539
+        24.61290897728284
+        131.2349051198752
+ 2.04e+10    
+        136.0697836621916
+        24.95780952279615
+        132.3304539764377
+        18.09289228920436
+        28.14781631958533
+         132.582415882273
+        13.98621137995042
+        18.25854970874962
+        24.86028662027295
+         131.736470351157
+ 2.05e+10    
+        136.5876538995037
+         25.2081083779745
+        132.8715486109054
+        18.19270222608103
+        28.40819230589519
+        133.1225028739668
+        13.98903351252843
+        18.35896382878483
+        25.10977609946759
+        132.2392504157522
+ 2.06e+10    
+         137.106782138174
+        25.46050329134072
+        133.4151808630556
+        18.29251819594234
+        28.66985469707426
+          133.66498525851
+        13.99058150739483
+        18.45938789077251
+        25.36134123696937
+        132.7432524600539
+ 2.07e+10    
+        137.6271726591522
+        25.71495792350127
+        133.9613144750741
+        18.39233735024741
+        28.93274259826489
+        134.2098274209191
+        13.99087238791866
+        18.55981918952074
+        25.61494590212562
+        133.2484833757136
+ 2.08e+10    
+        138.1488294991392
+        25.97143600288644
+        134.5099122798647
+        18.49215676494346
+        29.19679654006591
+        134.7569929636197
+        13.98992303771541
+        18.66025493907189
+        25.87055405238493
+        133.7549498162495
+ 2.09e+10    
+        138.6717564698306
+        26.22990136482466
+        135.0609362556678
+         18.5919734437072
+        29.46195849186367
+        135.3064447622307
+        13.98775019043684
+        18.76069227577495
+         26.1281297722252
+        134.2626582131897
+ 2.1e+10     
+        139.1959571765732
+        26.49031798875028
+        135.6143475799117
+        18.69178432090498
+        29.72817187178754
+        135.8581450204186
+        13.98437041993414
+        18.86112826108122
+        26.38763731019836
+        134.7716147917375
+ 2.11e+10    
+        139.7214350364362
+        26.75265003358976
+        136.1701066823103
+        18.79158626428357
+        29.99538155350918
+        136.4120553238373
+        13.97980013078725
+        18.96155988409077
+        26.64904111413819
+        135.2818255859618
+ 2.12e+10    
+        140.2481932956958
+        27.01686187137524
+         136.728173297235
+        18.89137607741949
+        30.26353387009641
+        136.9681366931624
+        13.97405554919197
+        19.06198406385714
+        26.91230586457696
+        135.7932964535119
+ 2.13e+10    
+        140.7762350467335
+        27.28291811913286
+         137.288506515377
+        18.99115050193486
+        30.53257661512574
+        137.5263496362378
+         13.9671527141979
+        19.16239765147948
+        27.17739650641904
+        136.3060330898543
+ 2.14e+10    
+        141.3055632443557
+        27.55078366909071
+        137.8510648347136
+        19.09090621949903
+        30.80245904124664
+        138.0866541993378
+        13.95910746928894
+        19.26279743198629
+        27.44427827891662
+        136.8200410420366
+ 2.15e+10    
+        141.8361807215326
+        27.82042371726046
+        138.4158062108051
+        19.19063985363375
+        31.07313185638751
+        138.6490100175668
+        13.94993545429914
+        19.36318012603348
+        27.71291674399997
+        137.3353257219783
+ 2.16e+10    
+        142.3680902045624
+        28.09180379043642
+        138.9826881064321
+        19.29034797133082
+        31.34454721778099
+        139.2133763643971
+        13.93965209765786
+        19.46354239143422
+        27.98327781300718
+         137.851892419295
+ 2.17e+10    
+        142.9012943276705
+        28.36488977166389
+        139.5516675405893
+        19.39002708450656
+        31.61665872398042
+        139.7797122003584
+        13.92827260895563
+        19.56388082452521
+         28.2553277718618
+        138.3697463136559
+ 2.18e+10    
+        143.4357956470422
+        28.63964792422209
+        140.1227011368483
+        19.48967365129431
+         31.8894214050306
+        140.3479762208884
+        13.91581197182534
+        19.66419196139516
+        28.52903330474825
+        138.8888924866793
+ 2.19e+10    
+        143.9715966543054
+        28.91604491417415
+        140.6957451711047
+        19.58928407720052
+        32.16279171094988
+        140.9181269033491
+        13.90228493713168
+        19.76447227898027
+         28.8043615163316
+        139.4093359333771
+ 2.2e+10     
+        144.5086997894578
+        29.19404783152793
+        141.2707556187145
+        19.68885471612692
+        32.43672749866938
+        141.4901225532156
+        13.88770601646207
+        19.86471819604359
+         29.0812799525696
+        139.9310815731451
+ 2.21e+10    
+        145.0471074532622
+        29.47362421005569
+        141.8476882010296
+        19.78838187127899
+         32.7111880175723
+        142.0639213494457
+        13.87208947591348
+         19.9649260740476
+        29.35975662016416
+        140.4541342603139
+ 2.22e+10    
+        145.5868220191036
+        29.75474204582284
+        142.4264984313438
+        19.88786179596293
+        32.98613389376385
+        142.6394813890282
+          13.855449330168
+        20.06509221793435
+         29.6397600046983
+        140.9784987942577
+ 2.23e+10    
+        146.1278458443283
+        30.03736981446638
+        143.0071416602503
+        19.98729069429279
+        33.26152711320076
+        143.2167607307209
+        13.83779933685237
+         20.1652128768208
+        29.92125908750488
+         141.504179929081
+ 2.24e+10    
+        146.6701812810664
+        30.32147648727224
+        143.5895731204096
+        20.08666472180735
+        33.53733100379589
+        143.7957174379726
+         13.8191529911746
+        20.26528424462359
+        30.20422336131244
+        142.0311823828739
+ 2.25e+10    
+        147.2138306865543
+        30.60703154609419
+        144.1737479707415
+        20.18597998601279
+        33.81351021661251
+        144.3763096210355
+        13.79952352083155
+        20.36530246061357
+        30.48862284471165
+        142.5595108465598
+ 2.26e+10    
+        147.7587964329586
+         30.8940049971578
+        144.7596213400292
+        20.28523254685783
+        34.09003070625235
+        144.9584954782653
+        13.77892388118339
+        20.46526360992381
+        30.77442809548692
+        143.0891699923338
+ 2.27e+10    
+        148.3050809167246
+        31.18236738379314
+        145.3471483699437
+          20.384418417149
+        34.36685971053699
+        145.5422333366069
+        13.75736675068756
+        20.56516372400344
+        31.06161022285479
+        143.6201644817008
+ 2.28e+10    
+        148.8526865674438
+        31.47208979813636
+        145.9362842574748
+        20.48353356291509
+        34.64396572957454
+         146.127481691267
+        13.73486452658764
+        20.66499878103559
+        31.35014089865201
+        144.1524989731255
+ 2.29e+10    
+        149.4016158562634
+        31.76314389184089
+        146.5269842967737
+        20.58257390372727
+        34.92131850429973
+        146.7141992445662
+        13.71142932085193
+        20.76476470632317
+        31.63999236751285
+        144.6861781293025
+ 2.3e+10     
+        149.9518713038475
+        32.05550188583928
+        147.1192039203952
+        20.68153531298097
+        35.19888899456706
+        147.3023449439698
+        13.68707295635542
+        20.86445737264732
+        31.93113745607575
+        145.2212066240498
+ 2.31e+10    
+        150.5034554878929
+        32.34913657919132
+        147.7128987399296
+        20.78041361814902
+        35.47664935687306
+        147.8918780192895
+        13.66180696330154
+        20.96407260060732
+        32.22354958125775
+        145.7575891488397
+ 2.32e+10    
+        151.0563710502168
+        32.64402135705839
+        148.3080245860239
+        20.87920460100315
+        35.75457292177862
+        148.4827580190537
+        13.63564257587654
+        21.06360615894588
+        32.51720275763668
+        146.2953304189771
+ 2.33e+10    
+         151.610620703431
+        32.94013019783819
+         148.904537547767
+        20.97790399782219
+        36.03263417109468
+        149.0749448460348
+        13.60859072913338
+        21.16305376486375
+        32.81207160397222
+        146.8344351794284
+ 2.34e+10    
+        152.1662072372044
+        33.23743767949637
+         149.502394011441
+         21.0765074995783
+        36.31080871489319
+        149.6683987919322
+        13.58066205609901
+         21.2624110843314
+        33.10813134890847
+        147.3749082103161
+ 2.35e+10    
+        152.7231335241326
+        33.53591898512774
+        150.1015506986168
+        21.17501075211575
+        36.58907326839952
+        150.2630805711995
+        13.55186688510066
+            21.3616737324
+        33.40535783588699
+         147.916754332085
+ 2.36e+10    
+         153.281402525221
+         33.8355499077795
+        150.7019647035754
+        21.27340935631765
+        36.86740562881353
+        150.8589513540051
+        13.52221523730521
+        21.46083727350987
+        33.70372752730505
+        148.4599784103473
+ 2.37e+10    
+        153.8410172949983
+        34.13630685457068
+        151.3035935300542
+        21.37169886827284
+        37.14578465211267
+        151.4559727983234
+        13.49171682446917
+        21.55989722181171
+        34.00321750795413
+        149.0045853604225
+ 2.38e+10    
+        154.4019809862645
+        34.43816685013508
+        151.9063951272812
+        21.46987479943774
+        37.42419022987401
+        152.0541070811435
+        13.46038104689217
+        21.65884904149328
+        34.30380548776583
+        149.5505801515727
+ 2.39e+10    
+        154.9642968544877
+        34.74110753941868
+        152.5103279252963
+        21.56793261680445
+        37.70260326615943
+         152.653316928786
+        13.42821699157114
+        21.75768814711503
+        34.60546980389807
+        150.0979678109474
+ 2.4e+10     
+        155.5279682618634
+        35.04510718985944
+        153.1153508695304
+        21.66586774306584
+        37.98100565449541
+        153.2535656463147
+        13.39523343054896
+        21.85640990396206
+        34.90818942219138
+        150.6467534272481
+ 2.41e+10    
+        156.0929986810436
+        35.35014469297793
+        153.7214234546261
+        21.76367555679363
+        38.25938025498301
+        153.8548171460432
+        13.36143881945497
+         21.9550096284082
+        35.21194393801986
+        151.1969421541155
+ 2.42e+10    
+        156.6593916985451
+         35.6561995654025
+        154.3285057574812
+        21.86135139262149
+          38.537710871566
+        154.4570359751115
+        13.32684129623161
+         22.0534825882971
+        35.51671357656782
+        151.7485392132528
+ 2.43e+10    
+        157.2271510178535
+        35.96325194935519
+        154.9365584694901
+        21.95889054143513
+        38.81598222948234
+        155.0601873421366
+         13.2914486800431
+        22.15182400334171
+        35.82247919255711
+        152.3015498972941
+ 2.44e+10    
+         157.796280462225
+        36.27128261262442
+        155.5455429279682
+        22.05628825057929
+        39.09417995292438
+        155.6642371429149
+        13.25526847036226
+        22.25002904553763
+        36.12922226944858
+        152.8559795724227
+ 2.45e+10    
+         158.366783977207
+        36.58027294804395
+         156.155421146729
+        22.15353972406902
+        39.37229054292611
+        156.2691519851756
+        13.21830784623075
+        22.34809283959961
+         36.4369249181451
+        153.4118336807529
+ 2.46e+10    
+        158.9386656328778
+        36.89020497250323
+        156.7661558458032
+        22.25064012281952
+        39.65030135549847
+        156.8748992123677
+        13.18057366568918
+        22.44601046341479
+        36.74556987521644
+        153.9691177424781
+ 2.47e+10    
+        159.5119296258184
+        37.20106132550819
+        157.3777104802639
+         22.3475845648863
+        39.92820058002513
+        157.4814469264747
+        13.14207246537196
+        22.54377694851233
+        37.05514050067091
+        154.5278373577964
+ 2.48e+10    
+        160.0865802808303
+        37.51282526731478
+        157.9900492681506
+         22.4443681257195
+        40.20597721793636
+        158.0887640098501
+        13.10281046026445
+        22.64138728055749
+        37.36562077529336
+        155.0879982086244
+ 2.49e+10    
+        160.6626220524055
+         37.8254806766527
+        158.6031372174614
+        22.54098583843258
+         40.4836210616688
+        158.6968201460546
+        13.06279354361639
+        22.73883639985718
+        37.67699529757189
+        155.6496060601004
+ 2.5e+10     
+        161.2400595259564
+        38.13901204805883
+        159.2169401521903
+        22.63743269408342
+        40.76112267392518
+        159.3055858397037
+        13.02202728700949
+         22.8361192018889
+        37.98924928023266
+        156.2126667618925
+ 2.51e+10    
+        161.8188974188186
+        38.45340448883875
+        159.8314247373969
+        22.73370364197083
+        41.03847336723799
+        159.9150324352936
+        12.98051694057441
+        22.93323053784591
+        38.30236854640108
+        156.7771862493097
+ 2.52e+10    
+         162.399140581035
+         38.7686437156713
+        160.4465585032791
+        22.82979358994552
+        41.31566518384704
+        160.5251321350265
+        12.93826743335335
+        23.03016521519498
+        38.61633952540944
+        157.3431705442375
+ 2.53e+10    
+        162.9807939959275
+        39.08471605087529
+        161.0623098682325
+        22.92569740473234
+        41.59269087589386
+        161.1358580156029
+        12.89528337380503
+        23.12691799825763
+        38.93114924826749
+        157.9106257558888
+ 2.54e+10    
+        163.5638627804683
+        39.40160841834958
+        161.6786481608771
+        23.02140991226504
+        41.86954388593753
+         161.747184043991
+        12.85156905044689
+        23.22348360879637
+        39.24678534281236
+        158.4795580813912
+ 2.55e+10    
+        164.1483521854574
+        39.71930833920683
+         162.295543641029
+        23.11692589803813
+        42.14621832779497
+         162.359085092163
+        12.80712843263333
+        23.31985672662267
+        39.56323602855648
+        159.0499738062096
+ 2.56e+10    
+        164.7342675955165
+        40.03780392710989
+        162.9129675196058
+        23.21224010746476
+        42.42270896770579
+        162.9715369507891
+        12.76196517146412
+        23.41603199021499
+        39.88049011124512
+        159.6218793044119
+ 2.57e+10    
+        165.3216145289021
+        40.35708388332786
+        163.5308919774405
+        23.30734724625085
+        42.69901120582363
+        163.5845163419002
+        12.71608260082034
+        23.51200399734446
+        40.19853697714527
+        160.1952810387941
+ 2.58e+10    
+        165.9103986371584
+        40.67713749152285
+         164.149290182992
+        23.40224198077649
+        42.97512105803177
+        164.1980009304966
+        12.66948373852456
+        23.60776730571488
+        40.51736658706979
+        160.7701855608482
+ 2.59e+10    
+         166.500625704596
+        40.99795461227943
+        164.7681363089383
+         23.4969189384882
+        43.25103513808325
+        164.8119693351198
+        12.62217128762166
+        23.70331643361144
+        40.83696947016315
+        161.3465995106124
+ 2.6e+10     
+         167.092301647632
+        41.31952567739214
+        165.3874055476352
+        23.59137270830183
+        43.52675064006288
+        165.4264011373731
+        12.57414763777664
+        23.79864586055341
+        41.15733671745062
+        161.9245296163768
+ 2.61e+10    
+        167.6854325139714
+        41.64184168391685
+        166.0070741254308
+        23.68559784101161
+        43.80226532116729
+        166.0412768904042
+        12.52541486678644
+        23.89375002795442
+        41.47845997517246
+        162.5039826942757
+ 2.62e+10    
+         168.280024481659
+        41.96489418800174
+        166.6271193158234
+        23.77958884970806
+        44.07757748480181
+        166.6565781263385
+        12.47597474220239
+        23.98862333978794
+        41.80033143790956
+        163.0849656477573
+ 2.63e+10    
+        168.8760838579917
+         42.2886752985055
+        167.2475194514536
+        23.87334021020109
+        44.35268596398824
+        167.2722873626739
+        12.42582872306023
+        24.08326016325564
+        42.12294384151534
+        163.6674854669419
+ 2.64e+10    
+        169.4736170783111
+        42.61317767041348
+        167.8682539349198
+         23.9668463614501
+        44.62759010508107
+        167.8883881076443
+        12.37497796171385
+         24.1776548294566
+        42.44629045586383
+        164.2515492278755
+ 2.65e+10    
+         170.072630704676
+        42.93839449806229
+        168.4893032484167
+        24.06010170599958
+         44.9022897517856
+        168.5048648645423
+        12.32342330577104
+        24.27180163405765
+         42.7703650774262
+         164.837164091686
+ 2.66e+10    
+        170.6731314244205
+        43.26431950818066
+        169.1106489621825
+         24.1531006104165
+         45.1767852294753
+        169.1217031350286
+        12.27116530012652
+        24.36569483796185
+         43.0951620216847
+        165.4243373036334
+ 2.67e+10    
+        171.2751260486081
+         43.5909469527567
+        169.7322737417623
+        24.24583740573278
+        45.45107732980119
+        169.7388894214134
+         12.2182041890906
+        24.45932866797739
+        43.42067611539549
+         166.013076192082
+ 2.68e+10    
+        171.8786215103862
+        43.91827160173901
+        170.3541613540734
+        24.33830638789064
+        45.72516729558881
+        170.3564112279374
+        12.16453991860975
+        24.55269731747729
+        43.74690268870976
+        166.6033881673814
+ 2.69e+10    
+        172.4836248632461
+        44.24628873558121
+        170.9762966722834
+        24.43050181818608
+        45.99905680601694
+        170.9742570610471
+        12.11017213857654
+         24.6457949470629
+        44.07383756716074
+        167.1952807206639
+ 2.7e+10     
+        173.0901432791912
+        44.57499413763753
+        171.5986656794986
+        24.52241792371898
+        46.27274796207272
+        171.5924164286886
+        12.05510020522576
+        24.73861568521097
+        44.40147706352968
+        167.7887614225718
+ 2.71e+10    
+        173.6981840468274
+        44.90438408641634
+        172.2212554712634
+        24.61404889783694
+        46.54624327227765
+        172.2108798386209
+        11.99932318361442
+        24.83115362892337
+         44.7298179695964
+        168.3838379219135
+ 2.72e+10    
+        174.3077545693726
+        45.23445534770181
+          172.84405425688
+        24.70538890058449
+         46.8195456386774
+        172.8296387957705
+        11.94283985018267
+        24.92340284436235
+        45.05885754778294
+        168.9805179442469
+ 2.73e+10    
+        174.9188623625939
+        45.56520516654625
+        173.4670513595538
+        24.79643205914677
+        47.09265834309087
+        173.4486857986358
+        11.88564869539238
+        25.01535736747793
+        45.38859352270005
+        169.5788092904036
+ 2.74e+10    
+        175.5315150526775
+        45.89663125914727
+        174.0902372153732
+        24.88717246829276
+        47.36558503361354
+        174.0680143347605
+        11.82774792644196
+        25.10701120462817
+        45.71902407260458
+        170.1787198349582
+ 2.75e+10    
+         176.145720374035
+        46.22873180460986
+        174.7136033711347
+        24.97760419081687
+        47.63832971136633
+        174.6876188752922
+        11.76913547005343
+        25.19835833318285
+        46.05014782077352
+        170.7802575246354
+ 2.76e+10    
+        176.7614861670507
+        46.56150543660464
+        175.3371424810249
+        25.06772125797703
+        47.91089671748831
+        175.3074948686435
+        11.70980897533049
+        25.28939270212081
+        46.38196382680432
+        171.3834303766731
+ 2.77e+10    
+         177.378820375781
+        46.89495123492887
+        175.9608483021776
+        25.15751766992783
+         48.1832907203655
+        175.9276387332743
+        11.64976581668397
+        25.38010823261137
+        46.71447157784748
+        171.9882464771337
+ 2.78e+10    
+        177.9977310455928
+        47.22906871697301
+        176.5847156891114
+         25.2469873961524
+        48.45551670308983
+        176.5480478496163
+        11.58900309682292
+        25.47049881858292
+        47.04767097977838
+        172.5947139791755
+ 2.79e+10    
+        178.6182263207692
+        47.56385782910481
+        177.2087405870796
+        25.33612437588934
+        48.72757995114539
+          177.16872055116
+        11.52751764980903
+        25.56055832727865
+        47.38156234831732
+        173.2028411012816
+ 2.8e+10     
+        179.2403144420626
+        47.89931893797272
+        177.8329200243409
+        25.42492251855089
+        48.99948604031497
+        177.7896561147259
+        11.46530604417103
+        25.65028059979734
+        47.71614640010085
+        173.8126361254524
+ 2.81e+10    
+        179.8640037442216
+        48.23545282173785
+        178.4572521033773
+        25.51337570414312
+        49.27124082480294
+         178.410854749942
+        11.40236458607826
+        25.73965945161936
+        48.05142424371405
+        174.4241073953688
+ 2.82e+10    
+        180.4893026534712
+        48.57226066123923
+        179.0817359910763
+        25.60147778367545
+        49.54285042556923
+        179.0323175879547
+        11.33868932256975
+        25.82868867311728
+        48.38739737068845
+        175.0372633145161
+ 2.83e+10    
+        181.1162196849758
+        48.90974403109823
+         179.706371907907
+        25.68922257956648
+        49.81432121887075
+         179.654046669392
+        11.27427604483761
+        25.91736203005062
+        48.72406764647233
+        175.6521123442906
+ 2.84e+10    
+        181.7447634402655
+         49.2479048907703
+        180.3311611161182
+        25.77660388604554
+        50.08565982500565
+        180.2760449316121
+        11.20912029156187
+        26.00567326404683
+        49.06143730137924
+        176.2686630020741
+ 2.85e+10    
+        182.3749426046446
+        49.58674557554619
+        180.9561059069677
+        25.86361546954397
+        50.35687309725498
+        180.8983161952515
+        11.14321735229495
+        26.09361609306398
+        49.39950892152009
+        176.8869238592907
+ 2.86e+10    
+        183.0067659445739
+        49.92626878751312
+        181.5812095870386
+        25.95025106908783
+         50.6279681110209
+        181.5208651501132
+        11.07656227089399
+        26.18118421183944
+        49.73828543972571
+        177.5069035394424
+ 2.87e+10    
+        183.6402423050483
+         50.2664775864784
+        182.2064764636477
+        26.03650439667823
+        50.89895215315437
+        182.1436973404112
+        11.00914984899832
+        26.26837129232092
+        50.07777012646388
+        178.1286107161316
+ 2.88e+10    
+        184.2753806069406
+        50.60737538086155
+        182.8319118293882
+        26.12236913766746
+        51.16983271147171
+         182.766819149406
+        10.94097464955026
+        26.35517098408386
+         50.4179665807577
+        178.7520541110625
+ 2.89e+10    
+        184.9121898443549
+        50.94896591856383
+        183.4575219458406
+          26.207838951132
+        51.44061746445472
+        183.3902377834523
+        10.87203100035814
+        26.44157691473133
+         50.7588787211096
+         179.377242492039
+ 2.9e+10     
+        185.5506790819533
+        51.29125327781443
+        184.0833140264744
+        26.29290747023742
+        51.71131427113296
+        184.0139612554981
+        10.80231299769833
+        26.52758269027896
+        51.10051077643623
+         180.004184670946
+ 2.91e+10    
+         186.190857452289
+        51.63424185800719
+        184.7092962187885
+        26.37756830259846
+        51.98193116114437
+        184.6379983680524
+        10.73181450995532
+        26.61318189552528
+        51.44286727701977
+        180.6328895017303
+ 2.92e+10    
+        186.8327341531279
+        51.97793637052626
+        185.3354775857091
+        26.46181503063114
+         52.2524763249711
+        185.2623586956599
+        10.66052918129749
+        26.69836809440676
+        51.78595304548021
+        181.2633658783668
+ 2.93e+10    
+        187.4763184447727
+         52.3223418295695
+        185.9618680862973
+        26.54564121190492
+        52.52295810435076
+        185.8870525669089
+        10.58845043538752
+        26.78313483033806
+        52.12977318777371
+        181.8956227328341
+ 2.94e+10    
+        188.1216196473878
+        52.66746354297519
+        186.5884785557865
+         26.6290403794855
+        52.79338498285677
+        186.5120910460008
+        10.51557147912462
+        26.86747562653865
+        52.47433308421988
+        182.5296690330736
+ 2.95e+10    
+        188.7686471383234
+         53.0133071030555
+        187.2153206849994
+        26.71200604227486
+        53.06376557664981
+         187.137485913913
+        10.44188530641786
+        26.95138398634551
+        52.81963838056558
+        183.1655137809629
+ 2.96e+10    
+        189.4174103494498
+        53.35987837744437
+        187.8424069991754
+        26.79453168534438
+         53.3341086253953
+        187.7632496491879
+        10.36738470198822
+        27.03485339351323
+        53.16569497908811
+        183.8031660102828
+ 2.97e+10    
+        190.0679187644963
+        53.70718349996363
+        188.4697508362494
+        26.87661077026885
+        53.60442298334817
+        188.3893954083713
+        10.29206224519869
+        27.11787731250246
+        53.51250902973949
+        184.4426347846902
+ 2.98e+10    
+        190.7201819163971
+        54.05522886151102
+        189.0973663246134
+        26.95823673545152
+        53.87471761059987
+        189.0159370061383
+        10.21591031390905
+        27.20044918875339
+        53.86008692134206
+        185.0839291956962
+ 2.99e+10    
+        191.3742093846517
+         54.4040211009794
+        189.7252683604131
+        27.03940299644814
+        54.14500156448995
+        189.6428888951305
+        10.13892108835589
+         27.2825624489522
+        54.20843527283318
+         185.727058360654
+ 3e+10       
+        192.0300107926962
+         54.7535670962071
+        190.3534725843985
+        27.12010294628776
+        54.41528399117749
+        190.2702661455347
+          10.061086555055
+         27.3642105012845
+         54.5575609245664
+        186.3720314207496
+ 3.01e+10    
+         192.687595805285
+        55.10387395496878
+        190.9819953583922
+        27.20032995579123
+        54.68557411737439
+        190.8980844244411
+        9.982398510724694
+        27.44538673567902
+        54.90747092967226
+        187.0188575390059
+ 3.02e+10    
+        193.3469741258964
+        55.45494900600774
+        191.6108537413874
+        27.28007737388564
+        54.95588124223707
+        191.5263599749967
+        9.902848566229451
+        27.52608452404388
+        55.25817254548247
+         187.667545898298
+ 3.03e+10    
+        194.0081554941439
+        55.80679979011691
+        192.2400654653324
+        27.35933852792046
+         55.2262147294165
+        192.1551095953925
+        9.822428150541477
+        27.60629722049256
+         55.6096732250197
+        188.3181056993772
+ 3.04e+10    
+        194.6711496832173
+        56.15943405127321
+        192.8696489106391
+        27.43810672397765
+         55.4965839992669
+        192.7843506177155
+        9.741128514719319
+        27.68601816156438
+        55.96198060855851
+        188.9705461589108
+ 3.05e+10    
+        195.3359664973349
+        56.51285972782699
+        193.4996230814412
+        27.51637524718617
+        55.76699852121033
+        193.4141008866827
+        9.658940735902423
+        27.76524066643652
+        56.31510251525991
+        189.6248765075383
+ 3.06e+10    
+        196.0026157692216
+        56.86708494375522
+        194.1300075806564
+        27.59413736202958
+        56.03746780625793
+         194.044378738296
+        9.575855721319192
+        27.84395803713179
+        56.66904693488194
+        190.2811059879379
+ 3.07e+10    
+        196.6711073576049
+        57.22211799997825
+        194.7608225848742
+         27.6713863126602
+        56.30800139968777
+        194.6752029784406
+        9.491864212309117
+        27.92216355872116
+        57.02382201956964
+        190.9392438529136
+ 3.08e+10    
+        197.3414511447382
+        57.57796736574765
+         195.392088819121
+        27.74811532321023
+        56.57860887387641
+        195.3065928614522
+        9.406956788355711
+        27.99985049951955
+        57.37943607572882
+        191.5992993634972
+ 3.09e+10    
+        198.0136570339461
+        57.93464167010801
+        196.0238275315284
+        27.82431759810215
+        56.84929982128654
+        195.9385680686831
+        9.321123871130331
+        28.07701211128381
+        57.73589755598401
+        192.2612817870704
+ 3.1e+10     
+        198.6877349471948
+        58.29214969343584
+        196.6560604679444
+        27.89998632236516
+        57.12008384760873
+        196.5711486870917
+        9.234355728545424
+        28.15364162940077
+        58.09321505122632
+        192.9252003955054
+ 3.11e+10    
+        199.3636948226884
+        58.65050035906174
+        197.2888098465237
+        27.97511466194896
+        57.39097056505769
+        197.2043551878814
+        9.146642478815632
+        28.22973227308111
+        58.45139728275056
+         193.591064463324
+ 3.12e+10    
+         200.041546612494
+        59.00970272497428
+        197.9220983323291
+        28.04969576404163
+        57.66196958582066
+        197.8382084052042
+        9.057974094525953
+        28.30527724554719
+        58.81045309448522
+        194.2588832658777
+ 3.13e+10    
+        200.7213002801887
+        59.36976597561791
+        198.5559490119806
+        28.12372275739123
+         57.9330905156624
+        198.4727295149751
+        8.968340406705874
+        28.38026973422234
+        59.17039144532067
+        194.9286660775515
+ 3.14e+10    
+         201.402965798545
+        59.73069941377826
+        199.1903853683794
+        28.19718875262799
+        58.20434294767962
+        199.1079400137907
+        8.877731108908215
+        28.45470291092188
+        59.53122140153211
+        195.6004221699854
+ 3.15e+10    
+        202.0865531472375
+        60.09251245256603
+        199.8254312555467
+         28.2700868425922
+        58.47573645621105
+        199.7438616979981
+        8.786135761291785
+        28.52856993204485
+        59.89295212930426
+         196.274160810324
+ 3.16e+10    
+        202.7720723105789
+        60.45521460749796
+        200.4611108736021
+        28.34241010266436
+          58.747280590899
+        200.3805166429245
+          8.6935437947062
+        28.60186393876736
+        60.25559288735705
+        196.9498912594798
+ 3.17e+10    
+        203.4595332752918
+        60.81881548867992
+        201.0974487439117
+        28.41415159110164
+        59.01898487090306
+        201.0179271822909
+        8.599944514779175
+         28.6745780572403
+        60.61915301967525
+        197.6276227704318
+ 3.18e+10    
+        204.1489460283072
+         61.1833247930939
+        201.7344696844363
+        28.48530434937675
+        59.29085877926605
+        201.6561158878305
+        8.505327106003929
+        28.74670539879098
+        60.98364194834376
+        198.3073645865379
+ 3.19e+10    
+        204.8403205545957
+        61.54875229699307
+        202.3721987853136
+        28.55586140252309
+         59.5629117574309
+        202.2951055491245
+        8.409680635826229
+        28.81823906012701
+        61.34906916648998
+        198.9891259398788
+ 3.2e+10     
+        205.5336668350307
+        61.91510784840489
+        203.0106613846838
+        28.62581575948596
+        59.83515319990946
+        202.9349191536868
+        8.312994058730673
+         28.8891721235489
+        61.71544423133308
+        199.6729160496223
+ 3.21e+10    
+        206.2289948442823
+        62.28240135974661
+         203.649883044805
+        28.69516041347786
+        60.10759244910127
+        203.5755798672996
+        8.215256220324166
+        28.95949765716476
+        62.08277675734613
+        200.3587441204143
+ 3.22e+10    
+        206.9263145487479
+        62.65064280055601
+        204.2898895284674
+          28.763888342342
+        60.38023879026305
+        204.2171110146289
+        8.116455861417121
+        29.02920871511511
+        62.45107640952574
+        201.0466193407952
+ 3.23e+10    
+         207.625635904509
+        63.01984219033692
+         204.930706775738
+        28.83199250891868
+        60.65310144662738
+        204.8595360601286
+        8.016581622099661
+        29.09829833780153
+        62.82035289677759
+        201.7365508816432
+ 3.24e+10    
+         208.326968855329
+        63.39000959152261
+        205.5723608810517
+        28.89946586142442
+        60.92618957467096
+        205.5028785892466
+        7.915622045814334
+        29.16675955212516
+        63.19061596541194
+         202.428547894642
+ 3.25e+10    
+        209.0303233306776
+        63.76115510256118
+        206.2148780706795
+        28.96630133383047
+        61.19951225953112
+        206.1471622899566
+        7.813565583421825
+        29.23458537173262
+         63.5618753927548
+        203.1226195107745
+ 3.26e+10    
+        209.7357092437941
+        64.13328885111849
+        206.8582846805763
+        29.03249184625397
+        61.47307851056993
+        206.7924109346145
+        7.710400597261291
+        29.30176879727084
+        63.93414098087424
+        203.8187748388462
+ 3.27e+10    
+        210.4431364897822
+        64.50642098740818
+         207.502607134645
+        29.09803030535525
+        61.74689725708586
+        207.4386483621671
+        7.606115365202957
+        29.36830281665062
+        64.30742255042182
+        204.5170229640303
+ 3.28e+10    
+        211.1526149437372
+        64.88056167764262
+         208.147871923427
+        29.16290960474098
+        62.02097734417105
+        208.0858984607077
+        7.500698084692567
+        29.43418040532008
+        64.68172993458887
+        205.2173729464446
+ 3.29e+10    
+        211.8641544589133
+        65.25572109761076
+         208.794105583227
+        29.22712262537739
+         62.2953275287151
+        208.7341851504065
+        7.394136876787375
+        29.49939452654827
+        65.05707297318227
+        205.9198338197515
+ 3.3e+10     
+        212.5777648649184
+        65.63190942638191
+        209.4413346757011
+        29.29066223601094
+        62.56995647555134
+        209.3835323668079
+        7.286419790182713
+        29.56393813171952
+        65.43346150681441
+        206.6244145897889
+ 3.31e+10    
+        213.2934559659471
+        66.00913684013604
+        210.0895857679128
+        29.35352129359453
+        62.84487275374913
+        210.0339640445206
+        7.177534805227531
+        29.62780416063773
+        65.81090537121098
+        207.3311242332239
+ 3.32e+10    
+        214.0112375390489
+        66.38741350612243
+        210.7388854128683
+        29.41569264372626
+        63.12008483304604
+        210.6855041012952
+        7.067469837929877
+        29.69098554184184
+        66.18941439163737
+        208.0399716962366
+ 3.33e+10    
+        214.7311193324304
+        66.76674957674692
+        211.3892601305504
+        29.47716912109285
+        63.39560108042307
+        211.3381764225007
+        6.956212743950202
+        29.75347519293298
+        66.56899837743975
+        208.7509658932321
+ 3.34e+10    
+        215.4531110637848
+        67.14715518378694
+        212.0407363894529
+        29.53794354992297
+        63.67142975681928
+        211.9920048460127
+         6.84375132258222
+        29.81526602091346
+        66.94966711670665
+        209.4641157055744
+ 3.35e+10    
+        216.1772224186711
+        67.52864043273688
+        212.6933405886274
+        29.59800874444974
+        63.94757901398491
+         212.647013147503
+        6.730073320721676
+        29.87635092253715
+        67.33143037104469
+        210.1794299803559
+ 3.36e+10    
+        216.9034630489144
+        67.91121539728211
+         213.347099040252
+        29.65735750937991
+        64.22405689147274
+        213.3032250261602
+        6.615166436819898
+        29.93672278467076
+        67.71429787047353
+        210.8969175291863
+ 3.37e+10    
+         217.631842571045
+        68.29489011390189
+        214.0020379527254
+        29.71598264037214
+        64.50087131376451
+        213.9606640908144
+        6.499018324824526
+        29.99637448466921
+        68.09827930843562
+        211.6165871270143
+ 3.38e+10    
+        218.3623705647742
+        68.67967457660149
+        214.6581834142961
+        29.77387692452474
+        64.77803008753308
+        214.6193538464971
+         6.38161659810457
+        30.05529889076183
+        68.48338433692315
+        212.3384475109743
+ 3.39e+10    
+        219.0950565715006
+        69.06557873177479
+        215.3155613772251
+         29.8310331408719
+        65.05554089903586
+        215.2793176814227
+        6.262948833360211
+        30.11348886245107
+        68.86962256172031
+        213.0625073792548
+ 3.4e+10     
+        219.8299100928536
+        69.45261247319308
+        215.9741976424941
+         29.8874440608859
+        65.33341131164281
+        215.9405788544019
+         6.14300257451624
+        30.17093725092325
+        69.25700353776102
+        213.7887753900092
+ 3.41e+10    
+        220.5669405892679
+        69.84078563712409
+        216.6341178450524
+        29.94310244899077
+        65.61164876349032
+        216.6031604826767
+         6.02176533659917
+        30.22763689947201
+        69.64553676460014
+        214.5172601602762
+ 3.42e+10    
+        221.3061574785961
+        70.23010799757685
+        217.2953474396123
+        29.99800106308236
+        65.89026056526636
+        217.2670855301957
+        5.899224609596859
+        30.28358064393364
+        70.03523168199965
+        215.2479702649344
+ 3.43e+10    
+        222.0475701347503
+        70.62058926167562
+        217.9579116869902
+        30.05213265505709
+        66.16925389812046
+        217.9323767963125
+        5.775367862300222
+        30.33876131313544
+        70.42609766562703
+        215.9809142356879
+ 3.44e+10    
+        222.7911878863804
+        71.01223906515766
+         218.621835640991
+        30.10548997135032
+        66.44863581169882
+        218.5990569049174
+        5.650182546127064
+        30.39317172935487
+        70.81814402286643
+        216.7161005600714
+ 3.45e+10    
+        223.5370200155839
+        71.40506696799838
+        219.2871441358392
+        30.15806575347828
+        66.72841322230084
+        219.2671482939908
+        5.523656098926097
+        30.44680470879118
+        71.21137998873948
+        217.4535376804848
+ 3.46e+10    
+        224.2850757566504
+        71.79908245015912
+        219.9538617741516
+        30.20985273859377
+         67.0085929111585
+         219.936673205596
+        5.395775948762756
+        30.49965306205063
+        71.60581472193894
+        218.1932339932543
+ 3.47e+10    
+        225.0353642948405
+        72.19429490746023
+        220.6220129154527
+        30.26084366004496
+        67.28918152283256
+        220.6076536762832
+        5.266529517683939
+         30.5517095946399
+        72.00145730096882
+        218.9351978477185
+ 3.48e+10    
+        225.7878947651903
+        72.59071364757381
+        221.2916216652231
+        30.31103124794302
+        67.57018556372607
+        221.2801115279196
+        5.135904225462923
+        30.60296710747478
+        72.39831672039406
+         219.679437545342
+ 3.49e+10    
+        226.5426762513572
+        72.98834788614003
+        221.9627118644833
+        30.36040822973777
+        67.85161140071295
+        221.9540683589437
+        5.003887493323145
+        30.65341839739758
+        72.79640188719807
+         220.425961338853
+ 3.5e+10     
+        227.2997177844933
+        73.38720674300127
+        222.6353070799038
+        30.40896733080009
+        68.13346525987897
+        222.6295455360249
+        4.870466747640688
+        30.70305625770679
+        73.19572161724361
+        221.1747774314075
+ 3.51e+10    
+        228.0590283421512
+        73.78729923855607
+        223.3094305944428
+        30.45670127501069
+        68.41575322537282
+        223.3065641861385
+         4.73562942362469
+        30.75187347869772
+        73.59628463184032
+         221.925893975778
+ 3.52e+10    
+        228.8206168472207
+        74.18863429022883
+        223.9851053984907
+        30.50360278535587
+        68.69848123836577
+        223.9851451890476
+         4.59936296897545
+        30.79986284821291
+        73.99809955441533
+         222.679319073569
+ 3.53e+10    
+        229.5844921668999
+        74.59122070905536
+        224.6623541815354
+        30.54966458452888
+        68.98165509611732
+        224.6653091701825
+        4.461654847519505
+        30.84701715220377
+        74.40117490728463
+        223.4350607744551
+ 3.54e+10    
+        230.3506631116958
+        74.99506719638357
+        225.3411993243243
+        30.59487939554018
+        69.26528045114487
+        225.3470764939192
+        4.322492542822022
+        30.89332917530174
+        74.80551910852705
+        224.1931270754458
+ 3.55e+10    
+        231.1191384344535
+        75.40018234068465
+        226.0216628915202
+        30.63923994232982
+        69.54936281049461
+        226.0304672572431
+        4.181863561774488
+        30.93879170139886
+        75.21114046895542
+        224.9535259201735
+ 3.56e+10    
+        231.8899268294178
+        75.80657461447632
+        226.7037666248542
+        30.68273895038821
+        69.83390753511273
+        226.7155012838043
+        4.039755438159029
+        30.98339751423838
+        75.61804718918788
+         225.716265198206
+ 3.57e+10    
+        232.6630369313287
+        76.21425237135483
+        227.3875319367434
+        30.72536914738153
+        70.11891983931268
+        227.4021981183452
+        3.896155736187687
+        31.02713939801425
+         76.0262473568134
+        226.4813527443829
+ 3.58e+10    
+        233.4384773145396
+        76.62322384313421
+        228.0729799043905
+        30.76712326378105
+        70.40440479033725
+        228.0905770214972
+         3.75105205401675
+        31.07001013797786
+        76.43574894365487
+        227.2487963381759
+ 3.59e+10    
+        234.2162564921721
+        77.03349713709176
+        228.7601312643384
+        30.80799403349994
+         70.6903673080145
+        228.7806569649513
+        3.604432027235699
+        31.11200252105596
+        76.84655980312311
+        228.0186037030737
+ 3.6e+10     
+        234.9963829152943
+        77.44508023331561
+        229.4490064074775
+        30.84797419453176
+        70.97681216450235
+        229.4724566269756
+        3.456283332330248
+        31.15310933647398
+        77.25868766766564
+        228.7907825059864
+ 3.61e+10    
+        235.7788649721305
+        77.85798098215793
+        230.1396253744943
+        30.88705648959522
+        71.26374398412165
+        230.1659943882913
+        3.306593690118946
+        31.19332337638676
+        77.67214014630369
+        229.5653403566783
+ 3.62e+10    
+        236.5637109873028
+        78.27220710178396
+        230.8320078517512
+        30.92523366678045
+        71.55116724327495
+        230.8612883282869
+        3.155350869163064
+        31.23263743651886
+        78.08692472225994
+        230.3422848072177
+ 3.63e+10    
+        237.3509292210958
+         78.6877661758229
+        231.5261731675886
+        30.96249848020281
+        71.83908627044846
+        231.5583562215708
+        3.002542689149756
+        31.27104431680829
+        78.50304875067303
+        231.1216233514528
+ 3.64e+10    
+        238.1405278687504
+        79.10466565111331
+        232.2221402890344
+        30.99884369065546
+        72.12750524629459
+        232.2572155348494
+        2.848157024247367
+         31.3085368220597
+        78.92051945639818
+          231.90336342451
+ 3.65e+10    
+        238.9325150597923
+        79.52291283554493
+        232.9199278189163
+        31.03426206626905
+        72.41642820379371
+        232.9578834241263
+        2.692181806433165
+        31.34510776260069
+        79.33934393189256
+        232.6875124023122
+ 3.66e+10    
+        239.7268988573705
+         79.9425148959909
+        233.6195539933625
+        31.06874638317038
+         72.7058590284915
+        233.6603767322148
+        2.534605028792281
+        31.38074995494571
+        79.75952913518316
+        233.4740776011152
+ 3.67e+10    
+        240.5236872576484
+        80.36347885633337
+        234.3210366796794
+        31.10228942614589
+        72.99580145881112
+        234.3647119865537
+        2.375414748788774
+         31.4154562224634
+        80.18108188791712
+        234.2630662770767
+ 3.68e+10    
+        241.3228881891951
+        80.78581159557629
+        235.0243933745948
+        31.13488398930662
+         73.2862590864362
+        235.0709053973151
+        2.214599091507058
+         31.4492193960491
+        80.60400887348979
+        235.0544856258333
+ 3.69e+10    
+         242.124509512421
+        81.20951984604609
+        235.7296412028628
+        31.16652287675419
+        73.57723535676456
+        235.7789728558095
+        2.052146252864386
+        31.48203231480225
+        81.02831663525376
+        235.8483427821064
+ 3.7e+10     
+        242.9285590190358
+        81.63461019167809
+        236.4367969162057
+        31.19719890324959
+        73.86873356942762
+        236.4889299331585
+        1.888044502793328
+        31.51388782670608
+        81.45401157480202
+        236.6446448193253
+ 3.71e+10    
+        243.7350444315225
+        82.06108906638374
+        237.1458768925941
+        31.22690489488042
+        74.16075687887599
+        237.2007918792491
+        1.722282188394042
+        31.54477878931156
+         81.8810999503286
+        237.4433987492719
+ 3.72e+10    
+        244.5439734026509
+        82.48896275250341
+        237.8568971358483
+        31.25563368973162
+        74.45330829502751
+        237.9145736219459
+        1.554847737056723
+        31.57469807042451
+        82.30958787506135
+        238.2446115217445
+ 3.73e+10    
+        245.3553535150052
+        82.91823737933468
+        238.5698732755482
+        31.28337813855605
+        74.74639068397602
+        238.6302897665614
+        1.385729659552396
+        31.60363854879369
+        82.73948131576734
+        239.0482900242407
+ 3.74e+10    
+        246.1691922805423
+        83.34891892174115
+         239.284820567249
+         31.3101311054428
+        75.04000676875751
+        239.3479545955665
+        1.214916553092997
+        31.63159311480216
+        83.17078609132882
+        239.8544410816615
+ 3.75e+10    
+        246.9854971401686
+        83.78101319883484
+        240.0017538929772
+        31.33588546848933
+        75.33415913017478
+        240.0675820685514
+        1.042397104360183
+        31.65855467116026
+        83.60350787138954
+        240.6630714560314
+ 3.76e+10    
+        247.8042754633494
+        84.21452587273494
+        240.7206877620117
+         31.3606341204686
+        75.62885020767422
+        240.7891858224048
+       0.8681600925016015
+        31.68451613359903
+         84.0376521750664
+        241.4741878462416
+ 3.77e+10    
+        248.6255345477311
+          84.649462447397
+        241.4416363119294
+        31.38436996949953
+        75.92408230027559
+        241.5127791717218
+       0.6921943920955718
+        31.70947043156419
+        84.47322436972917
+        242.2877968878059
+ 3.78e+10    
+        249.4492816187941
+        85.08582826751264
+        242.1646133099025
+        31.40708593971289
+        76.21985756755149
+        242.2383751094228
+       0.5144889760829336
+        31.73341050891194
+        84.91022966984332
+        243.1039051526391
+ 3.79e+10    
+        250.2755238295279
+        85.52362851748056
+        242.8896321542491
+         31.4287749719181
+        76.51617803065605
+        242.9659863075868
+       0.3350329186661929
+        31.75632932460286
+        85.34867313587921
+         243.922519148855
+ 3.8e+10     
+        251.1042682601251
+        85.96286822043901
+        243.6167058762096
+        31.44943002426672
+        76.81304557339777
+        243.6956251184701
+       0.1538153981751664
+         31.7782198533959
+        85.78855967327929
+        244.7436453205756
+ 3.81e+10    
+         251.935521917699
+        86.40355223736951
+        244.3458471419558
+        31.46904407291494
+         77.1104619433584
+        244.4273035757269
+      -0.0291743001004825
+        31.79907508654294
+        86.22989403148773
+        245.5672900477594
+ 3.82e+10    
+        252.7692917360246
+        86.84568526625949
+        245.0770682548053
+        31.48761011268294
+        77.40842875305248
+         245.161033395806
+      -0.2139467811129121
+        31.81888803247939
+        86.67268080304001
+        246.3934596460554
+ 3.83e+10    
+        253.6055845753004
+        87.28927184132989
+        245.8103811576468
+        31.50512115771255
+        77.70694748112814
+        245.8968259795251
+      -0.4005125372918066
+        31.83765171751536
+        87.11692442270753
+        247.2221603666593
+ 3.84e+10    
+        254.4444072219295
+         87.7343163323204
+         246.545797435556
+        31.52157024212005
+        78.00601947360627
+        246.6346924138147
+      -0.5888819458147658
+        31.85535918652372
+        87.56262916670117
+        248.0533983961977
+ 3.85e+10    
+        255.2857663883204
+        88.18082294383403
+        247.2833283185925
+        31.53695042064806
+        78.30564594515604
+        247.3746434736186
+      -0.7790652659122763
+        31.87200350362597
+         88.0097991519292
+        248.8871798566252
+ 3.86e+10    
+        256.1296687127179
+        88.62879571474167
+        248.0229846847787
+        31.55125476931275
+        78.60582798040512
+        248.1166896239494
+      -0.9710726362078583
+        31.88757775287566
+        88.45843833530726
+        249.7235108051336
+ 3.87e+10    
+         256.976120759039
+        89.07823851763547
+        248.7647770632338
+        31.56447638604731
+        78.90656653528393
+        248.8608410220899
+       -1.164914072094041
+        31.90207503893789
+        88.90855051312383
+        250.5623972340818
+ 3.88e+10    
+        257.8251290167382
+        89.52915505834272
+        249.5087156374739
+        31.57660839134129
+        79.20786243840097
+        249.6071075199338
+       -1.360599463143562
+        31.91548848776621
+        89.36013932045404
+          251.40384507094
+ 3.89e+10    
+        258.6766999006946
+          89.981548875489
+        250.2548102488506
+        31.58764392887607
+        79.50971639244727
+        250.3554986664567
+       -1.558138570557325
+        31.92781124727479
+         89.8132082306244
+        252.2478601782457
+ 3.9e+10     
+        259.5308397511048
+        90.43542334011191
+        251.0030704001299
+         31.5975761661557
+        79.81212897562988
+        251.1060237103136
+       -1.757541024648029
+        31.93903648800779
+        90.26776055472745
+        253.0944483535789
+ 3.91e+10    
+        260.3875548334134
+        90.89078165532568
+        251.7535052592024
+        31.60639829513265
+        80.11510064313173
+        251.8586916025545
+       -1.958816322361045
+         31.9491574038026
+        90.72379944118283
+        253.9436153295486
+ 3.92e+10    
+        261.2468513382445
+        91.34762685603266
+        252.5061236629119
+        31.61410353282851
+        80.41863172859674
+        252.6135109994535
+       -2.161973824832247
+         31.9581672124493
+        91.18132787534448
+        254.7953667737964
+ 3.93e+10    
+        262.1087353813628
+        91.80596180868345
+        253.2609341210004
+        31.62068512194996
+        80.72272244563806
+        253.3704902654411
+       -2.367022754982916
+        31.96605915634483
+        91.64034867915365
+        255.6497082890114
+ 3.94e+10    
+        262.9732130036465
+        92.26578921108016
+        254.0179448201526
+         31.6261363314988
+        81.02737288936916
+        254.1296374761408
+       -2.573972195152447
+        31.97282650314219
+        92.10086451083662
+        256.5066454129601
+ 3.95e+10    
+        263.8402901710795
+        92.72711159222429
+        254.7771636281406
+        31.63045045737606
+        81.33258303795414
+        254.8909604214899
+       -2.782831084769119
+        31.97846254639243
+        92.56287786464419
+        257.3661836185307
+ 3.96e+10    
+        264.7099727747628
+        93.18993131221001
+        255.5385980980615
+        31.63362082298027
+        81.63835275417978
+        255.6544666089609
+       -2.993608218058726
+        31.98296060618316
+        93.02639107063457
+         258.228328313788
+ 3.97e+10    
+        265.5822666309396
+        93.65425056215597
+         256.302255472652
+         31.6356407798007
+        81.94468178704341
+        256.4201632668572
+       -3.206312241792096
+        31.98631402976806
+        93.49140629449644
+        259.0930848420472
+ 3.98e+10    
+        266.4571774810368
+        94.12007136417834
+        257.0681426886811
+        31.63650370800215
+        82.25156977335843
+        257.1880573476832
+       -3.420951653071245
+         31.9885161921921
+         93.9579255374116
+        259.9604584819493
+ 3.99e+10    
+        267.3347109917268
+        94.58739557140406
+          257.83626638141
+        31.63620301700472
+         82.5590162393749
+        257.9581555315919
+       -3.637534797154572
+          31.989560496909
+         94.4259506359584
+        260.8304544475637
+ 4e+10       
+         268.214872755001
+        95.05622486802264
+        258.6066328891186
+        31.63473214605654
+         82.8670206024149
+        258.7304642298955
+       -3.856069865321685
+        31.98944037639193
+        94.89548326205087
+        261.7030778884899
+ 4.01e+10    
+        269.0976682882606
+         95.5265607693723
+        259.3792482576826
+        31.63208456479922
+        83.17558217252014
+        259.5049895886349
+       -4.076564892777785
+        31.98814929273624
+        95.36652492291688
+        262.5783338899797
+ 4.02e+10    
+        269.9831030344237
+        95.99840462206613
+        260.1541182452013
+        31.62825377382623
+        83.48470015411178
+        260.2817374922079
+       -4.299027756597847
+        31.98568073825682
+        95.83907696111116
+        263.4562274730662
+ 4.03e+10    
+        270.8711823620451
+        96.47175760414949
+        260.9312483266731
+        31.62323330523434
+        83.79437364766137
+        261.0607135670489
+       -4.523466173711613
+        31.98202823607476
+          96.313140554565
+        264.3367635947093
+ 4.04e+10    
+        271.7619115654539
+        96.94662072529417
+        261.7106436987027
+        31.61701672316737
+        84.10460165137056
+        261.8419231853498
+       -4.749887698928271
+        31.97718534069898
+        96.78871671666901
+        265.2199471479456
+ 4.05e+10    
+        272.6552958649012
+        97.42299482702423
+        262.4923092842495
+        31.60959762435194
+        84.41538306286081
+        262.6253714688317
+       -4.978299723002896
+        31.97114563859827
+        97.26580629639048
+        266.1057829620574
+ 4.06e+10    
+        273.5513404067286
+        97.90088058297481
+        263.2762497373931
+         31.6009696386264
+        84.72671668086851
+        263.4110632925438
+        -5.20870947074325
+        31.96390274876509
+        97.74440997842292
+        266.9942758027453
+ 4.07e+10    
+        274.4500502635433
+        98.38027849917994
+         264.062469448129
+        31.59112642946027
+        85.03860120694918
+        264.1990032887052
+       -5.441123999158607
+        31.95545032327102
+        98.22452828336868
+         267.885430372317
+ 4.08e+10    
+        275.3514304344152
+        98.86118891439513
+        264.8509725471821
+        31.58006169446751
+        85.35103524718627
+         264.989195850571
+       -5.675550195649375
+        31.94578204781448
+        98.70616156795134
+         268.779251309883
+ 4.09e+10    
+        276.2554858450757
+        99.34361200044411
+        265.6417629108234
+        31.56776916591022
+        85.66401731390432
+        265.7816451363238
+       -5.911994776239628
+        31.93489164225834
+        99.18931002525991
+        269.6757431915649
+ 4.1e+10     
+        277.1622213481438
+        99.82754776259941
+         266.434844165712
+        31.55424261119428
+        85.97754582738692
+        266.5763550729901
+       -6.150464283851173
+        31.92277286115963
+        99.67397368502222
+         270.574910530711
+ 4.11e+10    
+        278.0716417233529
+        100.3129960399868
+        267.2302196937226
+        31.53947583335629
+        86.29161911759759
+        267.3733293603725
+       -6.390965086620166
+          31.909419494289
+        100.1601524139079
+        271.4767577781244
+ 4.12e+10    
+        278.9837516777985
+        100.7999565060189
+        268.0278926367881
+        31.52346267154319
+        86.60623542590224
+        268.1725714749964
+       -6.633503376256819
+        31.89482536714222
+        100.6478459158593
+        272.3812893222977
+ 4.13e+10    
+        279.8985558461934
+        101.2884286688555
+        268.8278659017302
+        31.50619700148076
+        86.92139290679451
+        268.9740846740712
+       -6.878085166447556
+        31.87898434144162
+        101.1370537324507
+        273.2885094896646
+ 4.14e+10    
+        280.8160587911359
+        101.7784118718889
+         269.630142165087
+        31.48767273593626
+        87.23708962962058
+        269.7778719994551
+       -7.124716291300991
+        31.86189031562775
+        101.6277752432737
+        274.1984225448451
+ 4.15e+10    
+        281.7362650033946
+        102.2699052942543
+        270.4347238779267
+        31.46788382516941
+        87.55332358030502
+        270.5839362816302
+       -7.373402403836782
+        31.84353722534213
+        102.1200096663512
+        275.1110326909182
+ 4.16e+10    
+        282.6591789021961
+        102.7629079513655
+        271.2416132706503
+        31.44682425737638
+        87.87009266307589
+        271.3922801436761
+        -7.62414897451881
+         31.8239190438997
+        102.6137560585758
+        276.0263440696918
+ 4.17e+10    
+        283.5848048355327
+        103.2574186954741
+        272.0508123577773
+        31.42448805912289
+        88.18739470218783
+         272.202906005244
+       -7.876961289832162
+        31.80302978275192
+        103.1090133161735
+        276.9443607619837
+ 4.18e+10    
+        284.5131470804765
+        103.7534362162503
+        272.8623229427043
+        31.40086929576991
+        88.50522744364453
+         273.015816086531
+        -8.13184445090419
+        31.78086349193894
+        103.6057801751932
+        277.8650867879109
+ 4.19e+10    
+         285.444209843503
+        104.2509590413901
+        273.6761466224509
+        31.37596207188868
+        88.82358855691754
+        273.8310124122406
+       -8.388803372170379
+        31.75741426053305
+        104.1040552120201
+        278.7885261071879
+ 4.2e+10     
+         286.377997260834
+        104.7499855372407
+        274.4922847923747
+        31.34976053166714
+        89.14247563666338
+        274.6484968155471
+       -8.647842780084606
+        31.73267621707127
+        104.6038368439138
+        279.7146826194363
+ 4.21e+10    
+        287.3145133987798
+        105.2505139094517
+        275.3107386508576
+        31.32225885930645
+        89.46188620443564
+        275.4682709420373
+        -8.90896721187489
+        31.70664352997722
+        105.1051233295679
+        280.6435601644922
+ 4.22e+10    
+        288.2537622540974
+        105.7525422036419
+        276.1315092039621
+          31.293451279408
+        89.78181771039419
+        276.2903362536474
+       -9.172181014343902
+         31.6793104079742
+        105.6079127696947
+        281.5751625227335
+ 4.23e+10    
+        289.1957477543605
+        106.2560683060928
+        276.9545972700571
+         31.2633320573514
+        90.10226753500928
+        277.1146940325841
+       -9.437488342714982
+        31.65067110048631
+        106.1122031076306
+        282.5094934154062
+ 4.24e+10    
+        290.1404737583381
+        106.7610899444592
+        277.7800034844102
+        31.23189549966251
+        90.42323299076075
+        277.9413453852268
+       -9.704893159524136
+        31.62071989803022
+        106.6179921299651
+        283.4465565049624
+ 4.25e+10    
+        291.0879440563775
+        107.2676046884987
+        278.6077283037346
+        31.19913595437108
+         90.7447113238312
+        278.7702912460129
+       -9.974399233557726
+        31.58945113259607
+          107.12527746719
+        284.3863553954013
+ 4.26e+10    
+        292.0381623708057
+        107.7756099508235
+        279.4377720107119
+        31.16504781136011
+        91.06669971579478
+         279.601532381303
+       -10.24601013883613
+        31.55685917801793
+        107.6340565943714
+         285.328893632625
+ 4.27e+10    
+        292.9911323563299
+        108.2851029876682
+        280.2701347184594
+        31.12962550270388
+         91.3891952852976
+        280.4350693932242
+       -10.51972925364428
+        31.52293845033346
+        108.1443268318403
+        286.2741747047904
+ 4.28e+10    
+        293.9468576004619
+        108.7960808996807
+        281.1048163749708
+        31.09286350299763
+         91.7121950897334
+        281.2709027234881
+        -10.7955597596079
+        31.48768340813352
+        108.6560853459065
+        287.2222020426762
+ 4.29e+10    
+        294.9053416239324
+        109.3085406327238
+        281.9418167674993
+          31.054756329676
+        92.03569612691086
+        282.1090326571874
+       -11.07350464081758
+        31.45108855290044
+          109.16932914959
+        288.1729790200549
+ 4.3e+10     
+        295.8665878811287
+        109.8224789787043
+        282.7811355269127
+        31.01529854332237
+        92.35969533671425
+        282.9494593265627
+       -11.35356668299886
+        31.41314842933671
+        109.6840551033751
+        289.1265089540687
+ 4.31e+10    
+        296.8305997605361
+        110.3378925764114
+        283.6227721319837
+        30.97448474796854
+        92.68418960275588
+        283.7921827147451
+       -11.63574847273003
+        31.37385762568108
+        110.2002599159802
+        290.0827951056119
+ 4.32e+10    
+        297.7973805851869
+        110.8547779123786
+        284.4667259136556
+        30.93230959138303
+         93.0091757540212
+        284.6372026594642
+       -11.92005239670727
+        31.33321077401622
+        110.7179401451503
+        291.0418406797225
+ 4.33e+10    
+        298.7669336131166
+        111.3731313217581
+         285.312996059239
+        30.88876776535187
+        93.33465056650527
+        285.4845188567367
+       -12.20648064105698
+        31.29120255056431
+        111.2370921984671
+        292.0036488259775
+ 4.34e+10    
+        299.7392620378333
+        111.8929489892153
+        286.1615816165768
+        30.84385400594626
+        93.66061076484044
+        286.3341308645103
+       -12.49503519069654
+        31.24782767597155
+        111.7577123341771
+        292.9682226388946
+ 4.35e+10    
+        300.7143689887868
+        112.4142269498382
+          287.01248149815
+         30.7975630937833
+        93.98705302391602
+        287.1860381062902
+        -12.7857178287422
+        31.20308091558335
+        112.2797966620385
+        293.9355651583366
+ 4.36e+10    
+        301.6922575318529
+        112.9369610900635
+          287.86569448514
+        30.74988985427463
+        94.31397397048818
+        288.0402398747179
+       -13.07853013596564
+        31.15695707970748
+        112.8033411441871
+        294.9056793699292
+ 4.37e+10    
+        302.6729306698223
+        113.4611471486191
+        288.7212192314337
+        30.70082915786547
+        94.64137018478057
+        288.8967353351303
+       -13.37347349029877
+        31.10945102386714
+        113.3283415960191
+        295.8785682054776
+ 4.38e+10    
+        303.6563913428945
+         113.986780717482
+        289.5790542675849
+        30.65037592026435
+        94.96923820207705
+        289.7555235290762
+       -13.67054906638679
+        31.06055764904288
+        113.8547936870905
+        296.8542345433847
+ 4.39e+10    
+        304.6426424291842
+        114.5138572428529
+        290.4391980047183
+        30.59852510266261
+        95.29757451430264
+           290.6166033778
+       -13.96975783518986
+         31.0102719019043
+        114.3826929420373
+        297.8326812090885
+ 4.4e+10     
+        305.6316867452256
+        115.0423720261444
+        291.3016487383844
+        30.54527171194266
+        95.62637557159594
+        291.4799736856867
+       -14.27110056363371
+        30.95858877503052
+        114.9120347415096
+        298.8139109754925
+ 4.41e+10    
+        306.6235270464985
+        115.5723202249875
+        292.1664046523633
+        30.49061080087794
+        95.95563778387179
+        292.3456331436798
+       -14.57457781430922
+        30.90550330712031
+         115.442814323124
+        299.7979265634027
+ 4.42e+10    
+        307.6181660279436
+        116.1036968542502
+        293.0334638224122
+        30.43453746832187
+        96.28535752237377
+        293.2135803326505
+       -14.88018994522078
+        30.85101058319125
+        115.9750267824327
+        300.7847306419723
+ 4.43e+10    
+        308.6156063245007
+        116.6364967870734
+        293.9028242199644
+        30.37704685938676
+        96.61553112121501
+        294.0838137267386
+       -15.18793710958416
+        30.79510573476845
+        116.5086670739102
+        301.7743258291553
+ 4.44e+10    
+        309.6158505116376
+        117.1707147559209
+        294.7744837157751
+        30.31813416561366
+        96.94615487891191
+        294.9563316966533
+       -15.49781925567351
+        30.73778394006278
+        117.0437300119547
+        302.7667146921514
+ 4.45e+10    
+        310.6189011058995
+        117.7063453536437
+        295.6484400835089
+        30.25779462513064
+        97.27722505990364
+        295.8311325129337
+       -15.80983612671807
+         30.6790404241379
+        117.5802102719079
+        303.7618997478718
+ 4.46e+10    
+         311.624760565458
+        118.2433830345606
+        296.5246910032839
+          30.196023522803
+        97.60873789606424
+        296.7082143491759
+       -16.12398726084819
+        30.61887045906732
+        118.1181023910891
+        304.7598834633955
+ 4.47e+10    
+        312.6334312906624
+        118.7818221155512
+        297.4032340651563
+        30.13281619037187
+        97.94068958820233
+        297.5875752852176
+       -16.44027199109133
+        30.55726936408077
+        118.6574007698473
+        305.7606682564414
+ 4.48e+10    
+        313.6449156246071
+        119.3216567771655
+         298.284066772554
+        30.06816800658435
+        98.27307630755074
+        298.4692133102865
+       -16.75868944541782
+        30.49423250569965
+        119.1980996726272
+        306.7642564958358
+ 4.49e+10    
+        314.6592158536927
+        119.8628810647456
+        299.1671865456564
+         30.0020743973122
+         98.6058941972457
+        299.3531263261095
+       -17.07923854683639
+        30.42975529786299
+        119.7401932290527
+        307.7706505019883
+ 4.5e+10     
+        315.6763342082067
+        120.4054888895656
+        300.0525907247306
+        29.93453083566261
+        98.93913937379497
+        300.2393121499841
+       -17.40191801353977
+         30.3638332020419
+        120.2836754350257
+        308.7798525473724
+ 4.51e+10    
+        316.6962728628936
+        120.9494740299797
+        300.9402765733989
+        29.86553284207729
+        99.27280792853433
+        301.1277685178073
+       -17.72672635910074
+        30.29646172734417
+        120.8285401538403
+        309.7918648570071
+ 4.52e+10    
+         317.719033937546
+        121.4948301325907
+        301.8302412818747
+        29.79507598442299
+        99.60689592907536
+        302.0184930870726
+       -18.05366189271787
+        30.22763643060861
+        121.3747811173117
+        310.8066896089469
+ 4.53e+10    
+        318.7446194975909
+        122.0415507134295
+        302.7224819701289
+        29.72315587807187
+        99.94139942073944
+        302.9114834398212
+       -18.38272271951194
+        30.15735291648913
+        121.9223919269235
+        311.8243289347712
+ 4.54e+10    
+        319.7730315546849
+        122.5896291591479
+        303.6169956910185
+        29.64976818597226
+        100.2763144279838
+        303.8067370855578
+       -18.71390674087233
+        30.08560683752834
+        122.4713660549856
+        312.8447849200799
+ 4.55e+10    
+         320.804272067315
+        123.1390587282281
+        304.5137794333575
+        29.57490861870949
+        100.6116369558142
+        304.7042514641294
+       -19.04721165485425
+        30.01239389422093
+        123.0216968458125
+          313.86805960499
+ 4.56e+10    
+        321.8383429414037
+        123.6898325522034
+        305.4128301249402
+        29.49857293455782
+        100.9473629911881
+        305.6040239485601
+       -19.38263495662592
+        29.93770983506796
+        123.5733775169134
+        314.8941549846434
+ 4.57e+10    
+        322.8752460309172
+        124.2419436368954
+        306.3141446355145
+        29.42075693952185
+        101.2834885044064
+         306.506051847855
+       -19.72017393896682
+        29.86155045661918
+        124.1264011601986
+        315.9230730097083
+ 4.58e+10    
+        323.9149831384844
+        124.7953848636633
+        307.2177197797039
+        29.34145648736903
+        101.6200094504948
+        307.4103324097595
+       -20.05982569281601
+        29.78391160350715
+        124.6807607432007
+        316.9548155868891
+ 4.59e+10    
+        324.9575560160121
+         125.350148990668
+         308.123552319887
+        29.26066747965282
+        101.9569217705731
+        308.3168628234852
+       -20.40158710787106
+        29.70478916847089
+        125.2364491103109
+        317.9893845794418
+ 4.6e+10     
+        326.0029663653137
+          125.90622865415
+          309.03163896902
+        29.17838586572577
+        102.2942213932146
+         309.225640222392
+       -20.74545487323799
+        29.62417909236907
+        125.7934589840313
+          319.02678180769
+ 4.61e+10    
+        327.0512158387336
+        126.4636163697207
+         309.941976393419
+         29.0946076427441
+        102.6319042357947
+        310.1366616866436
+       -21.09142547813126
+        29.54207736418413
+          126.35178296624
+        320.0670090495404
+ 4.62e+10    
+        328.1023060397873
+        127.0223045336686
+        310.8545612154913
+        29.00932885566202
+        102.9699662058277
+        311.0499242458114
+       -21.43949521262492
+        29.45848002101656
+         126.911413539474
+         321.110068041014
+ 4.63e+10    
+        329.1562385237949
+        127.5822854242777
+        311.7693900164198
+         28.9225455972179
+         103.308403202294
+        311.9654248814533
+       -21.78966016845371
+        29.37338314806896
+        127.4723430682228
+        322.1559604767639
+ 4.64e+10    
+        330.2130147985252
+        128.1435512031628
+        312.6864593388066
+        28.83425400791009
+        103.6472111169557
+         312.883160529653
+       -22.14191623986544
+        29.28678287862161
+        128.0345638002426
+        323.2046880106103
+ 4.65e+10    
+        331.2726363248408
+        128.7060939166143
+        313.6057656892658
+        28.74445027596455
+        103.9863858356615
+        313.8031280835161
+       -22.49625912452344
+         29.1986753939974
+        128.5980678678798
+        324.2562522560711
+ 4.66e+10    
+        332.3351045173547
+        129.2699054969619
+         314.527305540972
+        28.65313063729342
+        104.3259232396422
+        314.7253243956425
+       -22.85268432445988
+        29.10905692351778
+        129.1628472894122
+        325.3106547868983
+ 4.67e+10    
+        333.4004207450805
+        129.8349777639484
+        315.4510753361699
+        28.56029137544297
+        104.6658192067926
+        315.6497462805518
+       -23.21118714707943
+        29.01792374444982
+        129.7288939704052
+        326.3678971376174
+ 4.68e+10    
+        334.4685863320944
+        130.4013024261179
+        316.3770714886335
+        28.46592882153536
+         105.006069612947
+        316.5763905170789
+       -23.57176270621337
+        28.92527218194311
+        130.2961997050805
+        327.4279808040656
+ 4.69e+10    
+        335.5396025581987
+        130.9688710822208
+        317.3052903860904
+        28.37003935419923
+        105.3466703331409
+        317.5052538507386
+       -23.93440592322421
+        28.83109860895829
+        130.8647561777035
+        328.4909072439416
+ 4.7e+10     
+        336.6134706595888
+        131.5376752226296
+         318.235728392596
+        28.27261939949251
+        105.6876172428627
+        318.4363329960456
+       -24.29911152816071
+        28.73539944618559
+          131.43455496398
+         329.556677877352
+ 4.71e+10    
+        337.6901918295277
+        132.1077062307705
+        319.1683818508761
+        28.17366543081624
+         106.028906219298
+        319.3696246388105
+       -24.66587406096283
+        28.63817116195548
+        132.0055875324728
+        330.6252940873582
+ 4.72e+10    
+        338.7697672190164
+        132.6789553845677
+        320.1032470846158
+        28.07317396882007
+         106.370533142558
+        320.3051254383958
+       -25.03468787271732
+        28.53941027213929
+        132.5778452460308
+        331.6967572205356
+ 4.73e+10    
+        339.8521979374804
+        133.2514138579028
+        321.0403204007212
+        27.97114158129878
+         106.712493896904
+         321.242832029945
+       -25.40554712696308
+        28.43911334004149
+        133.1513193632319
+        332.7710685875263
+ 4.74e+10    
+        340.9374850534463
+        133.8250727220891
+         321.979598091537
+        27.86756488308042
+        107.0547843719568
+        322.1827410265697
+       -25.77844580104665
+        28.33727697628318
+        133.7260010398423
+        333.8482294635963
+ 4.75e+10    
+         342.025629595235
+        134.3999229473573
+        322.9210764370243
+        27.76244053590617
+        107.3974004638991
+        323.1248490215161
+        -26.1533776875274
+        28.23389783867695
+        134.3018813302906
+        334.9282410892055
+ 4.76e+10    
+        343.1166325516485
+        134.9759554043584
+        323.8647517068991
+         27.6557652483018
+        107.7403380766657
+        324.0691525902902
+       -26.53033639563305
+         28.1289726320926
+        134.8789511891548
+        336.0111046705642
+ 4.77e+10    
+        344.2104948726645
+        135.5531608656779
+        324.8106201627395
+         27.5475357754405
+        108.0835931231249
+        325.0156482927562
+       -26.90931535276363
+        28.02249810831518
+        135.4572014726666
+        337.0968213802046
+ 4.78e+10    
+        345.3072174701391
+        136.1315300073678
+         325.758678060053
+        27.43774891899856
+        108.4271615262512
+        325.9643326752058
+       -27.29030780604634
+        27.91447106589424
+        136.0366229402286
+          338.18539235755
+ 4.79e+10    
+         346.406801218502
+        136.7110534104885
+        326.7089216503075
+        27.32640152700148
+        108.7710392202854
+          326.91520227239
+       -27.67330682393877
+        27.80488834998435
+        136.6172062559466
+        339.2768187094886
+ 4.8e+10     
+        347.5092469554716
+        137.2917215626698
+        327.6613471829295
+        27.21349049366338
+        109.1152221518877
+        327.8682536095325
+       -28.05830529788152
+        27.69374685217801
+        137.1989419901778
+        340.3711015109494
+ 4.81e+10    
+        348.6145554827507
+         137.873524859682
+        328.6159509072637
+        27.09901275921767
+        109.4597062812794
+        328.8234832043022
+       -28.44529594399989
+        27.58104351033028
+         137.781820621093
+        341.4682418054786
+ 4.82e+10    
+        349.7227275667517
+        138.4564536070236
+         329.572729074506
+        26.98296530974024
+        109.8044875833761
+        329.7808875687628
+       -28.83427130485432
+        27.46677530837496
+        138.3658325362532
+        342.5682406058227
+ 4.83e+10    
+        350.8337639393068
+        139.0404980215238
+        330.5316779395979
+        26.86534517696486
+        110.1495620489113
+        330.7404632112953
+       -29.22522375123967
+        27.35093927613342
+        138.9509680342011
+        343.6710988945104
+ 4.84e+10    
+        351.9476652983877
+        139.6256482329579
+        331.4927937630918
+        26.74614943809084
+        110.4949256855509
+        331.7022066384918
+       -29.61814548403226
+        27.23353248911543
+        139.5372173260709
+        344.7768176244438
+ 4.85e+10    
+        353.0644323088312
+         140.211894285679
+        332.4560728129821
+         26.6253752155831
+        110.8405745189968
+        332.6661143570147
+       -30.01302853608578
+        27.11455206831171
+        140.1245705372061
+        345.8853977194796
+ 4.86e+10    
+        354.1840656030608
+         140.799226140262
+        333.4215113665082
+        26.50301967696489
+         111.186504594085
+        333.6321828754426
+       -30.40986477417488
+         26.9939951799796
+        140.7130177087988
+        346.9968400750287
+ 4.87e+10    
+        355.3065657818229
+        141.3876336751654
+        334.3891057119271
+        26.37908003460314
+        111.5327119758702
+        334.6004087060784
+       -30.80864590098643
+        26.87185903542088
+        141.3025487995417
+        348.1111455586447
+ 4.88e+10    
+         356.431933414916
+        141.9771066884041
+        335.3588521502535
+        26.25355354548625
+         111.879192750705
+        335.5707883667374
+       -31.20936345715832
+        26.74814089075194
+         141.893153687293
+        349.2283150106246
+ 4.89e+10    
+        357.5601690419283
+        142.5676348992407
+        336.3307469969757
+        26.12643751099499
+        112.2259430273076
+        336.5433183825074
+       -31.61200882336542
+        26.62283804666682
+        142.4848221707595
+        350.3483492446066
+ 4.9e+10     
+        358.6912731729783
+        143.1592079498872
+        337.3047865837422
+        25.99772927666618
+        112.5729589378238
+        337.5179952874861
+       -32.01657322245269
+        26.49594784819354
+        143.0775439711934
+        351.4712490481744
+ 4.91e+10    
+        359.8252462894582
+        143.7518154072274
+        338.2809672600166
+        25.86742623194937
+        112.9202366388766
+        338.4948156264929
+       -32.42304772161449
+        26.36746768444213
+        143.6713087341035
+        352.5970151834603
+ 4.92e+10    
+        360.9620888447803
+        144.3454467645462
+        339.2592853947123
+        25.73552580995674
+        113.2677723126108
+        339.4737759567579
+        -32.8314232346209
+        26.23739498834655
+        144.2661060309821
+        353.7256483877524
+ 4.93e+10    
+        362.1018012651289
+        144.9400914432837
+         340.239737377797
+        25.60202548720603
+         113.615562167726
+        340.4548728495844
+       -33.24169052408933
+        26.10572723639981
+        144.8619253610483
+        354.8571493741089
+ 4.94e+10    
+        363.2443839502089
+        145.5357387947935
+        341.2223196218725
+         25.4669227833566
+        113.9636024405039
+        341.4381028919939
+       -33.65384020380268
+        25.97246194838165
+        145.4587561530037
+        355.9915188319676
+ 4.95e+10    
+        364.3898372740113
+        146.1323781021249
+          342.20702856373
+        25.33021526093993
+        114.3118893958254
+        342.4234626883457
+       -34.06786274107207
+        25.83759668707984
+        146.0565877668061
+        357.1287574277603
+ 4.96e+10    
+        365.5381615855642
+        146.7299985818156
+        343.1938606658833
+        25.19190052508195
+        114.6604193281805
+        343.4109488619328
+       -34.48374845914575
+        25.70112905800498
+        146.6554094954553
+        358.2688658055372
+ 4.97e+10    
+        366.6893572096998
+        147.3285893856996
+        344.1828124180716
+        25.05197622322035
+        115.0091885626691
+        344.4005580565576
+       -34.90148753966121
+        25.56305670909905
+        147.2552105667986
+        359.4118445875827
+ 4.98e+10    
+        367.8434244478283
+        147.9281396027328
+        345.1738803387508
+        24.91044004481554
+        115.3581934559959
+        345.3922869380932
+        -35.3210700251433
+        25.42337733043708
+        147.8559801453462
+        360.5576943750416
+ 4.99e+10    
+        369.0003635786941
+        148.5286382608297
+        346.1670609765519
+        24.76728972105435
+        115.7074303974546
+        346.3861321960142
+       -35.74248582154519
+        25.28208865392303
+        148.4577073341069
+        361.7064157485453
+ 5e+10       
+        370.1601748591618
+        149.1300743287199
+        347.1623509117193
+        24.62252302454895
+        116.0568958099061
+        347.3820905449117
+       -36.16572470083322
+        25.13918845297915
+        149.0603811764348
+        362.8580092688415
+ 5.01e+10    
+        371.3228585249881
+        149.7324367178163
+        348.1597467575356
+        24.47613776902923
+        116.4065861507487
+        348.3801587259906
+       -36.59077630361537
+        24.99467454222985
+        149.6639906578948
+        364.0124754774262
+ 5.02e+10    
+           372.4884147916
+        150.3357142841002
+        349.1592451617196
+         24.3281318090291
+        116.7564979128802
+        349.3803335085474
+       -37.01763014181178
+         24.8485447771796
+        150.2685247081416
+        365.1698148971798
+ 5.03e+10    
+        373.6568438548827
+        150.9398958300212
+        350.1608428078022
+        24.17850303956799
+        117.1066276256532
+        350.3826116914264
+       -37.44627560136854
+        24.70079705388449
+        150.8739722028148
+        366.3300280330038
+ 5.04e+10    
+        374.8281458919645
+        151.5449701064128
+        351.1645364164865
+        24.02724939582554
+        117.4569718558218
+        351.3869901044606
+       -37.87670194501254
+         24.5514293086186
+         151.480321965448
+        367.4931153724602
+ 5.05e+10    
+        376.0023210620079
+        152.1509258144237
+        352.1703227469944
+        23.87436885281194
+        117.8075272084824
+        352.3934656098966
+       -38.30889831504854
+        24.40043951753538
+        152.0875627693962
+        368.6590773864195
+ 5.06e+10    
+        377.1793695070015
+        152.7577516074636
+        353.1781985983805
+        23.71985942503181
+        118.1582903280054
+        353.4020351037939
+       -38.74285373619684
+        24.24782569632222
+        152.6956833397757
+        369.8279145297032
+ 5.07e+10    
+        378.3592913525613
+        153.3654360931648
+        354.1881608108438
+        23.56371916614416
+        118.5092578989627
+        354.4126955174219
+       -39.17855711847183
+        24.09358589985133
+        153.3046723554219
+        370.9996272417344
+ 5.08e+10    
+        379.5420867087257
+        153.9739678353606
+        355.2002062670118
+        23.40594616861587
+        118.8604266470441
+        355.4254438186248
+       -39.61599726010022
+        23.93771822182426
+        153.9145184508611
+        372.1742159471918
+ 5.09e+10    
+        380.7277556707628
+        154.5833353560763
+        356.2143318932113
+        23.24653856337062
+        119.2117933399698
+        356.4402770131813
+       -40.05516285047961
+        23.78022079441207
+         154.525210218297
+        373.3516810566617
+ 5.1e+10     
+        381.9162983199824
+        155.1935271375405
+        357.2305346607229
+        23.08549451943384
+        119.5633547883956
+        357.4571921461464
+       -40.49604247317544
+        23.62109178789012
+        155.1367362096165
+           374.5320229673
+ 5.11e+10    
+        383.1077147245364
+        155.8045316242057
+        358.2488115870245
+        22.92281224357122
+        119.9151078468097
+        358.4761863031757
+       -40.93862460895684
+        23.46032941026881
+        155.7490849384076
+        375.7152420634913
+ 5.12e+10    
+        384.3020049402421
+        156.4163372247911
+        359.2691597370069
+        22.75848997992389
+         120.267049414424
+        359.4972566118338
+       -41.38289763887079
+        23.29793190691849
+        156.3622448819923
+        376.9013387175132
+ 5.13e+10    
+        385.4991690113972
+        157.0289323143362
+        360.2915762241909
+         22.5925260096388
+        120.6191764360594
+        360.5204002428985
+        -41.8288498473533
+        23.13389756019146
+        156.9762044834807
+        378.0903132902062
+ 5.14e+10    
+        386.6992069716004
+        157.6423052362725
+        361.3160582119146
+        22.42491865049386
+        120.9714859030227
+        361.5456144116358
+       -42.27646942537825
+        22.96822468903751
+        157.5909521538328
+        379.2821661316414
+ 5.15e+10    
+        387.9021188445793
+        158.2564443045111
+        362.3426029145228
+        22.25566625652026
+        121.3239748539783
+        362.5728963790767
+       -42.72574447364183
+        22.80091164861754
+        158.2064762739436
+        380.4768975817961
+ 5.16e+10    
+        389.1079046450161
+        158.8713378055433
+        363.3712075985255
+        22.08476721761936
+        121.6766403758132
+        363.6022434532657
+       -43.17666300578377
+        22.63195682991082
+        158.8227651967374
+        381.6745079712307
+ 5.17e+10    
+         390.316564379381
+         159.486974000562
+        364.4018695837622
+        21.91221995917628
+        122.0294796044967
+        364.6336529905157
+       -43.62921295164315
+        22.46135865931985
+        159.4398072492834
+        382.8749976217678
+ 5.18e+10    
+        391.5280980467682
+        160.1033411275928
+        365.4345862445346
+        21.73802294166907
+        122.3824897259312
+        365.6671223966275
+       -44.08338216054923
+         22.2891155982707
+        160.0575907349226
+        384.0783668471761
+ 5.19e+10    
+        392.7425056397364
+         160.720427403647
+        366.4693550107473
+        21.56217466027489
+        122.7356679768001
+        366.7026491281188
+       -44.53915840464627
+         22.1152261428093
+        160.6761039354139
+         385.284615953859
+ 5.2e+10     
+        393.9597871451487
+        161.3382210268851
+        367.5061733690171
+         21.3846736444716
+        123.0890116454073
+        367.7402306934269
+       -44.99652938225191
+        21.93968882319501
+        161.2953351130937
+        386.4937452415419
+ 5.21e+10    
+        395.1799425450245
+        161.9567101788004
+        368.5450388637889
+        21.20551845763665
+        123.4425180725121
+        368.7798646541081
+       -45.45548272124817
+        21.76250220348971
+        161.9152725130508
+        387.7057550039665
+ 5.22e+10    
+        396.4029718173851
+         162.575883026416
+        369.5859490984257
+        21.02470769664237
+        123.7961846521572
+        369.8215486260243
+         -45.916005982505
+        21.58366488114418
+        162.5359043653208
+        388.9206455295883
+ 5.23e+10    
+        397.6288749371122
+        163.1957277244987
+        370.6289017363032
+        20.84223999144756
+        124.1500088324922
+        370.8652802805159
+       -46.37808666333507
+        21.40317548658149
+        163.1572188870923
+         390.138417102275
+ 5.24e+10    
+        398.8576518768031
+        163.8162324177883
+        371.6738945018791
+        20.65811400468657
+        124.5039881165893
+        371.9110573455702
+       -46.84171220097984
+         21.2210326827762
+        163.7792042849305
+        391.3590700020134
+ 5.25e+10    
+        400.0893026076344
+        164.4373852432435
+        372.7209251817653
+        20.47232843125529
+        124.8581200632558
+        372.9588776069743
+       -47.30686997612519
+        21.03723516483227
+        164.4018487570165
+        392.5826045056133
+ 5.26e+10    
+        401.3238271002252
+         165.059174332303
+        373.7699916257821
+        20.28488199789419
+        125.2124022878393
+        374.0087389094634
+       -47.77354731644734
+        20.85178165955658
+        165.0251404954037
+        393.8090208874214
+ 5.27e+10    
+        402.5612253255127
+        165.6815878131642
+        374.8210917480137
+         20.0957734627686
+        125.5668324630279
+        375.0606391578575
+       -48.24173150018741
+         20.6646709250307
+        165.6490676882868
+        395.0383194200286
+ 5.28e+10    
+        403.8014972556179
+        166.3046138130752
+        375.8742235278417
+        19.90500161504671
+        125.9214083196449
+        376.1145763181873
+       -48.71140975975366
+        20.47590175018037
+        166.2736185222913
+        396.2705003749992
+ 5.29e+10    
+        405.0446428647294
+        166.9282404606443
+        376.9293850109809
+        19.71256527447442
+        126.2761276474384
+         377.170548418817
+       -49.18256928535197
+        20.28547295434156
+        166.8987811847738
+        397.5055640235812
+ 5.3e+10     
+        406.2906621299809
+        167.5524558881677
+        377.9865743105093
+         19.5184632909496
+        126.6309882958656
+        378.2285535515524
+       -49.65519722864215
+         20.0933833868255
+         167.524543866142
+         398.743510637439
+ 5.31e+10    
+          407.53955503234
+        168.1772482339678
+        379.0457896078766
+        19.32269454409192
+        126.9859881748715
+        379.2885898727479
+       -50.12928070642121
+        19.89963192648068
+        168.1508947621895
+        399.9843404893781
+ 5.32e+10    
+         408.791321557494
+         168.802605644754
+         380.107029153921
+        19.12525794281267
+        127.3411252556629
+        380.3506556044009
+       -50.60480680433094
+        19.70421748125353
+        168.7778220764451
+         401.228053854079
+ 5.33e+10    
+        410.0459616967455
+        169.4285162779931
+        381.1702912698711
+        18.92615242488112
+        127.6963975714768
+        381.4147490352345
+       -51.08176258059069
+        19.50713898774693
+        169.4053140225397
+        402.4746510088365
+ 5.34e+10    
+        411.3034754479115
+        170.0549683043017
+        382.2355743483431
+        18.72537695649088
+        128.0518032183443
+         382.480868521789
+       -51.56013506975349
+        19.30839541077711
+        170.0333588265882
+        403.7241322342936
+ 5.35e+10    
+        412.5638628162217
+        170.6819499098496
+        383.3028768543321
+        18.52293053182304
+        128.4073403558499
+        383.5490124894917
+       -52.03991128648523
+        19.10798574292927
+        170.6619447295878
+        404.9764978151917
+ 5.36e+10    
+        413.8271238152266
+        171.3094492987826
+        384.3721973261972
+        18.31881217260894
+        128.7630072078847
+        384.6191794337209
+       -52.52107822936577
+        18.90590900411178
+        171.2910599898315
+        406.2317480411157
+ 5.37e+10    
+        415.0932584677069
+          171.93745469566
+        385.4435343766411
+        18.11302092769109
+        129.1188020633958
+         385.691367920874
+       -53.00362288471214
+        18.70216424110868
+        171.9206928853372
+         407.489883207246
+ 5.38e+10    
+        416.3622668065858
+        172.5659543479069
+        386.5168866936845
+        17.90555587258347
+        129.4747232771312
+        386.7655765894206
+       -53.48753223042151
+        18.49675052713176
+        172.5508317162949
+         408.750903615116
+ 5.39e+10    
+        417.6341488758533
+        173.1949365282868
+        387.5922530416365
+        17.69641610903033
+        129.8307692703785
+        387.8418041509522
+       -53.97279323983432
+        18.28966696137125
+        173.1814648075257
+        410.0148095733713
+ 5.4e+10     
+        418.9089047314827
+        173.8243895373845
+        388.6696322620585
+        17.48560076456451
+        130.1869385317016
+        388.9200493912291
+       -54.45939288561625
+        18.08091266854626
+        173.8125805109612
+        411.2816013985323
+ 5.41e+10    
+        420.1865344423596
+        174.4543017061073
+        389.7490232747225
+        17.27310899206485
+        130.5432296176695
+        390.0003111712151
+       -54.94731814365852
+        17.87048679845353
+        174.4441672081344
+        412.5512794157647
+ 5.42e+10    
+        421.4670380912134
+        175.0846613982058
+        390.8304250785708
+        17.05893996931296
+         130.899641153584
+        391.0825884281155
+       -55.43655599699517
+        17.65838852551735
+        175.0762133126904
+        413.8238439596506
+ 5.43e+10    
+        422.7504157755565
+        175.7154570128042
+        391.9138367526654
+        16.84309289855009
+        131.2561718342005
+        392.1668801764088
+       -55.92709343973692
+        17.44461704833707
+        175.7087072729088
+        415.0992953749652
+ 5.44e+10    
+         424.036667608618
+        176.3466769869517
+        392.9992574571377
+        16.62556700603324
+        131.6128204244458
+        393.2531855088644
+       -56.41891748102066
+        17.22917158923651
+        176.3416375742457
+        416.3776340174557
+ 5.45e+10    
+        425.3257937202922
+        176.9783097981856
+        394.0866864341292
+        16.40636154159096
+        131.9695857601306
+        394.3415035975706
+       -56.91201514897368
+         17.0120513938119
+        176.9749927418895
+        417.6588602546312
+ 5.46e+10    
+        426.6177942580879
+        177.6103439671161
+         395.176123008742
+        16.18547577818033
+        132.3264667486594
+        395.4318336949481
+       -57.40637349469167
+         16.7932557304803
+        177.6087613433313
+        418.9429744665463
+ 5.47e+10    
+        427.9126693880817
+          178.24276806002
+        396.2675665899655
+        15.96290901144264
+        132.6834623697341
+        396.5241751347613
+       -57.90197959622942
+        16.57278389002871
+        178.2429319909536
+        420.2299770465964
+ 5.48e+10    
+        429.2104192958733
+        178.8755706914558
+        397.3610166716231
+        15.73866055926042
+        133.0405716760551
+          397.61852733313
+       -58.39882056260461
+        16.35063518516273
+        178.8774933446327
+         421.519868402318
+ 5.49e+10    
+         430.511044187551
+        179.5087405268916
+        398.4564728332966
+        15.51272976131452
+        133.3977937940172
+        398.7148897895348
+       -58.89688353781131
+        16.12680895005697
+        179.5124341143576
+        422.8126489561872
+ 5.5e+10     
+        431.8145442906603
+        180.1422662853503
+        399.5539347412645
+        15.28511597864243
+        133.7551279244034
+        399.8132620878154
+        -59.3961557048452
+        15.90130453990504
+        180.1477430628652
+        424.1083191464297
+ 5.51e+10    
+        433.1209198551705
+        180.7761367420692
+         400.653402149422
+        15.05581859319637
+        134.1125733430711
+        400.9136438971748
+        -59.8966242897373
+        15.67412133047095
+        180.7834090082883
+        425.4068794278294
+ 5.52e+10    
+        434.4301711544556
+        181.4103407311774
+        401.7548749002153
+        14.82483700740327
+        134.4701294016395
+        402.0160349731729
+       -60.39827656559653
+        15.44525871764155
+        181.4194208268227
+         426.708330272544
+ 5.53e+10    
+        435.7422984862741
+        182.0448671483862
+        402.8583529255605
+         14.5921706437253
+        134.8277955281675
+         403.120435158721
+       -60.90109985665958
+        15.21471611697995
+        182.0557674554079
+        428.0126721709286
+ 5.54e+10    
+        437.0573021737544
+        182.6797049536982
+        403.9638362477708
+        14.35781894422185
+        135.1855712278332
+         404.226844385072
+       -61.40508154234807
+        14.98249296328052
+        182.6924378944234
+        429.3199056323568
+ 5.55e+10    
+        438.3751825663863
+        183.3148431741292
+        405.0713249804755
+          14.121781370113
+         135.543456083605
+        405.3352626728073
+       -61.91020906133042
+        14.74858871012508
+        183.3294212103993
+        430.6300311860493
+ 5.56e+10    
+        439.6959400410145
+        183.9502709064476
+          406.18081932954
+        13.88405740134439
+        135.9014497569123
+        406.4456901328288
+       -62.41646991558932
+        14.51300282944087
+        183.9667065387472
+        431.9430493819112
+ 5.57e+10    
+        441.0195750028403
+        184.5859773199295
+        407.2923195939874
+        13.64464653615391
+        136.2595519883116
+        407.5581269673372
+       -62.92385167449277
+        14.27573481106032
+        184.6042830864988
+        433.2589607913697
+ 5.58e+10    
+        442.3460878864276
+        185.2219516591262
+        408.4058261669126
+        13.40354829063985
+        136.6177625981473
+        408.6725734708156
+       -63.43234197886785
+        14.03678416228252
+        185.2421401350666
+         434.577766008214
+ 5.59e+10    
+         443.675479156708
+        185.8581832466531
+        409.5213395364051
+         13.1607621983317
+        136.9760814872115
+         409.789030031015
+       -63.94192854507667
+        13.79615040743752
+        185.8802670430171
+        435.8994656494476
+ 5.6e+10     
+         445.007749310001
+        186.4946614859866
+        410.6388602864602
+        12.91628780976296
+        137.3345086373994
+        410.9074971299265
+       -64.45259916909296
+        13.55383308745163
+         186.518653248858
+        437.2240603561378
+ 5.61e+10    
+        446.3428988750293
+        187.1313758642845
+        411.7583890978988
+        12.67012469204549
+        137.6930441123594
+         412.027975344763
+       -64.96434173057928
+        13.30983175941598
+        187.1572882738423
+        438.5515507942731
+ 5.62e+10    
+        447.6809284139449
+         187.768315955214
+        412.8799267492841
+        12.42227242844783
+        138.0516880581442
+        413.1504653489371
+       -65.47714419696243
+        13.06414599615811
+         187.796161724789
+        439.8819376556281
+ 5.63e+10    
+        449.0218385233585
+        188.4054714217997
+          414.00347411783
+        12.17273061797425
+        138.4104407038527
+        414.2749679130333
+        -65.9909946275077
+        12.81677538581464
+        188.4352632969158
+        441.2152216586301
+ 5.64e+10    
+        450.3656298353725
+         189.042832019287
+        415.1290321803269
+        11.92149887494858
+        138.7693023622731
+        415.4014839057806
+       -66.50588117738951
+        12.56771953140841
+         189.074582776687
+        442.5514035492249
+ 5.65e+10    
+        451.7123030186205
+        189.6803875980168
+         416.256602014049
+        11.66857682859925
+        139.1282734305214
+        416.5300142950313
+         -67.021792101759
+        12.31697805042781
+          189.71411004468
+        443.8904841017634
+ 5.66e+10    
+        453.0618587793139
+        190.3181281063205
+         417.386184797676
+        11.41396412264843
+        139.4873543906763
+        417.6605601487319
+       -67.53871575980634
+        12.06455057440919
+        190.3538350784623
+        445.2324641198725
+ 5.67e+10    
+        454.4142978622866
+        190.9560435934254
+        418.5177818122031
+        11.15766041490411
+        139.8465458104103
+        418.7931226358913
+       -68.05664061881663
+        11.81043674852319
+        190.9937479554871
+        446.5773444373514
+ 5.68e+10    
+        455.7696210520524
+        191.5941242123784
+        419.6513944418646
+        10.89966537685533
+        140.2058483436192
+        419.9277030275559
+       -68.57555525821999
+        11.55463623116403
+        191.6338388560002
+        447.9251259190549
+ 5.69e+10    
+        457.1278291738632
+        192.2323602229828
+        420.7870241750439
+        10.63997869327179
+        140.5652627310478
+        421.0643026977799
+       -69.09544837363313
+        11.29714869354222
+         192.274098065964
+        449.2758094617943
+ 5.7e+10     
+        458.4889230947733
+        192.8707419947503
+        421.9246726051946
+        10.37860006180551
+        140.9247898009114
+         422.202923124598
+       -69.61630878089247
+         11.0379738192822
+        192.9145159799981
+        450.6293959952396
+ 5.71e+10    
+        459.8529037247094
+        193.5092600098683
+        423.0643414317594
+        10.11552919259838
+        141.2844304695163
+        423.3435658909891
+       -70.13812542007737
+        10.77711130402177
+        193.5550831043262
+        451.9858864828176
+ 5.72e+10    
+        461.2197720175419
+        194.1479048661818
+         424.206032461085
+        9.850765807891845
+        141.6441857418756
+        424.4862326858558
+       -70.66088735952211
+        10.51456085501803
+        194.1957900597497
+         453.345281922635
+ 5.73e+10    
+         462.589528972168
+        194.7866672801903
+        425.3497476073479
+        9.584309641642015
+        142.0040567123231
+        425.6309253049894
+       -71.18458379981669
+        10.25032219075604
+        194.8366275846262
+        454.7075833483852
+ 5.74e+10    
+        463.9621756335961
+        195.4255380900573
+        426.4954888934695
+         9.31616043913861
+        142.3640445651233
+        426.7776456520405
+       -71.70920407779498
+        9.984395040561516
+        195.4775865378649
+        456.0727918302734
+ 5.75e+10    
+        465.3377130940328
+        196.0645082586374
+        427.6432584520452
+        9.046317956628044
+        142.7241505750799
+        427.9263957394932
+       -72.23473767050795
+        9.716779144219974
+        196.1186579019395
+        457.4409084759414
+ 5.76e+10    
+        466.7161424939787
+        196.7035688765147
+        428.7930585262578
+        8.774781960941537
+        143.0843761081394
+        429.0771776896335
+       -72.76117419918339
+        9.447474251598145
+        196.7598327859117
+        458.8119344314014
+ 5.77e+10    
+        468.0974650233316
+          197.34271116506
+        429.9448914708136
+        8.501552229127638
+        143.4447226219942
+        430.2299937355195
+       -73.28850343316901
+        9.176480122271705
+        197.4011024284692
+        460.1858708819686
+ 5.78e+10    
+        469.4816819224852
+        197.9819264794949
+        431.0987597528568
+        8.226628548090041
+        143.8051916666808
+        431.3848462219584
+       -73.81671529385937
+        8.903796525157723
+        198.0424582009801
+        461.5627190532044
+ 5.79e+10    
+        470.8687944834447
+        198.6212063119787
+        432.2546659529034
+        7.950010714229997
+        144.1657848851766
+        432.5417376064736
+       -74.34579985860415
+        8.629423238152189
+        198.6838916105597
+        462.9424802118651
+ 5.8e+10     
+        472.2588040509399
+        199.2605422947036
+        433.4126127657704
+        7.671698533094077
+        144.5265040139941
+        433.7006704602811
+       -74.87574736459877
+        8.353360047772057
+        199.3253943031506
+        464.3251556668497
+ 5.81e+10    
+        473.6517120235467
+        199.8999262030039
+        434.5726030015006
+        7.391691819027216
+        144.8873508837703
+        434.8616474692609
+        -75.4065482127542
+        8.075606748803899
+        199.9669580666173
+        465.7107467701561
+ 5.82e+10    
+        475.0475198548122
+        200.5393499584853
+         435.734639586302
+        7.109990394831728
+        145.2483274198571
+        436.0246714349342
+       -75.93819297154646
+        7.796163143957489
+        200.6085748338564
+        467.0992549178483
+ 5.83e+10    
+        476.4462290543824
+        201.1788056321581
+        436.8987255634722
+        6.826594091430417
+         145.609435642905
+        437.1897452754376
+       -76.47067238084433
+        7.515029043524894
+        201.2502366859171
+         468.490681551017
+ 5.84e+10    
+        477.8478411891456
+        201.8182854475934
+        438.0648640943398
+        6.541502747537608
+        145.9706776694468
+        438.3568720264983
+       -77.00397735571438
+        7.232204265045407
+        201.8919358551369
+         469.885028156752
+ 5.85e+10    
+        479.2523578843667
+        202.4577817840884
+        439.2330584592028
+        6.254716209334346
+        146.3320557124791
+        439.5260548424123
+       -77.53809899020187
+         6.94768863297724
+        202.5336647282919
+         471.282296269126
+ 5.86e+10    
+        480.6597808248355
+        203.0972871798438
+        440.4033120582585
+        5.966234330150364
+        146.6935720820382
+        440.6972969970233
+       -78.07302856108733
+        6.661481978374148
+        203.1754158497579
+        472.6824874701673
+ 5.87e+10    
+        482.0701117560188
+        203.7367943351592
+         441.575628412552
+        5.676056970152068
+        147.0552291857772
+           441.8706018847
+       -78.60875753161699
+        6.373584138569186
+         203.817181924687
+        474.0856033908518
+ 5.88e+10    
+        483.4833524852168
+        204.3762961156388
+        442.7500111649179
+        5.384183996036819
+         147.417029529538
+        443.0459730213182
+       -79.14527755520726
+        6.083994956864707
+        204.4589558221963
+        475.4916457120939
+ 5.89e+10    
+        484.8995048827248
+          205.01578555541
+        443.9264640809209
+        5.090615280733978
+        147.7789757179221
+        444.2234140452426
+       -79.68258047912012
+        5.792714282228303
+        205.1007305785702
+        476.9006161657459
+ 5.9e+10     
+        486.3185708829981
+        205.6552558603569
+        445.1049910498049
+        4.795350703111881
+        148.1410704548576
+        445.4029287183059
+       -80.22065834811168
+        5.499741968996236
+        205.7424994004748
+        478.3125165355975
+ 5.91e+10    
+        487.7405524858284
+        206.2947004113651
+        446.2855960854382
+        4.498390147692303
+        148.5033165441664
+        446.5845209267998
+       -80.75950340804937
+        5.205077876583339
+        206.3842556681854
+        479.7273486583824
+ 5.92e+10    
+         489.165451757511
+        206.9341127675818
+        447.4682833272727
+        4.199733504371164
+        148.8657168901262
+        447.7681946824529
+        -81.2991081094998
+        4.908721869199361
+         207.025992938828
+        481.1451144247948
+ 5.93e+10    
+        490.5932708320423
+        207.5734866696843
+        448.6530570412808
+        3.899380668146721
+        149.2282744980308
+        448.9539541234223
+       -81.83946511128426
+        4.610673815573563
+        207.6677049496313
+        482.5658157805022
+ 5.94e+10    
+        492.0240119122914
+        208.2128160431672
+        449.8399216209273
+        3.597331538854387
+        149.5909924747498
+        450.1418035152775
+       -82.38056728400214
+        4.310933588685018
+         208.309385621193
+        483.9894547271698
+ 5.95e+10    
+         493.457677271202
+        208.8520950016366
+        451.0288815881126
+        3.293586020909501
+         149.953874029284
+        451.3317472519939
+       -82.92240771352085
+        4.009501065501489
+        208.9510290607573
+          485.41603332349
+ 5.96e+10    
+        494.8942692529877
+        209.4913178501193
+        452.2199415941386
+        2.988144023056588
+        150.3169224733188
+        452.5237898569416
+       -83.46497970443083
+        3.706376126725637
+        209.5926295655055
+        486.8455536862094
+ 5.97e+10    
+        496.3337902743283
+         210.130479088385
+        453.4131064206688
+        2.681005458126918
+        150.6801412217767
+        453.7179359838775
+       -84.00827678346646
+         3.40155865654754
+        210.2341816258574
+        488.2780179911702
+ 5.98e+10    
+        497.7762428255897
+        210.7695734142791
+          454.60838098069
+        2.372170242803689
+        151.0435337933657
+        454.9141904179386
+       -84.55229270288861
+        3.095048542406737
+        210.8756799287866
+        489.7134284743511
+ 5.99e+10    
+        499.2216294720191
+        211.4085957270667
+        455.8057703194751
+        2.061638297394131
+        151.4071038111266
+        456.1125580766405
+       -85.09702144383223
+        2.786845674761249
+        211.5171193611476
+        491.1517874329182
+ 6e+10       
+        500.6699528549779
+        212.0475411307926
+        457.0052796155591
+        1.749409545610197
+        151.7708550029775
+        457.3130440108662
+       -85.64245721961427
+        2.476949946864078
+        212.1584950130099
+        492.5930972262668
+ 6.01e+10    
+        502.1212156931549
+        212.6864049376476
+        458.2069141816982
+        1.435483914357938
+        152.1347912022568
+        458.5156534058758
+        -86.1885944790034
+        2.165361254548632
+        212.7998021810126
+        494.0373602770892
+ 6.02e+10    
+        503.5754207837958
+        213.3251826713525
+        459.4106794658534
+        1.119861333533443
+        152.4989163482638
+        459.7203915822966
+       -86.73542790944867
+        1.852079496022615
+        213.4410363717221
+        495.4845790724335
+ 6.03e+10    
+        505.0325710039324
+        213.9638700705451
+        460.6165810521505
+       0.8025417358280595
+        152.8632344867959
+        460.9272639971297
+        -87.2829524402695
+        1.537104571668536
+         214.082193305005
+        496.9347561647648
+ 6.04e+10    
+        506.4926693116246
+        214.6024630921897
+        461.8246246618721
+       0.4835250565419038
+        153.2277497706856
+        462.1362762447519
+       -87.83116324580101
+         1.22043638385513
+        214.7232689174139
+        498.3878941730439
+ 6.05e+10    
+        507.9557187471973
+        215.2409579149877
+        463.0348161544241
+       0.1628112334059892
+        153.5924664603344
+        463.3474340579192
+       -88.38005574849942
+       0.9020748367550127
+        215.3642593655775
+        499.8439957837982
+ 6.06e+10    
+        509.4217224344883
+        215.8793509428056
+        464.2471615283241
+      -0.1595997935874873
+        153.9573889242444
+        464.5607433087744
+       -88.92962562200215
+        0.582019836172929
+         216.005161029612
+        501.3030637522056
+ 6.07e+10    
+        510.8906835820976
+        216.5176388081097
+        465.4616669221783
+      -0.4837080823460198
+        154.3225216395473
+        465.7762100098533
+       -89.47986879414441
+        0.260271289381393
+        216.6459705165324
+        502.7651009031761
+ 6.08e+10    
+         512.362605484646
+        217.1558183754158
+        466.6783386156743
+       -0.809513688828428
+        154.6878691925343
+        466.9938403150977
+       -90.03078144993067
+     -0.06317089503396645
+         217.286684663682
+        504.2301101324466
+ 6.09e+10    
+         513.837491524035
+        217.7938867447472
+        467.8971830305642
+        -1.13701666718792
+        155.0534362791795
+        468.2136405208605
+       -90.58236003445936
+      -0.3883068073199389
+        217.9273005421704
+        505.6980944076761
+ 6.1e+10     
+        515.3153451707051
+        218.4318412550999
+          469.11820673165
+       -1.466217069905891
+        155.4192277056638
+        469.4356170669237
+       -91.13460125580136
+      -0.7151365366931959
+        218.5678154603196
+        507.1690567695367
+ 6.11e+10    
+        516.7961699849168
+        219.0696794879276
+        470.3414164277878
+       -1.797114947916398
+        155.7852483888985
+        470.6597765375143
+       -91.68750208783067
+       -1.043660171467128
+        219.2082269671226
+        508.6430003328272
+ 6.12e+10    
+        518.2799696180173
+        219.7073992706252
+         471.566818972871
+       -2.129710350722437
+        156.1515033570417
+          471.88612566231
+       -92.24105977300654
+       -1.373877799170161
+        219.8485328557117
+         510.119928287574
+ 6.13e+10    
+        519.7667478137155
+        220.3449986800307
+        472.7944213668315
+       -2.464003326501111
+        156.5179977500184
+        473.1146713174671
+       -92.79527182510547
+       -1.705789506654339
+         220.488731166837
+        511.5998439001521
+ 6.14e+10    
+        521.2565084093758
+        220.9824760459335
+        474.0242307566349
+       -2.799993922200745
+        156.8847368200346
+        474.3454205266377
+       -93.35013603190488
+       -2.039395380194941
+        221.1288201923519
+        513.0827505143918
+ 6.15e+10    
+        522.7492553372961
+        221.6198299545935
+        475.2562544372881
+       -3.137682183627525
+        157.2517259320918
+        475.5783804619854
+       -93.90565045781403
+       -2.374695505579357
+        221.7687984787121
+        514.5686515527099
+ 6.16e+10    
+        524.2449926260014
+        222.2570592522679
+        476.4904998528331
+       -3.477068155523432
+        157.6189705644975
+        476.8135584452113
+       -94.46181344645457
+       -2.711689968187326
+        222.4086648304813
+        516.0575505172276
+ 6.17e+10    
+        525.7437244015466
+        222.8941630487512
+        477.7269745973588
+       -3.818151881633137
+        157.9864763093759
+        478.0509619485798
+       -95.01862362318772
+       -3.050378853060671
+        223.0484183138467
+        517.5494509909051
+ 6.18e+10    
+        527.2454548888059
+         223.531140720918
+        478.9656864160041
+       -4.160933404762172
+        158.3542488731754
+         479.290598595938
+       -95.57607989758876
+       -3.390762244963112
+        223.6880582601445
+         519.044356638678
+ 6.19e+10    
+        528.7501884127835
+        224.1679919162816
+        480.2066432059692
+         -4.5054127668249
+        158.7222940771741
+        480.5324761637494
+       -96.13418146586818
+       -3.732840228430621
+        224.3275842693919
+        520.5422712085859
+ 6.2e+10     
+        530.2579293999211
+        224.8047165565579
+        481.4498530175247
+       -4.851590008881837
+        159.0906178579832
+         481.776602582115
+       -96.69292781323679
+       -4.076612887811216
+        224.9669962138313
+        522.0431985329278
+ 6.21e+10    
+        531.7686823794148
+        225.4413148412382
+        482.6953240550267
+       -5.199465171167327
+        159.4592262680505
+        483.0229859358107
+       -97.25231871621682
+       -4.422080307294523
+        225.6062942414787
+        523.5471425293962
+ 6.22e+10    
+         533.282451984522
+        226.0777872511697
+        483.9430646779286
+       -5.549038293107291
+        159.8281254761592
+        484.2716344653138
+        -97.8123542448963
+       -4.769242570931258
+        226.2454787796851
+        525.0541072022376
+ 6.23e+10    
+        534.7992429538883
+        226.7141345521459
+        485.1930834018007
+       -5.900309413326095
+        160.1973217679264
+        485.5225565678359
+       -98.37303476512666
+       -5.118099762642384
+        226.8845505387018
+        526.5640966433984
+ 6.24e+10    
+        536.3190601328749
+        227.3503577985063
+        486.4453888993494
+       -6.253278569643575
+        160.5668215462993
+        486.7757607983594
+       -98.93436094066405
+       -5.468651966217676
+        227.5235105152568
+         528.077115033688
+ 6.25e+10    
+        537.8419084748779
+        227.9864583367386
+        487.6999900014355
+        -6.60794579906131
+        160.9366313320499
+        488.0312558706718
+        -99.4963337352508
+       -5.820899265303852
+        228.1623599961366
+        529.5931666439403
+ 6.26e+10    
+        539.3677930426688
+        228.6224378090949
+        488.9568956980968
+       -6.964311137737804
+        161.3067577642682
+        489.2890506584039
+       -100.0589544146395
+       -6.174841743382174
+        228.8011005617776
+        531.1122558361767
+ 6.27e+10    
+        540.8967190097264
+        229.2582981572119
+        490.2161151395744
+       -7.322374620955314
+        161.6772076008515
+        490.5491541960643
+       -100.6222245485581
+       -6.530479483735363
+        229.4397340898642
+        532.6343870647787
+ 6.28e+10    
+        542.4286916615738
+        229.8940416257386
+        491.4776576373384
+       -7.682136283072841
+        162.0479877189937
+        491.8115756800817
+       -101.1861460126133
+       -6.887812569403785
+        230.0782627589319
+        534.1595648776555
+ 6.29e+10    
+        543.9637163971281
+        230.5296707659724
+         492.741532665114
+       -8.043596157470477
+        162.4191051156747
+        493.0763244698516
+       -101.7507209901357
+       -7.246841083130477
+        230.7166890519829
+        535.6877939174273
+ 6.3e+10     
+        545.5017987300388
+        231.1651884395014
+        494.0077498599097
+       -8.406754276483058
+        162.7905669081414
+        494.3434100887641
+       -102.3159519739621
+       -7.607565107296287
+         231.355015760101
+        537.2190789225976
+ 6.31e+10    
+        547.0429442900443
+        231.8005978218527
+         495.276319023054
+       -8.771610671321469
+        163.1623803343953
+        495.6128422252636
+       -102.8818417681573
+       -7.969984723843252
+        231.9932459860797
+        538.7534247287396
+ 6.32e+10    
+         548.587158824319
+        232.4359024061496
+        496.5472501212215
+       -9.138165371984918
+        163.5345527536711
+        496.8846307338787
+       -103.4483934896728
+       -8.334100014186816
+        232.6313831480543
+        540.2908362696842
+ 6.33e+10    
+        550.1344481988348
+        233.0711060067711
+        497.8205532874709
+       -9.506418407160213
+        163.9070916469188
+        498.1587856362792
+       -104.0156105699432
+       -8.699911059118161
+        233.2694309831376
+        541.8313185787043
+ 6.34e+10    
+        551.6848183997145
+        233.7062127630221
+        499.0962388222788
+       -9.876369804112141
+        164.2800046172799
+        499.4353171223178
+       -104.5834967564196
+        -9.06741793869376
+        233.9073935510676
+        543.3748767897147
+ 6.35e+10    
+        553.2382755346048
+        234.3412271428073
+        500.3743171945792
+       -10.24801958856092
+         164.653299390565
+        500.7142355510767
+        -105.152056114039
+       -9.436620732115964
+        234.5452752378537
+        544.9215161384582
+ 6.36e+10    
+        554.7948258340261
+         234.976153946309
+        501.6547990427985
+       -10.62136778454976
+        165.0269838157271
+        501.9955514519179
+       -105.7212930266287
+       -9.807519517600188
+        235.1830807594347
+         546.471241963711
+ 6.37e+10    
+        556.3544756527587
+        235.6109983096736
+        502.9376951758969
+        -10.9964144143007
+        165.4010658653355
+        503.2792755255337
+       -106.2912121982476
+       -10.18011437223226
+        235.8208151653386
+        548.0240597084818
+ 6.38e+10    
+        557.9172314711985
+        236.2457657087017
+        504.2230165744103
+       -11.37315949805919
+        165.7755536360457
+        504.5654186449984
+       -106.8618186544608
+       -10.55440537181382
+        236.4584838423501
+        549.5799749212166
+ 6.39e+10    
+          559.48309989674
+        236.8804619625438
+        505.5107743914935
+       -11.75160305392771
+        166.1504553490691
+         505.853991856815
+       -107.4331177435495
+        -10.9303925906974
+        237.0960925181787
+        551.1389932570028
+ 6.4e+10     
+        561.0520876651498
+        237.5150932373995
+        506.8009799539597
+       -12.13174509768804
+        166.5257793506408
+        507.1450063819742
+       -108.0051151376541
+       -11.30807610160813
+        237.7336472651374
+        552.7011204787827
+ 6.41e+10    
+        562.6242016419477
+        238.1496660502241
+         508.093644763328
+       -12.51358564261198
+        166.9015341124829
+        508.4384736169999
+       -108.5778168338516
+       -11.68745597545659
+        238.3711545038208
+        554.2663624585598
+ 6.42e+10    
+        564.1994488237864
+        238.7841872724367
+        509.3887804968715
+       -12.89712469926064
+        167.2777282322727
+        509.7344051350132
+       -109.1512291551663
+       -12.06853228113833
+        239.0086210067915
+        555.8347251786184
+ 6.43e+10    
+        565.7778363398364
+        239.4186641336332
+        510.6863990086594
+       -13.28236227527295
+        167.6543704340998
+        511.0328126867763
+       -109.7253587515119
+       -12.45130508532239
+        239.6460539022663
+        557.4062147327375
+ 6.44e+10    
+         567.359371453174
+        240.0531042253053
+        511.9865123306056
+         -13.669298375142
+        168.0314695689304
+        512.3337082017532
+       -110.3002126005677
+       -12.83577445222897
+        240.2834606778109
+        558.9808373274088
+ 6.45e+10    
+        568.9440615621634
+        240.6875155045596
+        513.2891326735225
+       -14.05793299998004
+        168.4090346150637
+        513.6371037891688
+        -110.875798008586
+       -13.22194044339481
+        240.9208491840338
+        560.5585992830574
+ 6.46e+10    
+        570.5319142018575
+        241.3219062978439
+        514.5942724281631
+       -14.44826614727301
+        168.7870746785897
+        514.9430117390564
+       -111.4521226111319
+       -13.60980311742739
+        241.5582276382875
+         562.139507035269
+ 6.47e+10    
+        572.1229370453829
+        241.9562853046729
+        515.9019441662742
+       -14.84029781062187
+        169.1655989938444
+        516.2514445233253
+       -112.0291943737535
+       -13.99936252974781
+        242.1956046283699
+        563.7235671360085
+ 6.48e+10    
+        573.7171379053367
+        242.5906616013624
+        517.2121606416546
+       -15.23402797947367
+        169.5446169238628
+        517.5624147968072
+       -112.6070215925843
+       -14.39061873232094
+        242.8329891162305
+        565.3107862548499
+ 6.49e+10    
+        575.3145247351815
+        243.2250446447587
+        518.5249347911932
+       -15.62945663884123
+        169.9241379608306
+        518.8759353983219
+        -113.185612894877
+        -14.7835717733761
+        243.4703904416764
+        566.9011711802049
+ 6.5e+10     
+         576.915105630645
+        243.8594442759774
+        519.8402797359305
+       -16.02658376900956
+        170.3041717265343
+        520.1920193517324
+       -113.7649772394659
+       -15.17822169711382
+        244.1078183260856
+        568.4947288205501
+ 6.51e+10    
+        578.5188888311208
+        244.4938707241411
+        521.1582087821123
+       -16.42540934523332
+        170.6847279728101
+        521.5106798670025
+       -114.3451239171625
+       -15.57456854340247
+        244.7452828761187
+        570.0914662056631
+ 6.52e+10    
+        580.1258827210668
+        245.1283346101203
+        522.4787354222379
+        -16.8259333374207
+        171.0658165819889
+        522.8319303412566
+       -114.9260625510792
+       -15.97261234746306
+        245.3827945874325
+        571.6913904878496
+ 6.53e+10    
+        581.7360958314077
+         245.762846950274
+        523.8018733361137
+       -17.22815570980639
+        171.4474475673421
+         524.155784359837
+       -115.5078030968842
+       -16.37235313954186
+        246.0203643483975
+        573.2945089431814
+ 6.54e+10    
+        583.3495368409424
+        246.3974191601961
+        525.1276363919158
+       -17.63207642061308
+        171.8296310735252
+        525.4822556973648
+       -116.0903558429857
+       -16.77379094457199
+        246.6580034438161
+        574.9008289727333
+ 6.55e+10    
+        584.9662145777422
+        247.0320630584577
+        526.4560386472339
+       -18.03769542170194
+        172.2123773770174
+         526.811358318792
+       -116.6737314106466
+       -17.17692578182272
+        247.2957235586398
+        576.5103581038122
+ 6.56e+10    
+        586.5861380205629
+        247.6667908703547
+        527.7870943501323
+       -18.44501265820968
+         172.595696886563
+        528.1431063804728
+        -117.257940754028
+       -17.58175766453859
+        247.9335367816914
+        578.1231039912029
+ 6.57e+10    
+        588.2093163002518
+        248.3016152316564
+        529.1208179402037
+       -18.85402806817685
+        172.9796001436086
+        529.4775142312093
+       -117.8429951601633
+       -17.98828659956516
+        248.5714556093848
+        579.7390744184002
+ 6.58e+10    
+        589.8357587011485
+        248.9365491923487
+        530.4572240496199
+       -19.26474158216189
+        173.3640978227388
+        530.8145964133142
+       -118.4289062488591
+       -18.39651258696395
+        249.2094929494459
+        581.3582772988506
+ 6.59e+10    
+        591.4654746624996
+        249.5716062203866
+        531.7963275041939
+       -19.67715312284589
+        173.7492007321113
+        532.1543676636717
+       -119.0156859725299
+       -18.80643561961611
+        249.8476621246343
+        582.9807206771923
+ 6.6e+10     
+        593.0984737798678
+        250.2068002054394
+        533.1381433244292
+       -20.09126260462372
+        174.1349198138905
+        533.4968429147955
+       -119.6033466159573
+       -19.21805568281429
+        250.4859768764659
+        584.6064127304943
+ 6.61e+10    
+        594.7347658065371
+        250.8421454626393
+         534.482686726576
+       -20.50706993318602
+        174.5212661446762
+        534.8420372958802
+       -120.1919007959813
+       -19.63137275384249
+        251.1244513689319
+        586.2353617694959
+ 6.62e+10    
+        596.3743606549253
+        251.4776567363273
+        535.8299731236855
+       -20.92457500508789
+        174.9082509359353
+        536.1899661338629
+        -120.781361461121
+       -20.04638680154561
+        251.7631001922212
+        587.8675762398505
+ 6.63e+10    
+         598.017268397996
+        252.1133492038023
+        537.1800181266671
+       -21.34377770730675
+        175.2958855344285
+        537.5406449544799
+       -121.3717418911213
+       -20.46309778588553
+        252.4019383664392
+        589.5030647233637
+ 6.64e+10    
+        599.6634992706641
+        252.7492384790648
+        538.5328375453371
+       -21.76467791678904
+         175.684181422636
+         538.894089483323
+       -121.9630556964338
+       -20.88150565748849
+        253.0409813453261
+        591.1418359392312
+ 6.65e+10    
+        601.3130636712127
+        253.3853406165599
+         539.888447389473
+       -22.18727549998528
+        176.0731502191819
+        540.2503156468894
+        -122.555316817622
+       -21.30161035717769
+        253.6802450199765
+        592.7838987452905
+ 6.66e+10    
+        602.9659721626913
+        254.0216721149232
+        541.2468638698726
+       -22.61157031237385
+        176.4628036792571
+        541.6093395736463
+       -123.1485395246987
+       -21.72341181549785
+        254.3197457225522
+        594.4292621392497
+ 6.67e+10    
+        604.6222354743425
+        254.6582499207195
+        542.6081033993991
+       -23.03756219797388
+          176.85315369504
+        542.9711775950738
+       -123.7427384163934
+       -22.14690995222606
+        254.9595002299985
+        596.0779352599349
+ 6.68e+10    
+        606.2818645029989
+        255.2950914321832
+        543.9721825940378
+       -23.46525098884536
+        177.2442122961153
+         544.335846246727
+       -124.3379284193449
+       -22.57210467587188
+        255.5995257677541
+        597.7299273885285
+ 6.69e+10    
+        607.9448703144939
+        255.9322145029514
+        545.3391182739408
+       -23.89463650458067
+        177.6359916498915
+        545.7033622692819
+       -124.9341247872295
+       -22.99899588316712
+        256.2398400134624
+        599.3852479498048
+ 6.7e+10     
+        609.6112641450774
+        256.5696374458042
+        546.7089274644874
+       -24.32571855178224
+        178.0285040620166
+        547.0737426095898
+       -125.5313430998139
+        -23.4275834585428
+        256.8804611006764
+        601.0439065133739
+ 6.71e+10    
+        611.2810574028132
+        257.2073790363882
+        548.0816273973215
+         -24.758496923531
+        178.4217619767924
+        548.4470044217262
+       -126.1295992619402
+       -23.85786727359649
+        257.5214076225639
+         602.705912794919
+ 6.72e+10    
+        612.9542616689965
+         257.845458516952
+        549.4572355114121
+       -25.19297139884241
+        178.8157779775867
+        549.8231650680405
+       -126.7289095024408
+       -24.28984718654707
+        258.1626986356077
+        604.3712766574308
+ 6.73e+10    
+        614.6308886995494
+        258.4838956000639
+        550.8357694540886
+       -25.62914174211272
+        179.2105647872429
+        551.2022421202018
+       -127.3292903729833
+       -24.72352304168005
+        258.8043536633014
+        606.0400081124423
+ 6.74e+10    
+        616.3109504264348
+        259.1227104723378
+        552.2172470820975
+       -26.06700770255327
+        179.6061352684906
+        552.5842533602483
+       -127.9307587468451
+          -25.15889466878
+        259.4463926998449
+        607.7121173212657
+ 6.75e+10    
+        617.9944589590558
+        259.7619237981488
+        553.6016864626442
+        -26.5065690136137
+        180.0025024243517
+        553.9692167816313
+       -128.5333318176194
+       -25.59596188255323
+        260.0888362138322
+        609.3876145962286
+ 6.76e+10    
+        619.6814265856563
+        260.4015567233434
+        554.9891058744303
+       -26.94782539239633
+        180.3996793985453
+        555.3571505902549
+       -129.1370270978531
+       -26.03472448203996
+        260.7317051519362
+        611.0665104018966
+ 6.77e+10    
+        621.3718657747246
+         261.041630878951
+         556.379523808706
+       -27.39077653905712
+        180.7976794758932
+        556.7480732055271
+       -129.7418624176126
+       -26.47518225001398
+        261.3750209425917
+        612.7488153563158
+ 6.78e+10    
+        623.0657891763954
+        261.6821683848859
+        557.7729589703058
+       -27.83542213619696
+        181.1965160827203
+        558.1420032613923
+       -130.3478559229841
+       -26.91733495237312
+        262.0188054996667
+        614.4345402322286
+ 6.79e+10    
+        624.7632096238382
+        262.3231918536453
+        559.1694302786914
+       -28.28176184824351
+        181.5962027872552
+        559.5389596073705
+       -130.9550260745048
+       -27.36118233751835
+        262.6630812261363
+        616.1236959583111
+ 6.8e+10     
+        626.4641401346628
+        262.9647243940023
+        560.5689568689829
+       -28.72979532082026
+        181.9967533000306
+        560.9389613096039
+        -131.563391645525
+        -27.8067241357224
+        263.3078710177466
+         617.816293620391
+ 6.81e+10    
+        628.1685939123045
+        263.6067896146927
+        561.9715580930038
+        -29.1795221801073
+        182.3981814742764
+        562.3420276518754
+       -132.1729717205035
+       -28.25396005848769
+        263.9531982666721
+        619.5123444626713
+ 6.82e+10    
+        629.8765843474258
+         264.249411628098
+        563.3772535203092
+       -29.63094203218945
+          182.80050130632
+         563.748178136664
+       -132.7837856932353
+       -28.70288979789371
+         264.599086865173
+        621.2118598889533
+ 6.83e+10    
+        631.5881250192929
+        264.8926150539188
+        564.7860629392227
+        -30.0840544623963
+        183.2037269359751
+        565.1574324861562
+       -133.3958532650128
+       -29.15351302593443
+        265.2455612092378
+        622.9148514638505
+ 6.84e+10    
+        633.3032296971726
+        265.5364250228441
+        566.1980063578656
+       -30.53885903463039
+        183.6078726469365
+        566.5698106432867
+       -134.0091944427206
+       -29.60582939384507
+        265.8926462022275
+        624.6213309140101
+ 6.85e+10    
+        635.0219123417113
+        266.1808671802133
+        567.6131040051857
+       -30.99535529068568
+        184.0129528671686
+        567.9853327727624
+       -134.6238295368618
+       -30.05983853141853
+        266.5403672585049
+        626.3313101293143
+ 6.86e+10    
+         636.744187106319
+        266.8259676896691
+        569.0313763319824
+        -31.4535427495563
+        184.4189821692952
+        569.4040192620907
+       -135.2397791595222
+       -30.51554004631197
+        267.1887503070664
+        628.0448011641065
+ 6.87e+10    
+        638.4700683385479
+        267.4717532368084
+        570.4528440119356
+        -31.9134209067351
+        184.8259752709843
+         570.825890722597
+       -135.8570642222674
+       -30.97293352334353
+        267.8378217951552
+        629.7618162383803
+ 6.88e+10    
+        640.1995705814655
+        268.1182510328189
+        571.8775279426281
+       -32.37498923350153
+        185.2339470353349
+        572.2509679904516
+        -136.475705933973
+       -31.43201852377802
+        268.4876086918786
+         631.482367739002
+ 6.89e+10    
+        641.9327085750319
+        268.7654888181112
+        573.3054492465581
+       -32.83824717620133
+        185.6429124712589
+        573.6792721276809
+       -137.0957257985944
+       -31.89279458460429
+        269.1381384918044
+        633.2064682208916
+ 6.9e+10     
+        643.6694972574664
+        269.4134948659449
+        574.7366292721675
+       -33.30319415551489
+        186.0528867338636
+        575.1108244231903
+       -137.7171456128694
+       -32.35526121780151
+        269.7894392185634
+        634.9341304082387
+ 6.91e+10    
+        645.4099517666116
+        270.0622979860391
+        576.1710895948488
+       -33.76982956571726
+        186.4638851248307
+         576.545646393771
+       -138.3399874639594
+       -32.81941790959692
+        270.4415394284296
+        636.6653671956838
+ 6.92e+10    
+        647.1540874413034
+         270.711927528183
+        577.6088520179632
+       -34.23815277392762
+        186.8759230927956
+        577.9837597851168
+       -138.9642737270265
+       -33.28526411971276
+        271.0944682139011
+        638.4001916495148
+ 6.93e+10    
+        648.9019198227227
+        271.3624133858309
+        579.0499385738498
+       -34.70816311935054
+        187.2890162337224
+        579.4251865728266
+       -139.5900270627492
+        -33.7527992806052
+         271.748255207268
+         640.138617008851
+ 6.94e+10    
+         650.653464655757
+        272.0137859996888
+         580.494371524829
+       -35.17985991250641
+         187.703180291279
+        580.8699489634074
+       -140.2172704147748
+       -34.22202279669228
+        272.4029305841697
+        641.8806566868279
+ 6.95e+10    
+        652.4087378903448
+        272.6660763612945
+        581.9421733642112
+       -35.65324243445426
+        188.1184311572115
+        582.3180693952867
+       -140.8460270071122
+       -34.69293404357467
+        273.0585250671467
+        643.6263242717719
+ 6.96e+10    
+        654.1677556828304
+         273.319316016585
+        583.3933668172982
+       -36.12830993600421
+        188.5347848717134
+        583.7695705397981
+       -141.4763203414633
+       -35.16553236724459
+        273.7150699291774
+        645.3756335283821
+ 6.97e+10    
+        655.9305343973056
+        273.9735370694526
+        584.8479748423807
+       -36.60506163692239
+        188.9522576237972
+        585.2244753021864
+       -142.1081741944944
+       -35.63981708328862
+        274.3725969972085
+        647.1285983988926
+ 6.98e+10    
+        657.6970906069436
+        274.6287721852935
+        586.3060206317319
+       -37.08349672512547
+        189.3708657516595
+        586.6828068225946
+       -142.7416126150479
+       -36.11578747607965
+        275.0311386556716
+        648.8852330042441
+ 6.99e+10    
+        659.4674410953395
+        275.2850545945431
+         587.767527612604
+       -37.56361435586733
+        189.7906257430509
+        588.1445884770611
+       -143.3766599212957
+       -36.59344279796058
+        275.6907278499929
+        650.6455516452429
+ 7e+10       
+        661.2416028578411
+         275.942418096203
+        589.2325194482166
+       -38.04541365091759
+        190.2115542356375
+        589.6098438784957
+       -144.0133406978339
+       -37.07278226841991
+        276.3513980900868
+        652.4095688037188
* NOTE: Solution at 1e+08 Hz used as DC point.

.model l_m4lines_HFSS_W_1 sp N=4 SPACING=nonuniform VALTYPE=real
+ INTERPOLATION=spline
+ INFINITY =
+    4.771275496612187e-07
+    1.992620892018445e-07
+    4.599493106995181e-07
+    6.333700301101069e-08
+    1.283548577953231e-07
+    4.599264508819013e-07
+    2.830257265266555e-08
+    6.339692795622215e-08
+    1.993667267423742e-07
+    4.775330895971331e-07
+ DATA = 700
+ 0           
+    4.187375639716964e-07
+    1.499780296080442e-07
+    4.160104447847029e-07
+    4.559175281127766e-08
+      9.3362516970571e-08
+    4.159107655224221e-07
+    2.474797370846747e-08
+    4.559883258452768e-08
+    1.500178654245671e-07
+     4.18915896522694e-07
+ 2e+08       
+    4.152409295458201e-07
+    1.496357305871249e-07
+    4.124619577225161e-07
+    4.548151148332848e-08
+      9.2913481972087e-08
+    4.123676835644636e-07
+    2.471316967566081e-08
+    4.548809260884237e-08
+    1.496823467245008e-07
+    4.154633204210293e-07
+ 3e+08       
+    4.136486656757639e-07
+    1.495163480809376e-07
+    4.108544222836318e-07
+    4.542229773637365e-08
+    9.271611584391797e-08
+    4.107642254925401e-07
+    2.469173623432938e-08
+    4.542794895367581e-08
+    1.495623570531414e-07
+    4.138979002356905e-07
+ 4e+08       
+    4.127491121110181e-07
+    1.494674564879319e-07
+    4.099434383939512e-07
+    4.539229528127803e-08
+    9.260776279126221e-08
+    4.098566144861343e-07
+    2.468312840559359e-08
+    4.539725852963568e-08
+    1.495126419631506e-07
+    4.130184879975287e-07
+ 5e+08       
+    4.121313746128284e-07
+    1.494315581240394e-07
+    4.093168219391762e-07
+    4.537387643230625e-08
+    9.253361250161293e-08
+    4.092328666957902e-07
+    2.467882915622239e-08
+    4.537829677420827e-08
+    1.494763879888115e-07
+    4.124167743840308e-07
+ 6e+08       
+    4.116606371114502e-07
+    1.493998803351824e-07
+    4.088397915546797e-07
+     4.53606269268681e-08
+    9.247712803445569e-08
+    4.087582166247306e-07
+    2.467580053249492e-08
+    4.536458521887698e-08
+    1.494446090073347e-07
+     4.11959011756301e-07
+ 7e+08       
+    4.112849431016661e-07
+    1.493727465672836e-07
+    4.084597465168611e-07
+    4.535032585077475e-08
+    9.243225166966005e-08
+    4.083801157525448e-07
+    2.467331398647141e-08
+    4.535388116828527e-08
+    1.494174616029349e-07
+    4.115940282130534e-07
+ 8e+08       
+    4.109786239826518e-07
+     1.49350648695808e-07
+    4.081501796886804e-07
+    4.534212976387202e-08
+    9.239595057502099e-08
+    4.080721446939833e-07
+    2.467133421986299e-08
+    4.534533432088021e-08
+    1.493953604773808e-07
+    4.112967749299486e-07
+ 9e+08       
+    4.107254835411902e-07
+    1.493331689259142e-07
+    4.078942439898151e-07
+    4.533562699302215e-08
+    9.236622925020992e-08
+    4.078175450740826e-07
+    2.466995580577002e-08
+     4.53385281155439e-08
+    1.493778561619893e-07
+    4.110514931708178e-07
+ 1e+09       
+    4.105136024924595e-07
+    1.493193440705552e-07
+    4.076796662179595e-07
+    4.533053841996527e-08
+    9.234158265688879e-08
+    4.076041127226923e-07
+     2.46692448524731e-08
+    4.533317717036472e-08
+    1.493639705729949e-07
+    4.108465377447294e-07
+ 1.1e+09     
+    4.103023716928628e-07
+     1.49313947387997e-07
+    4.074380291582628e-07
+    4.531980943518837e-08
+    9.231461011155443e-08
+    4.073634695051537e-07
+    2.466308647032362e-08
+    4.532241960162495e-08
+    1.493587597973719e-07
+    4.106421840425814e-07
+ 1.2e+09     
+    4.101179800860868e-07
+    1.493093538467062e-07
+    4.072374741600299e-07
+    4.531139755840584e-08
+    9.229081786787945e-08
+     4.07163855472372e-07
+    2.465802306187109e-08
+    4.531396376427121e-08
+    1.493543421667787e-07
+     4.10464305303107e-07
+ 1.3e+09     
+    4.099576930813259e-07
+    1.493054659480915e-07
+    4.070701907588902e-07
+    4.530517538927157e-08
+    9.227005509960278e-08
+    4.069974460116692e-07
+    2.465405391307196e-08
+    4.530768109316568e-08
+    1.493506134246402e-07
+     4.10310109727224e-07
+ 1.4e+09     
+    4.098185415518215e-07
+    1.493021952857321e-07
+    4.069296716684634e-07
+    4.530099964468045e-08
+    9.225207118843113e-08
+    4.068577274532445e-07
+    2.465116019412628e-08
+    4.530342740541275e-08
+     1.49347480516876e-07
+    4.101765986322123e-07
+ 1.5e+09     
+    4.096976163832522e-07
+     1.49299464978453e-07
+    4.068106135835024e-07
+    4.529872465546234e-08
+    9.223659425171136e-08
+    4.067393950881482e-07
+     2.46493124160821e-08
+    4.530105642140413e-08
+    1.493448639131783e-07
+    4.100608545173434e-07
+ 1.6e+09     
+    4.095922298660851e-07
+    1.492972120491388e-07
+    4.067087528225239e-07
+    4.529820805724975e-08
+    9.222336745289981e-08
+    4.066381869523635e-07
+    2.464847531937749e-08
+    4.530042547353725e-08
+    1.493426996926803e-07
+     4.09960196803909e-07
+ 1.7e+09     
+    4.094999904521203e-07
+    1.492953887664738e-07
+     4.06620691619622e-07
+     4.52993123139985e-08
+    9.221216327266082e-08
+    4.065507088881004e-07
+    2.464861089323851e-08
+    4.530139705186902e-08
+    1.493409405237129e-07
+    4.098722519137703e-07
+ 1.8e+09     
+    4.094188243047893e-07
+    1.492939627485588e-07
+    4.065437386507315e-07
+    4.530190416035827e-08
+    9.220278675277345e-08
+    4.064742742538015e-07
+    2.464968009371305e-08
+    4.530383827659352e-08
+    1.493395554067979e-07
+    4.097949710907745e-07
+ 1.9e+09     
+    4.093469662317995e-07
+    1.492929160288452e-07
+     4.06475771754273e-07
+    4.530585316550455e-08
+    9.219507359464662e-08
+     4.06406766101025e-07
+    2.465164369859237e-08
+    4.530761949868568e-08
+    1.493385284189872e-07
+     4.09726618451859e-07
+ 2e+09       
+    4.092829345740905e-07
+    1.492922434206536e-07
+    4.064151236971854e-07
+    4.531103012501526e-08
+     9.21888861896109e-08
+    4.063465225779688e-07
+    2.465446262747277e-08
+    4.531261273070195e-08
+    1.493378568117296e-07
+    4.096657437132563e-07
+ 2.1e+09     
+    4.092254990762207e-07
+    1.492919505113622e-07
+    4.063604889247688e-07
+    4.531730570836218e-08
+    9.218410914652992e-08
+    4.062922434396572e-07
+     2.46580979683341e-08
+    4.531869032854262e-08
+    1.493375487960881e-07
+     4.09611148486786e-07
+ 2.2e+09     
+    4.091736470856249e-07
+     1.49292051554243e-07
+    4.063108483017992e-07
+    4.532454962793395e-08
+    9.218064507628079e-08
+     4.06242914634344e-07
+    2.466251088553173e-08
+     4.53257241820517e-08
+    1.493376212788093e-07
+    4.095618513738323e-07
+ 2.3e+09     
+    4.091265510695991e-07
+    1.492925674495874e-07
+    4.062654088022628e-07
+    4.533263049362978e-08
+    9.217841096745592e-08
+    4.061977478984043e-07
+    2.466766253329167e-08
+     4.53335855700811e-08
+    1.493380977330648e-07
+    4.095170547413185e-07
+ 2.4e+09     
+    4.090835389694563e-07
+    1.492935239372434e-07
+    4.062235554051074e-07
+    4.534141644202661e-08
+     9.21773352659368e-08
+    4.061561326000178e-07
+    2.467351405901589e-08
+    4.534214576124277e-08
+    1.493390063171503e-07
+     4.09476114611151e-07
+ 2.5e+09     
+    4.090440680228954e-07
+    1.492949500665817e-07
+    4.061848128573086e-07
+    4.535077656270183e-08
+    9.217735565666241e-08
+    4.061175974809551e-07
+    2.468002674818133e-08
+    4.535127737693859e-08
+    1.493403782986581e-07
+    4.094385142223174e-07
+ 2.6e+09     
+    4.090077021681668e-07
+    1.492968769675921e-07
+    4.061488153660386e-07
+    4.536058307775446e-08
+    9.217841748726707e-08
+    4.060817803495908e-07
+    2.468716233474853e-08
+     4.53608564697281e-08
+    1.493422468003602e-07
+    4.094038413219091e-07
+ 2.7e+09     
+    4.089740928580227e-07
+     1.49299336916312e-07
+    4.061152826376026e-07
+    4.537071416190985e-08
+    9.218047274296577e-08
+    4.060484041363018e-07
+    2.469488347639809e-08
+    4.537076520554781e-08
+    1.493446458548759e-07
+    4.093717689685063e-07
+ 2.8e+09     
+     4.08942962967895e-07
+    1.493023626667046e-07
+    4.060840009812158e-07
+    4.538105722294484e-08
+    9.218347946633779e-08
+    4.060172580242864e-07
+    2.470315437231024e-08
+    4.538089497548056e-08
+    1.493476097355371e-07
+    4.093420394985364e-07
+ 2.9e+09     
+    4.089140934242439e-07
+    1.493059870074902e-07
+     4.06054808442822e-07
+    4.539151240234282e-08
+    9.218740150822103e-08
+    4.059881826169183e-07
+    2.471194148323646e-08
+    4.539114970788544e-08
+    1.493511725185679e-07
+    4.093144512565695e-07
+ 3e+09       
+    4.088873121700225e-07
+    1.493102424948618e-07
+    4.060275831350117e-07
+    4.540199601295551e-08
+    9.219220849461252e-08
+    4.059610583043086e-07
+    2.472121430049433e-08
+    4.540144911275184e-08
+    1.493553678252855e-07
+    4.092888476885899e-07
+ 3.1e+09     
+    4.088624851029855e-07
+    1.493151613096188e-07
+    4.060022340917775e-07
+    4.541244361276308e-08
+    9.219787589905706e-08
+      4.0593579615498e-07
+    2.473094610357646e-08
+    4.541173157503836e-08
+    1.493602286915321e-07
+    4.092651084215351e-07
+ 3.2e+09     
+    4.088395086559701e-07
+    1.493207751893492e-07
+    4.059786941089321e-07
+    4.542281242795748e-08
+    9.220438512085534e-08
+    4.059123307911434e-07
+    2.474111464625371e-08
+    4.542195642813171e-08
+    1.493657875142982e-07
+    4.092431419899407e-07
+ 3.3e+09     
+     4.08818303728453e-07
+    1.493271153922281e-07
+    4.059569141387934e-07
+    4.543308288639115e-08
+    9.221172348652262e-08
+    4.058906148144183e-07
+    2.475170271848867e-08
+    4.543210538399082e-08
+    1.493720760318011e-07
+    4.092228799136224e-07
+ 3.4e+09     
+    4.087988107208695e-07
+    1.493342126579206e-07
+    4.059368588962374e-07
+    4.544325910015766e-08
+    9.221988411436768e-08
+    4.058706144379019e-07
+    2.476269854519164e-08
+    4.544218296939753e-08
+    1.493791253023401e-07
+    4.092042718744959e-07
+ 3.5e+09     
+    4.087809854643483e-07
+    1.493420971418513e-07
+    4.059185034060719e-07
+    4.545336823428701e-08
+    9.222886560791143e-08
+    4.058523060539962e-07
+    2.477409600079297e-08
+    4.545221590939256e-08
+    1.493869656579751e-07
+    4.091872817830727e-07
+ 3.6e+09     
+    4.087647958767149e-07
+    1.493507983104362e-07
+     4.05901830281544e-07
+    4.546345880387122e-08
+    9.223867157040068e-08
+     4.05835673527847e-07
+    2.478589463796759e-08
+    4.546225149712845e-08
+    1.493956266202531e-07
+     4.09171884564078e-07
+ 3.7e+09     
+    4.087502192095283e-07
+    1.493603447954113e-07
+    4.058868275725229e-07
+    4.547359803952307e-08
+    9.224930995689621e-08
+    4.058207060555269e-07
+    2.479809954657845e-08
+    4.547235508044201e-08
+     1.49405136775563e-07
+    4.091580635249641e-07
+ 3.8e+09     
+    4.087372397797132e-07
+    1.493707642139923e-07
+    4.058734870608567e-07
+    4.548386853772584e-08
+    9.226079229963914e-08
+    4.058073964653985e-07
+    2.481072107237752e-08
+    4.548260686732339e-08
+    1.494155236161578e-07
+    4.091458082001356e-07
+ 3.9e+09     
+    4.087258471027816e-07
+    1.493820829675042e-07
+     4.05861802910825e-07
+    4.549436445935751e-08
+    9.227313285481481e-08
+    4.057957398717618e-07
+    2.482377443249762e-08
+    4.549309829677787e-08
+    1.494268133587345e-07
+    4.091351125873177e-07
+ 4e+09       
+    4.087160343627817e-07
+    1.493943260340238e-07
+    4.058517706056025e-07
+    4.550518755306532e-08
+    9.228634772377323e-08
+    4.057857326128654e-07
+    2.483727926579862e-08
+    4.550392823511257e-08
+    1.494390307554059e-07
+    4.091259737108543e-07
+ 4.1e+09     
+      4.0870779716755e-07
+    1.494075167706951e-07
+    4.058433861174505e-07
+    4.551644326258927e-08
+    9.230045399975272e-08
+    4.057773714220819e-07
+    2.485125915142909e-08
+    4.551519924237481e-08
+     1.49452198912161e-07
+    4.091183904604241e-07
+ 4.2e+09     
+    4.087011325473754e-07
+    1.494216767392689e-07
+    4.058366452711766e-07
+    4.552823713531653e-08
+    9.231546898364392e-08
+    4.057706527926061e-07
+    2.486574112018972e-08
+    4.552701411560095e-08
+    1.494663391279866e-07
+    4.091123626634329e-07
+ 4.3e+09     
+    4.086960381617356e-07
+    1.494368255648687e-07
+    4.058315432685033e-07
+    4.554067169261696e-08
+    9.233140950131012e-08
+    4.057655725038818e-07
+    2.488075517261178e-08
+    4.553947286315046e-08
+    1.494814707645036e-07
+    4.091078903561924e-07
+ 4.4e+09     
+    4.086925116832874e-07
+    1.494529808338191e-07
+    4.058280743464211e-07
+    4.555384386050909e-08
+    9.234829134252738e-08
+    4.057621252831136e-07
+    2.489633380726949e-08
+    4.555267020661588e-08
+    1.494976111519988e-07
+    4.091049732237159e-07
+ 4.5e+09     
+    4.086905503315881e-07
+    1.494701580323015e-07
+    4.058262315463816e-07
+    4.556784300029692e-08
+    9.236612882953408e-08
+    4.057603045787683e-07
+    2.491251155453083e-08
+    4.556669365139024e-08
+     1.49514775533836e-07
+     4.09103610181438e-07
+ 4.6e+09     
+    4.086901505316665e-07
+    1.494883705241404e-07
+    4.058260065739285e-07
+    4.558274952896952e-08
+    9.238493451280149e-08
+    4.057601024255448e-07
+     2.49293245058738e-08
+    4.558162211963202e-08
+    1.495329770478755e-07
+    4.091037990749024e-07
+ 4.7e+09     
+     4.08691307675033e-07
+    1.495076295634664e-07
+    4.058273897306645e-07
+    4.559863408163281e-08
+    9.240471898370507e-08
+    4.057615093824734e-07
+    2.494680982748013e-08
+    4.559752510327294e-08
+    1.495522267410389e-07
+    4.091055364759525e-07
+ 4.8e+09     
+    4.086940159631406e-07
+    1.495279443364396e-07
+    4.058303699025274e-07
+    4.561555714386565e-08
+    9.242549078853013e-08
+    4.057645145278554e-07
+    2.496500524882297e-08
+    4.561446227082643e-08
+    1.495725336115965e-07
+    4.091088175563502e-07
+ 4.9e+09     
+    4.086982683158349e-07
+    1.495493220255619e-07
+    4.058349345903738e-07
+    4.563356906960552e-08
+    9.244725642549882e-08
+    4.057691054967551e-07
+    2.498394852161705e-08
+     4.56324834492293e-08
+    1.495939046730801e-07
+    4.091136360221986e-07
+ 5e+09       
+    4.087040563298485e-07
+    1.495717678901985e-07
+    4.058410699708904e-07
+    4.565271039781611e-08
+    9.247002040586535e-08
+    4.057752685488218e-07
+    2.500367685073171e-08
+    4.565162889887471e-08
+    1.496163450337679e-07
+    4.091199840949648e-07
+ 5.1e+09     
+    4.087113702749138e-07
+    1.495952853575524e-07
+    4.058487609778119e-07
+    4.567301238608263e-08
+    9.249378536104272e-08
+    4.057829886562276e-07
+    2.502422630529658e-08
+    4.567192980393569e-08
+    1.496398579862442e-07
+    4.091278525272889e-07
+ 5.2e+09     
+    4.087201991173942e-07
+    1.496198761192551e-07
+    4.058579913952957e-07
+    4.569449768881112e-08
+     9.25185521796722e-08
+    4.057922496034325e-07
+    2.504563122418165e-08
+    4.569340890858603e-08
+     1.49664445102409e-07
+     4.09137230644002e-07
+ 5.3e+09     
+    4.087305305634822e-07
+    1.496455402298021e-07
+    4.058687439570582e-07
+    4.571718111958277e-08
+    9.254432016105533e-08
+    4.058030340922708e-07
+    2.506792363445185e-08
+    4.571608124065117e-08
+    1.496901063303053e-07
+    4.091481064008032e-07
+ 5.4e+09     
+     4.08742351115848e-07
+    1.496722762040862e-07
+    4.058810004463853e-07
+    4.574107044966891e-08
+    9.257108717405958e-08
+    4.058153238474461e-07
+    2.509113270375001e-08
+    4.573995487586395e-08
+    1.497168400901184e-07
+    4.091604664547982e-07
+ 5.5e+09     
+    4.087556461391599e-07
+    1.497000811122043e-07
+    4.058947417934993e-07
+    4.576616720650743e-08
+    9.259884981321986e-08
+    4.058290997188821e-07
+    2.511528424765979e-08
+    4.576503170705702e-08
+    1.497446433675838e-07
+    4.091742962425735e-07
+ 5.6e+09     
+    4.087703999311363e-07
+    1.497289506704714e-07
+    4.059099481678613e-07
+    4.579246744634822e-08
+    9.262760354612205e-08
+    4.058443417785236e-07
+     2.51404003110706e-08
+    4.579130819255288e-08
+    1.497735118037636e-07
+    4.091895800626527e-07
+ 5.7e+09     
+     4.08786595796733e-07
+    1.497588793281389e-07
+    4.059265990638981e-07
+    4.581996248392159e-08
+    9.265734284817594e-08
+    4.058610294101015e-07
+    2.516649883879037e-08
+    4.581877606635003e-08
+    1.498034397806982e-07
+    4.092063011600717e-07
+ 5.8e+09     
+    4.088042161237542e-07
+    1.497898603497163e-07
+    4.059446733793668e-07
+    4.584863956883056e-08
+     9.26880613225412e-08
+    4.058791413911031e-07
+    2.519359344567799e-08
+    4.584742299934712e-08
+    1.498344205028275e-07
+    4.092244418114831e-07
+ 5.9e+09     
+    4.088232424586879e-07
+    1.498218858930391e-07
+    4.059641494860891e-07
+    4.587848250352758e-08
+    9.271975180426359e-08
+    4.058986559667225e-07
+    2.522169329101265e-08
+    4.587723320591379e-08
+    1.498664460743107e-07
+     4.09243983409668e-07
+ 6e+09       
+     4.08843655581888e-07
+    1.498549470833588e-07
+     4.05985005293207e-07
+    4.590947220143908e-08
+    9.275240644865199e-08
+    4.059195509159714e-07
+    2.525080305627562e-08
+     4.59081879937904e-08
+    1.498995075724995e-07
+     4.09264906546641e-07
+ 6.1e+09     
+    4.088654355814573e-07
+    1.498890340837741e-07
+    4.060072183033707e-07
+    4.594158718632147e-08
+     9.27860168046155e-08
+    4.059418036103954e-07
+    2.528092302049932e-08
+    4.594026625783644e-08
+    1.499335951178655e-07
+    4.092871910947592e-07
+ 6.2e+09     
+     4.08888561925329e-07
+    1.499241361623148e-07
+    4.060307656624437e-07
+    4.597480403554252e-08
+    9.282057387414623e-08
+      4.0596539106602e-07
+    2.531204922321252e-08
+    4.597344491980281e-08
+    1.499686979406736e-07
+    4.093108162853767e-07
+ 6.3e+09     
+    4.089130135311413e-07
+    1.499602417559577e-07
+    4.060556242034325e-07
+    4.600909777091332e-08
+     9.28560681594108e-08
+    4.059902899892424e-07
+    2.534417370199207e-08
+    4.600769931729583e-08
+    1.500048044446616e-07
+    4.093357607846805e-07
+ 6.4e+09     
+    4.089387688335738e-07
+    1.499973385317989e-07
+    4.060817704853572e-07
+    4.604444220115463e-08
+     9.28924896990565e-08
+    4.060164768174306e-07
+    2.537728478979841e-08
+    4.604300354562842e-08
+    1.500419022679331e-07
+    4.093620027664066e-07
+ 6.5e+09     
+     4.08965805848884e-07
+    1.500354134455695e-07
+    4.061091808278247e-07
+    4.608081022023591e-08
+     9.29298280953765e-08
+    4.060439277549805e-07
+    2.541136745656806e-08
+    4.607933075646776e-08
+    1.500799783412387e-07
+    4.093895199812102e-07
+ 6.6e+09     
+    4.089941022364158e-07
+     1.50074452797637e-07
+    4.061378313419925e-07
+    4.611817406576593e-08
+    9.296807253394164e-08
+    4.060726188055647e-07
+    2.544640367981455e-08
+    4.611665341719362e-08
+    1.501190189437733e-07
+    4.094182898224932e-07
+ 6.7e+09     
+    4.090236353569304e-07
+    1.501144422866095e-07
+    4.061676979586043e-07
+    4.615650554144875e-08
+    9.300721179722216e-08
+    4.061025258012419e-07
+    2.548237283005278e-08
+    4.615494353477252e-08
+    1.501590097565998e-07
+    4.094482893885663e-07
+ 6.8e+09     
+    4.090543823276525e-07
+    1.501553670606445e-07
+    4.061987564536813e-07
+    4.619577620739048e-08
+    9.304723427360412e-08
+    4.061336244290366e-07
+    2.551925205848422e-08
+    4.619417284776397e-08
+    1.501999359137906e-07
+    4.094794955410699e-07
+ 6.9e+09     
+    4.090863200739828e-07
+     1.50197211766552e-07
+    4.062309824724133e-07
+    4.623595754178163e-08
+    9.308812796307063e-08
+      4.0616589025554e-07
+    2.555701667634095e-08
+    4.623431298985994e-08
+    1.502417820513722e-07
+    4.095118849596264e-07
+ 7e+09       
+    4.091194253778715e-07
+    1.502399605967805e-07
+    4.062643515517032e-07
+    4.627702107721447e-08
+    9.312988048067161e-08
+    4.061992987499885e-07
+    2.559564051739545e-08
+     4.62753356281208e-08
+    1.502845323541574e-07
+    4.095454341927563e-07
+ 7.1e+09     
+    4.091536749229059e-07
+    1.502835973343767e-07
+    4.062988391417628e-07
+    4.631893851463319e-08
+    9.317247905876234e-08
+    4.062338253062354e-07
+    2.563509627723434e-08
+    4.631721257883865e-08
+    1.503281706005506e-07
+    4.095801197051273e-07
+ 7.2e+09     
+    4.091890453361963e-07
+    1.503281053960073e-07
+    4.063344206270744e-07
+    4.636168181765734e-08
+    9.321591054884491e-08
+    4.062694452639319e-07
+    2.567535582485402e-08
+    4.635991590371834e-08
+     1.50372680205415e-07
+    4.096159179212484e-07
+ 7.3e+09     
+     4.09225513227173e-07
+    1.503734678731384e-07
+    4.063710713469844e-07
+    4.640522328977838e-08
+    9.326016142371515e-08
+    4.063061339291975e-07
+    2.571639048388156e-08
+     4.64034179888445e-08
+    1.504180442610924e-07
+    4.096528052657544e-07
+ 7.4e+09     
+     4.09263055223445e-07
+    1.504196675714618e-07
+    4.064087666161274e-07
+    4.644953563669083e-08
+    9.330521778048422e-08
+    4.063438665949833e-07
+    2.575817128220942e-08
+    4.644769160867584e-08
+    1.504642455766691e-07
+    4.096907582004434e-07
+ 7.5e+09     
+    4.093016480038708e-07
+    1.504666870486607e-07
+    4.064474817448227e-07
+    4.649459201580439e-08
+    9.335106534493106e-08
+     4.06382618561285e-07
+    2.580066917004663e-08
+    4.649270997710046e-08
+    1.505112667155742e-07
+    4.097297532582552e-07
+ 7.6e+09     
+    4.093412683290212e-07
+    1.505145086505982e-07
+    4.064871920595507e-07
+    4.654036607476662e-08
+    9.339768947753066e-08
+    4.064223651553169e-07
+    2.584385520732878e-08
+     4.65384467873787e-08
+    1.505590900315992e-07
+    4.097697670743768e-07
+ 7.7e+09     
+    4.093818930691949e-07
+    1.505631145460101e-07
+    4.065278729235625e-07
+    4.658683198063408e-08
+    9.344507518140755e-08
+    4.064630817517151e-07
+    2.588770072212457e-08
+    4.658487624261038e-08
+    1.506076977034163e-07
+    4.098107764146785e-07
+ 7.8e+09     
+    4.094234992301695e-07
+    1.506124867597694e-07
+    4.065694997576392e-07
+    4.663396444113976e-08
+    9.349320711237451e-08
+    4.065047437928005e-07
+     2.59321774421494e-08
+    4.663197307817828e-08
+    1.506570717676685e-07
+    4.098527582016644e-07
+ 7.9e+09     
+     4.09466063976852e-07
+    1.506626072047908e-07
+    4.066120480610056e-07
+    4.668173871933467e-08
+    9.354206959114264e-08
+    4.065473268089055e-07
+    2.597725760178579e-08
+     4.66797125774515e-08
+    1.507071941506948e-07
+    4.098956895381357e-07
+ 8e+09       
+    4.095095646549858e-07
+    1.507134577126219e-07
+    4.066554934323488e-07
+    4.673013064271968e-08
+    9.359164661771718e-08
+    4.065908064387412e-07
+    2.602291402714708e-08
+    4.672807058187167e-08
+    1.507580466989438e-07
+     4.09939547728735e-07
+ 8.1e+09     
+    4.095539788110642e-07
+    1.507650200627699e-07
+    4.066998115908974e-07
+    4.677911660783963e-08
+    9.364192188793899e-08
+    4.066351584497625e-07
+    2.606912020174195e-08
+    4.677702349640046e-08
+    1.508096112081211e-07
+    4.099843102995499e-07
+ 8.2e+09     
+    4.095992842105896e-07
+     1.50817276010796e-07
+    4.067449783974861e-07
+    4.682867358117538e-08
+    9.369287881208014e-08
+    4.066803587584695e-07
+     2.61158503152284e-08
+    4.682654829117494e-08
+    1.508618694511066e-07
+    4.100299550159166e-07
+ 8.3e+09     
+    4.096454588548041e-07
+    1.508702073152068e-07
+    4.067909698755239e-07
+    4.687877909705131e-08
+    9.374450053536018e-08
+    4.067263834505783e-07
+    2.616307929761546e-08
+    4.687662250009402e-08
+    1.509148032046701e-07
+    4.100764598985899e-07
+ 8.4e+09     
+    4.096924809960057e-07
+    1.509237957631612e-07
+    4.068377622317759e-07
+    4.692941125316841e-08
+    9.379676996021844e-08
+    4.067732088009722e-07
+    2.621078284109996e-08
+    4.692722421695417e-08
+    1.509683942750069e-07
+    4.101238032383813e-07
+ 8.5e+09     
+    4.097403291515504e-07
+    1.509780231950098e-07
+    4.068853318768631e-07
+    4.698054870427608e-08
+    9.384966977015024e-08
+    4.068208112933618e-07
+    2.625893741153012e-08
+    4.697833208965507e-08
+    1.510226245221077e-07
+    4.101719636094075e-07
+ 8.6e+09     
+    4.097889821166368e-07
+    1.510328715276751e-07
+     4.06933655445379e-07
+    4.703217065441212e-08
+    9.390318245489355e-08
+    4.068691676395518e-07
+    2.630752025128259e-08
+    4.702992531291289e-08
+    1.510774758829763e-07
+    4.102209198810404e-07
+ 8.7e+09     
+    4.098384189759521e-07
+    1.510883227768804e-07
+    4.069827098155319e-07
+    4.708425684806859e-08
+    9.395729033674382e-08
+    4.069182547982351e-07
+    2.635650937513359e-08
+    4.708198361984226e-08
+     1.51132930393701e-07
+    4.102706512286601e-07
+ 8.8e+09     
+    4.098886191142523e-07
+    1.511443590782343e-07
+    4.070324721282128e-07
+    4.713678756057562e-08
+    9.401197559776236e-08
+    4.069680499932281e-07
+    2.640588356050616e-08
+    4.713448727270853e-08
+    1.511889702103876e-07
+    4.103211371432947e-07
+ 8.9e+09     
+    4.099395622259458e-07
+    1.512009627071723e-07
+    4.070829198054021e-07
+    4.718974358794179e-08
+    9.406722030764335e-08
+    4.070185307310572e-07
+    2.645562233328745e-08
+    4.718741705309061e-08
+    1.512455776289568e-07
+    4.103723574402242e-07
+ 9e+09       
+    4.099912283237327e-07
+     1.51258116097762e-07
+    4.071340305678304e-07
+    4.724310623634306e-08
+    9.412300645200678e-08
+    4.070696748178313e-07
+    2.650570595023788e-08
+    4.724075425165388e-08
+    1.513027351038139e-07
+    4.104242922666153e-07
+ 9.1e+09     
+    4.100435977463604e-07
+    1.513158018603783e-07
+    4.071857824518138e-07
+    4.729685731141286e-08
+    9.417931596088833e-08
+    4.071214603753202e-07
+    2.655611537885728e-08
+     4.72944806576883e-08
+    1.513604252653941e-07
+    4.104769221082523e-07
+ 9.2e+09     
+    4.100966511655329e-07
+    1.513740027982518e-07
+    4.072381538252013e-07
+    4.735097910745172e-08
+    9.423613073720851e-08
+    4.071738658561775e-07
+    2.660683227543256e-08
+    4.734857854853653e-08
+    1.514186309365926e-07
+    4.105302277954164e-07
+ 9.3e+09     
+    4.101503695920231e-07
+    1.514327019229045e-07
+    4.072911234023685e-07
+    4.740545439665075e-08
+    9.429343268501347e-08
+     4.07226870058257e-07
+    2.665783896186884e-08
+    4.740303067900519e-08
+     1.51477335148088e-07
+    4.105841905079644e-07
+ 9.4e+09     
+    4.102047343810276e-07
+    1.514918824684806e-07
+    4.073446702582091e-07
+    4.746026641839615e-08
+    9.435120373729601e-08
+    4.072804521379695e-07
+    2.670911840179807e-08
+    4.745782027083518e-08
+    1.515365211525713e-07
+      4.1063879177966e-07
+ 9.5e+09     
+     4.10259727236799e-07
+    1.515515279049893e-07
+    4.073987738410824e-07
+    4.751539886870773e-08
+    9.440942588321931e-08
+    4.073345916226469e-07
+    2.676065417636549e-08
+    4.751293100228207e-08
+    1.515961724378955e-07
+    4.106940135017867e-07
+ 9.6e+09     
+    4.103153302165837e-07
+     1.51611621950475e-07
+    4.074534139846855e-07
+    4.757083588984545e-08
+    9.446808119458403e-08
+    4.073892684218797e-07
+    2.681243046001507e-08
+    4.756834699784688e-08
+    1.516562727391621e-07
+    4.107498379260969e-07
+ 9.7e+09     
+    4.103715257339109e-07
+    1.516721485821379e-07
+    4.075085709188285e-07
+    4.762656206011265e-08
+    9.452715185139992e-08
+    4.074444628378082e-07
+    2.686443199652798e-08
+    4.762405281818373e-08
+    1.517168060497662e-07
+    4.108062476671217e-07
+ 9.8e+09     
+    4.104282965612489e-07
+    1.517330920464252e-07
+    4.075642252790959e-07
+    4.768256238386538e-08
+    9.458662016643636e-08
+     4.07500155574356e-07
+    2.691664407550927e-08
+    4.768003345020094e-08
+    1.517777566314223e-07
+    4.108632257038848e-07
+ 9.9e+09     
+    4.104856258320639e-07
+    1.517944368681214e-07
+    4.076203581153923e-07
+    4.773882228174192e-08
+    9.464646860865137e-08
+    4.075563277453989e-07
+    2.696905250947286e-08
+    4.773627429736629e-08
+     1.51839109023197e-07
+     4.10920755381047e-07
+ 1e+10       
+    4.105434970423134e-07
+    1.518561678584655e-07
+     4.07676950899373e-07
+    4.779532758111034e-08
+    9.470667982541157e-08
+    4.076129608818726e-07
+    2.702164361163332e-08
+    4.779276117022086e-08
+    1.519008480495785e-07
+     4.10978820409516e-07
+ 1.01e+10    
+    4.106018940513929e-07
+    1.519182701223255e-07
+    4.077339855307753e-07
+    4.785206450673752e-08
+    9.476723666343854e-08
+    4.076700369378309e-07
+    2.707440417448178e-08
+    4.784948027709978e-08
+    1.519629588276101e-07
+     4.11037404866548e-07
+ 1.02e+10    
+    4.106608010825639e-07
+    1.519807290644633e-07
+    4.077914443426578e-07
+    4.790901967166982e-08
+    9.482812218842873e-08
+    4.077275382954651e-07
+    2.712732144919635e-08
+     4.79064182150601e-08
+    1.520254267731251e-07
+    4.110964931953747e-07
+ 1.03e+10    
+    4.107202027229009e-07
+    1.520435303949276e-07
+    4.078493101055853e-07
+    4.796618006832695e-08
+    9.488931970331614e-08
+    4.077854477691136e-07
+    2.718038312591675e-08
+    4.796356196100885e-08
+    1.520882376061131e-07
+    4.111560702043745e-07
+ 1.04e+10    
+     4.10780083922759e-07
+     1.52106660133606e-07
+    4.079075660307748e-07
+    4.802353305979488e-08
+    9.495081276515762e-08
+    4.078437486082878e-07
+    2.723357731489474e-08
+    4.802089886302565e-08
+    1.521513773552581e-07
+    4.112161210658241e-07
+ 1.05e+10    
+    4.108404299948143e-07
+    1.521701046139797e-07
+    4.079661957722508e-07
+    4.808106637131548e-08
+    9.501258520063645e-08
+     4.07902424499739e-07
+    2.728689252852028e-08
+    4.807841663187453e-08
+     1.52214832361682e-07
+    4.112766313142489e-07
+ 1.06e+10    
+     4.10901226612678e-07
+    1.522338504861151e-07
+    4.080251834280366e-07
+    4.813876808196186e-08
+    9.507462112019244e-08
+    4.079614595686145e-07
+     2.73403176642109e-08
+    4.813610333269569e-08
+    1.522785892819332e-07
+    4.113375868443972e-07
+ 1.07e+10    
+    4.109624598091233e-07
+    1.522978847189328e-07
+    4.080845135404301e-07
+    4.819662661649455e-08
+    9.513690493079712e-08
+    4.080208383787319e-07
+     2.73938419881462e-08
+    4.819394737687312e-08
+    1.523426350902604e-07
+    4.113989739088693e-07
+ 1.08e+10    
+    4.110241159739395e-07
+    1.523621946017932e-07
+    4.081441710954067e-07
+    4.825463073738814e-08
+    9.519942134740279e-08
+    4.080805459320188e-07
+    2.744745511982117e-08
+    4.825193751406838e-08
+    1.524069570802066e-07
+    4.114607791154133e-07
+ 1.09e+10    
+    4.110861818514417e-07
+    1.524267677454398e-07
+    4.082041415212027e-07
+    4.831276953702557e-08
+     9.52621554031031e-08
+    4.081405676671641e-07
+    2.750114701739022e-08
+     4.83100628244178e-08
+    1.524715428655667e-07
+    4.115229894239205e-07
+ 1.1e+10     
+    4.111486445376545e-07
+    1.524915920823363e-07
+    4.082644106861161e-07
+    4.837103243004916e-08
+    9.532509245804842e-08
+    4.082008894575199e-07
+    2.755490796376862e-08
+    4.836831271088424e-08
+    1.525363803807447e-07
+    4.115855921431346e-07
+ 1.11e+10    
+    4.112114914771957e-07
+    1.525566558664385e-07
+    4.083249648955858e-07
+    4.842940914586769e-08
+    9.538821820716585e-08
+    4.082614976083093e-07
+    2.760872855345833e-08
+    4.842667689175947e-08
+    1.526014578805492e-07
+     4.11648574927102e-07
+ 1.12e+10    
+    4.112747104598761e-07
+    1.526219476724379e-07
+    4.083857908885954e-07
+    4.848788972131008e-08
+    9.545151868673858e-08
+    4.083223788531812e-07
+    2.766259968006294e-08
+    4.848514539331417e-08
+    1.526667639394661e-07
+    4.117119257713752e-07
+ 1.13e+10    
+    4.113382896170397e-07
+    1.526874563945161e-07
+    4.084468758334531e-07
+    4.854646449342542e-08
+     9.55149802799016e-08
+    4.083835203501646e-07
+    2.771651252445698e-08
+    4.854370854258851e-08
+    1.527322874504437e-07
+    4.117756330089999e-07
+ 1.14e+10    
+    4.114022174176651e-07
+    1.527531712446437e-07
+    4.085082073229958e-07
+    4.860512409242154e-08
+    9.557858972111363e-08
+    4.084449096770658e-07
+    2.777045854357465e-08
+    4.860235696032256e-08
+    1.527980176232276e-07
+    4.118396853062939e-07
+ 1.15e+10    
+    4.114664826642429e-07
+    1.528190817504601e-07
+    4.085697733692694e-07
+    4.866385943474172e-08
+    9.564233409966507e-08
+    4.085065348263604e-07
+     2.78244294597837e-08
+     4.86610815540205e-08
+    1.528639439822787e-07
+    4.119040716584415e-07
+ 1.16e+10    
+    4.115310744884541e-07
+      1.5288517775277e-07
+    4.086315623977377e-07
+    4.872266171627429e-08
+    9.570620086228562e-08
+    4.085683841996211e-07
+    2.787841725081196e-08
+    4.871987351114947e-08
+    1.529300563643091e-07
+    4.119687813849228e-07
+ 1.17e+10    
+    4.115959823466641e-07
+    1.529514494026847e-07
+    4.086935632410553e-07
+    4.878152240569507e-08
+    9.577017781490989e-08
+    4.086304466015305e-07
+    2.793241414019399e-08
+    4.877872429246702e-08
+    1.529963449154673e-07
+    4.120338041247869e-07
+ 1.18e+10    
+    4.116611960152454e-07
+     1.53017887158444e-07
+    4.087557651324654e-07
+    4.884043323793721e-08
+    9.583425312366283e-08
+    4.086927112335197e-07
+    2.798641258820753e-08
+    4.883762562547789e-08
+    1.530628000882036e-07
+    4.120991298317938e-07
+ 1.19e+10    
+    4.117267055857602e-07
+    1.530844817819457e-07
+    4.088181576988567e-07
+    4.889938620778824e-08
+    9.589841531512161e-08
+    4.087551676870735e-07
+    2.804040528327052e-08
+    4.889656949801538e-08
+    1.531294126378458e-07
+    4.121647487694333e-07
+ 1.2e+10     
+    4.117925014600003e-07
+    1.531512243350112e-07
+     4.08880730953522e-07
+    4.895837356361285e-08
+    9.596265327591249e-08
+    4.088178059367495e-07
+    2.809438513377105e-08
+    4.895554815194911e-08
+    1.531961736189122e-07
+    4.122306515058406e-07
+ 1.21e+10    
+    4.118585743449126e-07
+    1.532181061754156e-07
+    4.089434752886655e-07
+    4.901738780119718e-08
+    9.602695625169394e-08
+    4.088806163329398e-07
+    2.814834526030374e-08
+    4.901455407701339e-08
+    1.532630743811885e-07
+    4.122968289086181e-07
+ 1.22e+10    
+    4.119249152474234e-07
+    1.532851189527055e-07
+    4.090063814676881e-07
+    4.907642165771596e-08
+    9.609131384557966e-08
+    4.089435895944168e-07
+    2.820227898828822e-08
+    4.907358000475782e-08
+    1.533301065655944e-07
+    4.123632721395784e-07
+ 1.23e+10    
+     4.11991515469169e-07
+    1.533522546038293e-07
+     4.09069440617293e-07
+    4.913546810581758e-08
+    9.615571601604802e-08
+    4.090067168006977e-07
+    2.825617984094609e-08
+    4.913261890261735e-08
+     1.53397262099863e-07
+    4.124299726494242e-07
+ 1.24e+10    
+     4.12058366601153e-07
+     1.53419505348602e-07
+    4.091326442194426e-07
+    4.919452034782817e-08
+    9.622015307438515e-08
+    4.090699893842594e-07
+    2.831004153261443e-08
+    4.919166396809923e-08
+    1.534645331940529e-07
+    4.124969221723684e-07
+ 1.25e+10    
+     4.12125460518339e-07
+     1.53486863685026e-07
+    4.091959841031992e-07
+    4.925357181007178e-08
+    9.628461568170228e-08
+    4.091333991226319e-07
+     2.83638579623757e-08
+    4.925070862308747e-08
+    1.535319123359184e-07
+    4.125641127207153e-07
+ 1.26e+10    
+    4.121927893741902e-07
+    1.535543223844852e-07
+    4.092594524364763e-07
+    4.931261613730428e-08
+    9.634909484556752e-08
+    4.091969381304006e-07
+    2.841762320798431e-08
+    4.930974650826045e-08
+    1.535993922861516e-07
+    4.126315365794059e-07
+ 1.27e+10    
+    4.122603455951746e-07
+    1.536218744868346e-07
+    4.093230417177313e-07
+    4.937164718726064e-08
+    9.641358191628886e-08
+    4.092605988511432e-07
+    2.847133152007225e-08
+    4.936877147762258e-08
+    1.536669660735186e-07
+    4.126991863005422e-07
+ 1.28e+10    
+    4.123281218752314e-07
+    1.536895132953967e-07
+    4.093867447676226e-07
+    4.943065902531303e-08
+    9.647806858288098e-08
+    4.093243740493262e-07
+    2.852497731661687e-08
+    4.942777759314728e-08
+    1.537346269899035e-07
+    4.127670546978951e-07
+ 1.29e+10    
+    4.123961111702256e-07
+    1.537572323718852e-07
+    4.094505547206527e-07
+    4.948964591923795e-08
+    9.654254686874649e-08
+    4.093882568021811e-07
+    2.857855517765491e-08
+    4.948675911952746e-08
+    1.538023685852774e-07
+    4.128351348414091e-07
+ 1.3e+10     
+    4.124643066923876e-07
+    1.538250255312672e-07
+    4.095144650168236e-07
+    4.954860233409005e-08
+    9.660700912710009e-08
+    4.094522404915791e-07
+    2.863205984022828e-08
+    4.954571051903597e-08
+     1.53870184662605e-07
+    4.129034200517093e-07
+ 1.31e+10    
+    4.125327019047519e-07
+    1.538928868365785e-07
+    4.095784693933146e-07
+     4.96075229271818e-08
+    9.667144803616009e-08
+    4.095163187959306e-07
+    2.868548619354804e-08
+    4.960462644648995e-08
+    1.539380692727041e-07
+    4.129719038946168e-07
+ 1.32e+10    
+    4.126012905156066e-07
+    1.539608105937035e-07
+    4.096425618762084e-07
+    4.966640254316659e-08
+    9.673585659413167e-08
+    4.095804856821166e-07
+     2.87388292743636e-08
+     4.96635017443192e-08
+    1.540060167090672e-07
+    4.130405801756839e-07
+ 1.33e+10    
+    4.126700664729481e-07
+     1.54028791346131e-07
+    4.097067367722774e-07
+     4.97252362092222e-08
+    9.680022811400136e-08
+    4.096447353974754e-07
+    2.879208426252508e-08
+    4.972233143773668e-08
+    1.540740215026583e-07
+    4.131094429347509e-07
+ 1.34e+10    
+    4.127390239589665e-07
+    1.540968238696968e-07
+    4.097709886608421e-07
+    4.978401913033421e-08
+    9.686455621816239e-08
+    4.097090624618493e-07
+    2.884524647672838e-08
+     4.97811107300081e-08
+    1.541420784166952e-07
+    4.131784864405359e-07
+ 1.35e+10    
+    4.128081573845527e-07
+    1.541649031673205e-07
+    4.098353123857204e-07
+    4.984274668467645e-08
+    9.692883483288856e-08
+     4.09773461659715e-07
+    2.889831137043173e-08
+    4.983983499781931e-08
+    1.542101824414241e-07
+    4.132477051852541e-07
+ 1.36e+10    
+    4.128774613838419e-07
+    1.542330244637477e-07
+    4.098997030472696e-07
+    4.990141441908651e-08
+    9.699305818267069e-08
+    4.098379280323984e-07
+    2.895127452793475e-08
+    4.989849978673894e-08
+    1.542783287888981e-07
+     4.13317093879285e-07
+ 1.37e+10    
+    4.129469308087969e-07
+    1.543011832003031e-07
+    4.099641559945404e-07
+    4.996001804463402e-08
+    9.705722078443182e-08
+    4.099024568703893e-07
+    2.900413166061075e-08
+     4.99571008067755e-08
+    1.543465128877648e-07
+    4.133866474458786e-07
+ 1.38e+10    
+    4.130165607238333e-07
+    1.543693750296612e-07
+     4.10028666817542e-07
+    5.001855343228084e-08
+    9.712131744163193e-08
+    4.099670437057591e-07
+    2.905687860328374e-08
+    5.001563392802447e-08
+    1.544147303780711e-07
+    4.134563610159142e-07
+ 1.39e+10    
+    4.130863464004969e-07
+    1.544375958106444e-07
+    4.100932313396359e-07
+    5.007701660862914e-08
+    9.718534323827662e-08
+    4.100316843046985e-07
+    2.910951131074239e-08
+    5.007409517640638e-08
+     1.54482977106092e-07
+    4.135262299227112e-07
+ 1.4e+10     
+    4.131562833121948e-07
+    1.545058416030501e-07
+    4.101578456100552e-07
+    5.013540375175802e-08
+    9.724929353283816e-08
+    4.100963746601692e-07
+    2.916202585438392e-08
+    5.013248072949166e-08
+     1.54551249119187e-07
+    4.135962496968988e-07
+ 1.41e+10    
+    4.132263671289812e-07
+     1.54574108662514e-07
+     4.10222505896559e-07
+    5.019371118714377e-08
+    9.731316395210085e-08
+    4.101611109846858e-07
+     2.92144184189804e-08
+    5.019078691241097e-08
+    1.546195426606934e-07
+    4.136664160613442e-07
+ 1.42e+10    
+    4.132965937124081e-07
+    1.546423934354144e-07
+    4.102872086782269e-07
+    5.025193538366502e-08
+    9.737695038493935e-08
+    4.102258897032227e-07
+    2.926668529956174e-08
+     5.02490101938497e-08
+    1.546878541648553e-07
+    4.137367249261437e-07
+ 1.43e+10    
+     4.13366959110438e-07
+    1.547106925538225e-07
+     4.10351950638398e-07
+    5.031007294968803e-08
+     9.74406489760401e-08
+     4.10290707446263e-07
+    2.931882289840892e-08
+    5.030714718212453e-08
+    1.547561802517989e-07
+    4.138071723836822e-07
+ 1.44e+10    
+    4.134374595524238e-07
+    1.547790028304989e-07
+    4.104167286577501e-07
+    5.036812062923279e-08
+    9.750425611957266e-08
+    4.103555610429757e-07
+    2.937082772215206e-08
+    5.036519462133949e-08
+    1.548245177225537e-07
+    4.138777547037572e-07
+ 1.45e+10    
+    4.135080914441615e-07
+    1.548473212539455e-07
+    4.104815398075357e-07
+    5.042607529821697e-08
+    9.756776845282163e-08
+    4.104204475145406e-07
+    2.942269637896823e-08
+    5.042314938762154e-08
+    1.548928635541239e-07
+    4.139484683287787e-07
+ 1.46e+10    
+    4.135788513630106e-07
+    1.549156449835101e-07
+    4.105463813429587e-07
+    5.048393396077601e-08
+    9.763118284978396e-08
+    4.104853640676079e-07
+    2.947442557587351e-08
+    5.048100848543194e-08
+    1.549612148946142e-07
+    4.140193098690323e-07
+ 1.47e+10    
+    4.136497360530923e-07
+    1.549839713445504e-07
+    4.106112506967068e-07
+      5.0541693745659e-08
+    9.769449641474284e-08
+    4.105503080879077e-07
+    2.952601211610563e-08
+    5.053876904395395e-08
+    1.550295690584123e-07
+    4.140902760980261e-07
+ 1.48e+10    
+    4.137207424205643e-07
+     1.55052297823659e-07
+    4.106761454726366e-07
+    5.059935190269738e-08
+    9.775770647582319e-08
+    4.106152771339974e-07
+    2.957745289659202e-08
+    5.059642831355414e-08
+    1.550979235214298e-07
+    4.141613639479058e-07
+ 1.49e+10    
+    4.137918675289676e-07
+    1.551206220639503e-07
+    4.107410634396058e-07
+    5.065690579934602e-08
+    9.782081057853777e-08
+    4.106802689311584e-07
+    2.962874490549965e-08
+    5.065398366231604e-08
+    1.551662759164056e-07
+    4.142325705049499e-07
+ 1.5e+10     
+    4.138631085946608e-07
+    1.551889418604128e-07
+    4.108060025254641e-07
+    5.071435291729575e-08
+    9.788380647932982e-08
+    4.107452813654355e-07
+    2.967988521986284e-08
+    5.071143257264504e-08
+    1.552346240282708e-07
+     4.14303893005139e-07
+ 1.51e+10    
+    4.139344629823253e-07
+    1.552572551553277e-07
+    4.108709608111872e-07
+    5.077169084915491e-08
+    9.794669213912096e-08
+    4.108103124778211e-07
+    2.973087100328549e-08
+    5.076877263794352e-08
+     1.55302965789581e-07
+    4.143753288298067e-07
+ 1.52e+10    
+      4.1400592820056e-07
+    1.553255600337562e-07
+    4.109359365251683e-07
+    5.082891729519929e-08
+    9.800946571687075e-08
+    4.108753604585855e-07
+    2.978169950371421e-08
+     5.08260015593548e-08
+    1.553712992760141e-07
+    4.144468755013675e-07
+ 1.53e+10    
+    4.140775018975491e-07
+    1.553938547190956e-07
+     4.11000928037656e-07
+    5.088603006018969e-08
+    9.807212556315479e-08
+    4.109404236417475e-07
+    2.983236805127925e-08
+     5.08831171425741e-08
+    1.554396227019364e-07
+    4.145185306791231e-07
+ 1.54e+10    
+    4.141491818568201e-07
+     1.55462137568707e-07
+    4.110659338553411e-07
+     5.09430270502564e-08
+    9.813467021376915e-08
+    4.110055004996915e-07
+    2.988287405620073e-08
+    5.094011729472698e-08
+    1.555079344160392e-07
+    4.145902921551521e-07
+ 1.55e+10    
+    4.142209659930788e-07
+    1.555304070696148e-07
+    4.111309526160905e-07
+    5.099990626984772e-08
+     9.81970983833674e-08
+    4.110705896379233e-07
+     2.99332150067565e-08
+    5.099700002131293e-08
+    1.555762328970445e-07
+    4.146621578502741e-07
+ 1.56e+10    
+    4.142928523481292e-07
+    1.555986618342783e-07
+    4.111959830838282e-07
+    5.105666581874439e-08
+    9.825940895913746e-08
+    4.111356897899679e-07
+    2.998338846730991e-08
+     5.10537634232137e-08
+    1.556445167494842e-07
+    4.147341258100998e-07
+ 1.57e+10    
+    4.143648390868772e-07
+    1.556669005964379e-07
+    4.112610241435552e-07
+    5.111330388913599e-08
+    9.832160099452475e-08
+    4.112007998124044e-07
+    3.003339207639433e-08
+    5.111040569376543e-08
+    1.557127846995502e-07
+    4.148061942011559e-07
+ 1.58e+10    
+    4.144369244934146e-07
+     1.55735122207035e-07
+    4.113260747965182e-07
+    5.116981876276157e-08
+    9.838367370300853e-08
+    4.112659186800411e-07
+    3.008322354485264e-08
+    5.116692511589402e-08
+    1.557810355910191e-07
+    4.148783613070942e-07
+ 1.59e+10    
+    4.145091069671897e-07
+    1.558033256302074e-07
+    4.113911341555131e-07
+    5.122620880811123e-08
+    9.844562645193775e-08
+    4.113310454812238e-07
+      3.0132880654029e-08
+    5.122332005931227e-08
+    1.558492683812501e-07
+    4.149506255249786e-07
+ 1.6e+10     
+    4.145813850192561e-07
+    1.558715099393595e-07
+    4.114562014403281e-07
+    5.128247247768878e-08
+    9.850745875643207e-08
+    4.113961794132769e-07
+    3.018236125401118e-08
+    5.127958897777855e-08
+    1.559174821372571e-07
+     4.15022985361649e-07
+ 1.61e+10    
+    4.146537572686082e-07
+    1.559396743133083e-07
+    4.115212759733207e-07
+    5.133860830533576e-08
+    9.856917027335566e-08
+    4.114613197780797e-07
+    3.023166326192124e-08
+    5.133573040641578e-08
+    1.559856760318564e-07
+    4.150954394301688e-07
+ 1.62e+10    
+    4.147262224385943e-07
+    1.560078180325067e-07
+    4.115863571751326e-07
+    5.139461490361415e-08
+    9.863076079536786e-08
+    4.115264659777701e-07
+    3.028078466025311e-08
+    5.139174295909133e-08
+    1.560538493398897e-07
+    4.151679864463488e-07
+ 1.63e+10    
+    4.147987793534145e-07
+    1.560759404753416e-07
+    4.116514445605317e-07
+    5.145049096124815e-08
+    9.869223024505748e-08
+    4.115916175105761e-07
+    3.032972349525455e-08
+    5.144762532585465e-08
+    1.561220014345217e-07
+    4.152406252253479e-07
+ 1.64e+10    
+    4.148714269346962e-07
+    1.561440411145091e-07
+     4.11716537734383e-07
+     5.15062352406253e-08
+    9.875357866916569e-08
+    4.116567739667737e-07
+    3.037847787535279e-08
+    5.150337627043479e-08
+    1.561901317836139e-07
+    4.153133546783531e-07
+ 1.65e+10    
+     4.14944164198154e-07
+    1.562121195134667e-07
+    4.117816363877501e-07
+    5.156184657535394e-08
+    9.881480623290297e-08
+    4.117219350247684e-07
+    3.042704596962144e-08
+    5.155899462779471e-08
+    1.562582399461747e-07
+    4.153861738093348e-07
+ 1.66e+10    
+    4.150169902503231e-07
+    1.562801753229607e-07
+    4.118467402941148e-07
+    5.161732386787864e-08
+    9.887591321436405e-08
+    4.117871004472976e-07
+    3.047542600628777e-08
+    5.161447930174386e-08
+    1.563263255688844e-07
+    4.154590817118801e-07
+ 1.67e+10    
+    4.150899042853767e-07
+    1.563482082776319e-07
+    4.119118493057249e-07
+    5.167266608715157e-08
+    9.893689999904653e-08
+     4.11852270077751e-07
+    3.052361627127847e-08
+    5.166982926260605e-08
+    1.563943883826965e-07
+    4.155320775660979e-07
+ 1.68e+10    
+     4.15162905582017e-07
+    1.564162181926952e-07
+    4.119769633500543e-07
+    5.172787226635983e-08
+     9.89977670744765e-08
+    4.119174438366109e-07
+    3.057161510680302e-08
+    5.172504354494426e-08
+    1.564624281995151e-07
+    4.156051606356023e-07
+ 1.69e+10    
+    4.152359935004453e-07
+     1.56484204960698e-07
+    4.120420824263872e-07
+    5.178294150070735e-08
+    9.905851502494551e-08
+    4.119826217180032e-07
+    3.061942090997292e-08
+    5.178012124534035e-08
+    1.565304449089465e-07
+     4.15678330264567e-07
+ 1.7e+10     
+    4.153091674794079e-07
+    1.565521685483518e-07
+    4.121072066025109e-07
+    5.183787294525195e-08
+    9.911914452636174e-08
+    4.120478037863617e-07
+    3.066703213145597e-08
+     5.18350615202292e-08
+    1.565984384751271e-07
+    4.157515858748529e-07
+ 1.71e+10    
+    4.153824270333163e-07
+    1.566201089934407e-07
+    4.121723360115207e-07
+    5.189266581279572e-08
+    9.917965634121987e-08
+    4.121129901732055e-07
+    3.071444727416417e-08
+    5.188986358378681e-08
+    1.566664089336266e-07
+    4.158249269632074e-07
+ 1.72e+10    
+      4.1545577174944e-07
+    1.566880264018048e-07
+     4.12237470848739e-07
+    5.194731937182818e-08
+    9.924005131369076e-08
+    4.121781810740168e-07
+    3.076166489197424e-08
+     5.19445267058717e-08
+    1.567343563884241e-07
+    4.158983530985347e-07
+ 1.73e+10    
+     4.15529201285175e-07
+    1.567559209443979e-07
+    4.123026113687368e-07
+    5.200183294452277e-08
+    9.930033036483545e-08
+    4.122433767452315e-07
+    3.080868358847974e-08
+      5.1999050210019e-08
+    1.568022810089607e-07
+    4.159718639192352e-07
+ 1.74e+10    
+    4.156027153653817e-07
+    1.568237928544194e-07
+     4.12367757882459e-07
+     5.20562059047843e-08
+    9.936049448794344e-08
+    4.123085775013268e-07
+    3.085550201577381e-08
+     5.20534334714862e-08
+    1.568701830272636e-07
+     4.16045459130616e-07
+ 1.75e+10    
+    4.156763137797937e-07
+    1.568916424245196e-07
+    4.124329107544549e-07
+    5.211043767634741e-08
+    9.942054474399926e-08
+    4.123737837120124e-07
+    3.090211887326133e-08
+    5.210767591535026e-08
+    1.569380627351455e-07
+    4.161191385023636e-07
+ 1.76e+10    
+    4.157499963804987e-07
+    1.569594700040786e-07
+    4.124980704002058e-07
+    5.216452773092603e-08
+    9.948048225727696e-08
+    4.124389957995177e-07
+    3.094853290650008e-08
+    5.216177701465476e-08
+    1.570059204814746e-07
+     4.16192901866091e-07
+ 1.77e+10    
+    4.158237630794831e-07
+    1.570272759965561e-07
+    4.125632372835488e-07
+     5.22184755864119e-08
+    9.954030821106488e-08
+    4.125042142359745e-07
+    3.099474290606947e-08
+     5.22157362886075e-08
+     1.57073756669518e-07
+    4.162667491129421e-07
+ 1.78e+10    
+    4.158976138462497e-07
+    1.570950608569149e-07
+    4.126284119141981e-07
+    5.227228080512196e-08
+    9.960002384352129e-08
+    4.125694395408951e-07
+    3.104074770646634e-08
+     5.22695533008264e-08
+    1.571415717543564e-07
+    4.163406801912671e-07
+ 1.79e+10    
+    4.159715487054953e-07
+    1.571628250891133e-07
+    4.126935948453542e-07
+    5.232594299209391e-08
+    9.965963044366104e-08
+    4.126346722787392e-07
+     3.10865461850271e-08
+    5.232322765763391e-08
+    1.572093662403684e-07
+    4.164146951043587e-07
+ 1.8e+10     
+    4.160455677348574e-07
+    1.572305692436681e-07
+    4.127587866714046e-07
+    5.237946179342955e-08
+    9.971912934747357e-08
+    4.126999130565681e-07
+    3.113213726087514e-08
+    5.237675900639894e-08
+    1.572771406787858e-07
+    4.164887939082486e-07
+ 1.81e+10    
+    4.161196710627245e-07
+    1.572982939152883e-07
+    4.128239880257134e-07
+    5.243283689468413e-08
+      9.9778521934173e-08
+    4.127651625217905e-07
+    3.117751989389308e-08
+    5.243014703392569e-08
+    1.573448956653178e-07
+    4.165629767095689e-07
+ 1.82e+10    
+    4.161938588661059e-07
+     1.57365999740575e-07
+    4.128891995784918e-07
+    5.248606801930139e-08
+    9.983780962257821e-08
+    4.128304213599839e-07
+    3.122269308371886e-08
+    5.248339146488739e-08
+    1.574126318378426e-07
+    4.166372436634715e-07
+ 1.83e+10    
+     4.16268131368567e-07
+      1.5743368739579e-07
+    4.129544220347515e-07
+    5.253915492709442e-08
+    9.989699386762436e-08
+    4.128956902928045e-07
+    3.126765586876544e-08
+    5.253649206030675e-08
+    1.574803498741678e-07
+    4.167115949716056e-07
+ 1.84e+10    
+    4.163424888382204e-07
+    1.575013575946917e-07
+     4.13019656132344e-07
+    5.259209741276985e-08
+    9.995607615700359e-08
+    4.129609700759734e-07
+    3.131240732526286e-08
+    5.258944861607904e-08
+    1.575480504898558e-07
+    4.167860308801549e-07
+ 1.85e+10    
+    4.164169315857802e-07
+    1.575690110864354e-07
+    4.130849026400677e-07
+    5.264489530449593e-08
+    1.000150580079342e-07
+    4.130262614973398e-07
+    3.135694656632272e-08
+       5.264226096154e-08
+    1.576157344361159e-07
+    4.168605516779293e-07
+ 1.86e+10    
+    4.164914599626697e-07
+    1.576366486535381e-07
+    4.131501623558569e-07
+    5.269754846251291e-08
+    1.000739409640566e-07
+    4.130915653750195e-07
+    3.140127274102381e-08
+    5.269492895807529e-08
+    1.576834024977606e-07
+    4.169351576945144e-07
+ 1.87e+10    
+    4.165660743591896e-07
+    1.577042711099088e-07
+     4.13215436105044e-07
+    5.275005677778502e-08
+    1.001327265924559e-07
+    4.131568825556041e-07
+    3.144538503351888e-08
+    5.274745249777264e-08
+    1.577510554912253e-07
+    4.170098492984736e-07
+ 1.88e+10    
+    4.166407752027378e-07
+    1.577718792989394e-07
+    4.132807247386883e-07
+    5.280242017069368e-08
+    1.001914164808072e-07
+    4.132222139124437e-07
+    3.148928266216155e-08
+    5.279983150211412e-08
+    1.578186942626507e-07
+    4.170846268956036e-07
+ 1.89e+10    
+    4.167155629560883e-07
+    1.578394740916587e-07
+    4.133460291319764e-07
+    5.285463858977052e-08
+    1.002500122346439e-07
+    4.132875603439952e-07
+    3.153296487865342e-08
+    5.285206592070965e-08
+    1.578863196860273e-07
+    4.171594909272438e-07
+ 1.9e+10     
+    4.167904381157171e-07
+    1.579070563849451e-07
+    4.134113501826888e-07
+    5.290671201046964e-08
+    1.003085154747451e-07
+    4.133529227722364e-07
+    3.157643096720987e-08
+    5.290415573006821e-08
+     1.57953932661399e-07
+    4.172344418686324e-07
+ 1.91e+10    
+     4.16865401210184e-07
+    1.579746270998011e-07
+    4.134766888097288e-07
+    5.295864043397775e-08
+    1.003669278346412e-07
+    4.134183021411469e-07
+    3.161968024374522e-08
+    5.295610093240894e-08
+    1.580215341131278e-07
+    4.173094802273191e-07
+ 1.92e+10    
+    4.169404527985644e-07
+     1.58042187179684e-07
+    4.135420459517161e-07
+    5.301042388606284e-08
+    1.004252509582344e-07
+    4.134836994152463e-07
+    3.166271205507599e-08
+    5.300790155450886e-08
+    1.580891249882155e-07
+    4.173846065416192e-07
+ 1.93e+10    
+    4.170155934689295e-07
+    1.581097375888947e-07
+    4.136074225656385e-07
+    5.306206241595828e-08
+    1.004834864975334e-07
+    4.135491155781966e-07
+    3.170552577814202e-08
+    5.305955764658782e-08
+    1.581567062546829e-07
+    4.174598213791215e-07
+ 1.94e+10    
+    4.170908238368742e-07
+    1.581772793110224e-07
+    4.136728196255602e-07
+    5.311355609528313e-08
+    1.005416361104962e-07
+    4.136145516314579e-07
+    3.174812081924497e-08
+    5.311106928122869e-08
+    1.582242789000054e-07
+    4.175351253352391e-07
+ 1.95e+10    
+    4.171661445440962e-07
+    1.582448133474443e-07
+    4.137382381213902e-07
+    5.316490501699801e-08
+    1.005997014589827e-07
+    4.136800085930048e-07
+    3.179049661330399e-08
+    5.316243655233322e-08
+    1.582918439296032e-07
+    4.176105190318065e-07
+ 1.96e+10    
+    4.172415562570152e-07
+    1.583123407158789e-07
+    4.138036790577003e-07
+    5.321610929439375e-08
+    1.006576842068111e-07
+     4.13745487496093e-07
+    3.183265262312781e-08
+    5.321365957411155e-08
+    1.583594023653854e-07
+    4.176860031157232e-07
+ 1.97e+10    
+    4.173170596654416e-07
+     1.58379862448991e-07
+    4.138691434525976e-07
+    5.326716906011466e-08
+    1.007155860179171e-07
+    4.138109893880781e-07
+    3.187458833870297e-08
+    5.326473848010505e-08
+    1.584269552443465e-07
+    4.177615782576376e-07
+ 1.98e+10    
+    4.173926554812879e-07
+    1.584473795930502e-07
+    4.139346323366462e-07
+    5.331808446521276e-08
+    1.007734085546113e-07
+    4.138765153292855e-07
+    3.191630327649792e-08
+    5.331567342224189e-08
+     1.58494503617214e-07
+     4.17837245150674e-07
+ 1.99e+10    
+    4.174683444373212e-07
+    1.585148932066369e-07
+    4.140001467518353e-07
+    5.336885567823483e-08
+    1.008311534759346e-07
+    4.139420663919293e-07
+    3.195779697878256e-08
+    5.336646456992383e-08
+    1.585620485471473e-07
+    4.179130045092045e-07
+ 2e+10       
+    4.175441272859599e-07
+    1.585824043593996e-07
+    4.140656877505978e-07
+    5.341948288433946e-08
+    1.008888224361056e-07
+    4.140076436590745e-07
+    3.199906901296267e-08
+    5.341711210914424e-08
+     1.58629591108485e-07
+    4.179888570676564e-07
+ 2.01e+10    
+    4.176200047981087e-07
+    1.586499141308588e-07
+     4.14131256394869e-07
+    5.346996628444411e-08
+    1.009464170830596e-07
+    4.140732482236474e-07
+    3.204011897092907e-08
+     5.34676162416354e-08
+    1.586971323855397e-07
+     4.18064803579361e-07
+ 2.02e+10    
+    4.176959777620353e-07
+    1.587174236092574e-07
+    4.141968537551901e-07
+    5.352030609440142e-08
+    1.010039390570744e-07
+     4.14138881187488e-07
+    3.208094646842119e-08
+    5.351797718404586e-08
+    1.587646734714409e-07
+     4.18140844815442e-07
+ 2.03e+10    
+    4.177720469822851e-07
+    1.587849338904586e-07
+    4.142624809098545e-07
+    5.357050254420368e-08
+    1.010613899894816e-07
+    4.142045436604403e-07
+    3.212155114440452e-08
+    5.356819516714526e-08
+    1.588322154670217e-07
+    4.182169815637387e-07
+ 2.04e+10    
+    4.178482132786306e-07
+    1.588524460768844e-07
+    4.143281389440889e-07
+    5.362055587721509e-08
+    1.011187715014586e-07
+    4.142702367594887e-07
+    3.216193266046185e-08
+    5.361827043505743e-08
+    1.588997594797514e-07
+    4.182932146277678e-07
+ 2.05e+10    
+    4.179244774850616e-07
+    1.589199612765012e-07
+    4.143938289492756e-07
+    5.367046634943042e-08
+    1.011760852028999e-07
+    4.143359616079265e-07
+    3.220209070019766e-08
+    5.366820324451965e-08
+    1.589673066227107e-07
+    4.183695448257192e-07
+ 2.06e+10    
+    4.180008404488104e-07
+    1.589874806018453e-07
+    4.144595520222128e-07
+    5.372023422875941e-08
+    1.012333326913646e-07
+    4.144017193345641e-07
+    3.224202496865585e-08
+    5.371799386416843e-08
+    1.590348580136095e-07
+    4.184459729894867e-07
+ 2.07e+10    
+    4.180773030294066e-07
+    1.590550051690888e-07
+    4.145253092644016e-07
+    5.376985979433751e-08
+    1.012905155510958e-07
+    4.144675110729724e-07
+    3.228173519174998e-08
+    5.376764257385026e-08
+    1.591024147738449e-07
+    4.185224999637349e-07
+ 2.08e+10    
+    4.181538660977736e-07
+    1.591225360971475e-07
+    4.145911017813758e-07
+    5.381934333585979e-08
+    1.013476353521113e-07
+    4.145333379607576e-07
+    3.232122111570611e-08
+     5.38171496639569e-08
+    1.591699780275999e-07
+    4.185991266049939e-07
+ 2.09e+10    
+    4.182305305353503e-07
+    1.591900745068246e-07
+    4.146569306820584e-07
+     5.38686851529393e-08
+    1.014046936493604e-07
+    4.145992011388712e-07
+    3.236048250651766e-08
+    5.386651543478467e-08
+    1.592375489009801e-07
+    4.186758537807884e-07
+ 2.1e+10     
+    4.183072972332488e-07
+    1.592576215199943e-07
+    4.147227970781462e-07
+    5.391788555448845e-08
+    1.014616919819464e-07
+    4.146651017509474e-07
+     3.23995191494124e-08
+    5.391574019591633e-08
+    1.593051285211887e-07
+     4.18752682368801e-07
+ 2.11e+10    
+    4.183841670914448e-07
+    1.593251782588204e-07
+    4.147887020835288e-07
+    5.396694485812247e-08
+      1.0151863187241e-07
+    4.147310409426733e-07
+    3.243833084833089e-08
+    5.396482426562611e-08
+    1.593727180157375e-07
+    4.188296132560586e-07
+ 2.12e+10    
+    4.184611410179905e-07
+    1.593927458450104e-07
+    4.148546468137299e-07
+    5.401586338958474e-08
+    1.015755148260719e-07
+    4.147970198611856e-07
+    3.247691742541637e-08
+     5.40137679703053e-08
+     1.59440318511694e-07
+    4.189066473381544e-07
+ 2.13e+10    
+    4.185382199282661e-07
+    1.594603253991044e-07
+    4.149206323853796e-07
+    5.406464148219322e-08
+     1.01632342330433e-07
+     4.14863039654494e-07
+    3.251527872051584e-08
+    5.406257164391022e-08
+    1.595079311349617e-07
+    4.189837855184963e-07
+ 2.14e+10    
+    4.186154047442539e-07
+    1.595279180397965e-07
+    4.149866599157064e-07
+    5.411327947630672e-08
+    1.016891158546265e-07
+    4.149291014709308e-07
+    3.255341459069184e-08
+    5.411123562742936e-08
+    1.595755570095956e-07
+    4.190610287075807e-07
+ 2.15e+10    
+      4.1869269639384e-07
+    1.595955248832889e-07
+    4.150527305220572e-07
+    5.416177771881164e-08
+    1.017458368489236e-07
+    4.149952064586266e-07
+    3.259132490974504e-08
+    5.415976026837057e-08
+    1.596431972571479e-07
+    4.191383778222975e-07
+ 2.16e+10    
+    4.187700958101454e-07
+    1.596631470426767e-07
+    4.151188453214391e-07
+    5.421013656262673e-08
+    1.018025067442869e-07
+    4.150613557650056e-07
+    3.262900956774721e-08
+    5.420814592026796e-08
+    1.597108529960462e-07
+    4.192158337852564e-07
+ 2.17e+10    
+    4.188476039308821e-07
+     1.59730785627363e-07
+    4.151850054300797e-07
+    5.425835636622777e-08
+    1.018591269519714e-07
+    4.151275505363084e-07
+    3.266646847058433e-08
+    5.425639294220623e-08
+    1.597785253410025e-07
+     4.19293397524144e-07
+ 2.18e+10    
+    4.189252216977325e-07
+    1.597984417425034e-07
+    4.152512119630118e-07
+    5.430643749318841e-08
+    1.019156988631683e-07
+    4.151937919171317e-07
+    3.270370153950965e-08
+    5.430450169836366e-08
+    1.598462154024499e-07
+    4.193710699710997e-07
+ 2.19e+10    
+    4.190029500557564e-07
+    1.598661164884774e-07
+    4.153174660336744e-07
+     5.43543803117397e-08
+     1.01972223848693e-07
+    4.152600810499915e-07
+    3.274070871070652e-08
+    5.435247255757193e-08
+     1.59913924286009e-07
+    4.194488520621206e-07
+ 2.2e+10     
+    4.190807899528193e-07
+    1.599338109603894e-07
+    4.153837687535339e-07
+    5.440218519434563e-08
+    1.020287032587117e-07
+    4.153264190749028e-07
+    3.277748993486082e-08
+     5.44003058928931e-08
+    1.599816530919809e-07
+    4.195267447364868e-07
+ 2.21e+10    
+    4.191587423390437e-07
+    1.600015262475933e-07
+    4.154501212317214e-07
+    5.444985251729495e-08
+     1.02085138422506e-07
+    4.153928071289807e-07
+    3.281404517674249e-08
+    5.444800208121212e-08
+    1.600494029148675e-07
+    4.196047489362098e-07
+ 2.22e+10    
+     4.19236808166285e-07
+    1.600692634332442e-07
+    4.155165245746868e-07
+    5.449738266030864e-08
+    1.021415306482738e-07
+    4.154592463460567e-07
+    3.285037441479655e-08
+    5.449556150284547e-08
+    1.601171748429157e-07
+    4.196828656055016e-07
+ 2.23e+10    
+    4.193149883876265e-07
+    1.601370235938741e-07
+    4.155829798858685e-07
+    5.454477600616285e-08
+     1.02197881222964e-07
+    4.155257378563145e-07
+    3.288647764074262e-08
+    5.454298454116485e-08
+    1.601849699576887e-07
+    4.197610956902687e-07
+ 2.24e+10    
+    4.193932839568964e-07
+    1.602048077989905e-07
+    4.156494882653765e-07
+    5.459203294032565e-08
+    1.022541914121428e-07
+    4.155922827859371e-07
+    3.292235485918372e-08
+    5.459027158223535e-08
+     1.60252789333659e-07
+    4.198394401376229e-07
+ 2.25e+10    
+    4.194716958282048e-07
+    1.602726171106994e-07
+    4.157160508096921e-07
+    5.463915385060879e-08
+    1.023104624598909e-07
+    4.156588822567755e-07
+    3.295800608722296e-08
+    5.463742301446743e-08
+     1.60320634037825e-07
+    4.199178998954115e-07
+ 2.26e+10    
+    4.195502249555001e-07
+    1.603404525833481e-07
+    4.157826686113765e-07
+    5.468613912683244e-08
+    1.023666955887278e-07
+    4.157255373860243e-07
+    3.299343135408928e-08
+    5.468443922828323e-08
+    1.603885051293504e-07
+    4.199964759117718e-07
+ 2.27e+10    
+    4.196288722921468e-07
+    1.604083152631914e-07
+    4.158493427587973e-07
+    5.473298916050355e-08
+     1.02422891999565e-07
+    4.157922492859184e-07
+     3.30286307007709e-08
+    5.473132061579539e-08
+    1.604564036592235e-07
+    4.200751691346986e-07
+ 2.28e+10    
+    4.197076387905158e-07
+    1.604762061880752e-07
+    4.159160743358593e-07
+    5.477970434450647e-08
+    1.024790528716818e-07
+    4.158590190634372e-07
+    3.306360417965701e-08
+    5.477806757049865e-08
+    1.605243306699386e-07
+    4.201539805116324e-07
+ 2.29e+10    
+    4.197865254015999e-07
+    1.605441263871425e-07
+    4.159828644217527e-07
+     5.48262850728064e-08
+    1.025351793627271e-07
+    4.159258478200231e-07
+     3.30983518541873e-08
+    5.482468048697429e-08
+    1.605922871951961e-07
+    4.202329109890672e-07
+ 2.3e+10     
+    4.198655330746421e-07
+     1.60612076880557e-07
+     4.16049714090708e-07
+    5.487273174016422e-08
+     1.02591272608741e-07
+    4.159927366513137e-07
+     3.31328737985092e-08
+    5.487115976060554e-08
+    1.606602742596217e-07
+    4.203119615121702e-07
+ 2.31e+10    
+    4.199446627567798e-07
+    1.606800586792438e-07
+    4.161166244117602e-07
+     5.49190447418633e-08
+    1.026473337241988e-07
+    4.160596866468807e-07
+    3.316717009714253e-08
+    5.491750578730503e-08
+    1.607282928785042e-07
+    4.203911330244223e-07
+ 2.32e+10    
+    4.200239153927087e-07
+    1.607480727846492e-07
+     4.16183596448526e-07
+    5.496522447344668e-08
+    1.027033638020738e-07
+    4.161266988899847e-07
+     3.32012408446517e-08
+    5.496371896325314e-08
+    1.607963440575509e-07
+    4.204704264672725e-07
+ 2.33e+10    
+    4.201032919243594e-07
+    1.608161201885157e-07
+    4.162506312589833e-07
+    5.501127133046562e-08
+    1.027593639139171e-07
+    4.161937744573346e-07
+      3.3235086145325e-08
+    5.500979968464679e-08
+    1.608644287926592e-07
+    4.205498427798087e-07
+ 2.34e+10    
+    4.201827932905905e-07
+    1.608842018726736e-07
+    4.163177298952635e-07
+    5.505718570823813e-08
+    1.028153351099558e-07
+    4.162609144188631e-07
+    3.326870611286108e-08
+     5.50557483474587e-08
+    1.609325480697056e-07
+    4.206293828984435e-07
+ 2.35e+10    
+    4.202624204268954e-07
+    1.609523188088484e-07
+    4.163848934034496e-07
+    5.510296800161743e-08
+    1.028712784192055e-07
+    4.163281198375045e-07
+    3.330210087006224e-08
+    5.510156534720676e-08
+    1.610007028643487e-07
+    4.207090477566119e-07
+ 2.36e+10    
+    4.203421742651231e-07
+    1.610204719584817e-07
+    4.164521228233822e-07
+    5.514861860477003e-08
+    1.029271948495973e-07
+    4.163953917689865e-07
+    3.333527054853453e-08
+    5.514725107873209e-08
+    1.610688941418487e-07
+    4.207888382844862e-07
+ 2.37e+10    
+    4.204220557332155e-07
+     1.61088662272567e-07
+    4.165194191884684e-07
+    5.519413791096331e-08
+    1.029830853881187e-07
+    4.164627312616276e-07
+    3.336821528839468e-08
+    5.519280593598753e-08
+    1.611371228569001e-07
+    4.208687554087034e-07
+ 2.38e+10    
+    4.205020657549513e-07
+     1.61156890691499e-07
+    4.165867835255032e-07
+    5.523952631236148e-08
+    1.030389510009667e-07
+    4.165301393561433e-07
+    3.340093523798315e-08
+    5.523823031183414e-08
+    1.612053899534787e-07
+    4.209488000521047e-07
+ 2.39e+10    
+     4.20582205249711e-07
+     1.61225158144935e-07
+    4.166542168544899e-07
+    5.528478419983106e-08
+    1.030947926337112e-07
+      4.1659761708546e-07
+    3.343343055358408e-08
+    5.528352459784665e-08
+    1.612736963647012e-07
+    4.210289731334876e-07
+ 2.4e+10     
+    4.206624751322462e-07
+    1.612934655516704e-07
+    4.167217201884733e-07
+    5.532991196275381e-08
+    1.031506112114706e-07
+    4.166651654745367e-07
+    3.346570139915094e-08
+    5.532868918412706e-08
+    1.613420430126984e-07
+    4.211092755673724e-07
+ 2.41e+10    
+     4.20742876312467e-07
+    1.613618138195236e-07
+    4.167892945333694e-07
+    5.537490998884798e-08
+    1.032064076390946e-07
+    4.167327855401907e-07
+    3.349774794603875e-08
+    5.537372445912627e-08
+    1.614104308084993e-07
+    4.211897082637774e-07
+ 2.42e+10    
+    4.208234096952373e-07
+    1.614302038452342e-07
+    4.168569408878076e-07
+    5.541977866399787e-08
+    1.032621828013582e-07
+    4.168004782909344e-07
+    3.352957037274202e-08
+     5.54186308094734e-08
+    1.614788606519272e-07
+    4.212702721280069e-07
+ 2.43e+10    
+    4.209040761801809e-07
+     1.61498636514371e-07
+     4.16924660242974e-07
+    5.546451837208977e-08
+    1.033179375631615e-07
+    4.168682447268163e-07
+    3.356116886463869e-08
+    5.546340861981264e-08
+    1.615473334315072e-07
+     4.21350968060451e-07
+ 2.44e+10    
+    4.209848766615011e-07
+    1.615671127012506e-07
+    4.169924535824585e-07
+    5.550912949485635e-08
+    1.033736727697375e-07
+     4.16936085839266e-07
+     3.35925436137398e-08
+    5.550805827264697e-08
+    1.616158500243838e-07
+    4.214317969563943e-07
+ 2.45e+10    
+    4.210658120278072e-07
+    1.616356332688658e-07
+    4.170603218821079e-07
+    5.555361241172682e-08
+    1.034293892468664e-07
+    4.170040026109499e-07
+    3.362369481844472e-08
+    5.555258014818908e-08
+    1.616844112962486e-07
+    4.215127597058364e-07
+ 2.46e+10    
+    4.211468831619535e-07
+    1.617041990688234e-07
+     4.17128266109883e-07
+    5.559796749968482e-08
+    1.034850878010956e-07
+    4.170719960156278e-07
+    3.365462268330214e-08
+    5.559697462421903e-08
+    1.617530181012778e-07
+    4.215938571933204e-07
+ 2.47e+10    
+     4.21228090940886e-07
+    1.617728109412913e-07
+    4.171962872257154e-07
+    5.564219513313217e-08
+    1.035407692199643e-07
+    4.171400670180186e-07
+    3.368532741877617e-08
+    5.564124207594783e-08
+    1.618216712820789e-07
+    4.216750902977732e-07
+ 2.48e+10    
+    4.213094362354985e-07
+    1.618414697149526e-07
+    4.172643861813747e-07
+    5.568629568375905e-08
+    1.035964342722334e-07
+    4.172082165736708e-07
+    3.371580924101792e-08
+    5.568538287588783e-08
+    1.618903716696461e-07
+    4.217564598923527e-07
+ 2.49e+10    
+    4.213909199104999e-07
+    1.619101762069708e-07
+    4.173325639203328e-07
+    5.573026952042044e-08
+    1.036520837081189e-07
+    4.172764456288336e-07
+    3.374606837164233e-08
+    5.572939739372865e-08
+    1.619591200833236e-07
+    4.218379668443057e-07
+ 2.5e+10     
+     4.21472542824286e-07
+    1.619789312229589e-07
+    4.174008213776359e-07
+     5.57741170090178e-08
+    1.037077182595287e-07
+    4.173447551203422e-07
+    3.377610503750995e-08
+    5.577328599621902e-08
+    1.620279173307783e-07
+    4.219196120148333e-07
+ 2.51e+10    
+    4.215543058288225e-07
+    1.620477355569602e-07
+    4.174691594797768e-07
+    5.581783851238706e-08
+    1.037633386403025e-07
+    4.174131459754976e-07
+    3.380591947051383e-08
+     5.58170490470544e-08
+    1.620967642079778e-07
+    4.220013962589639e-07
+ 2.52e+10    
+    4.216362097695356e-07
+     1.62116589991432e-07
+    4.175375791445742e-07
+    5.586143439019162e-08
+    1.038189455464548e-07
+    4.174816191119602e-07
+    3.383551190737134e-08
+    5.586068690676955e-08
+    1.621656614991784e-07
+    4.220833204254376e-07
+ 2.53e+10    
+    4.217182554852088e-07
+    1.621854952972386e-07
+    4.176060812810487e-07
+    5.590490499882073e-08
+    1.038745396564183e-07
+    4.175501754376414e-07
+    3.386488258942052e-08
+    5.590419993263671e-08
+    1.622346099769173e-07
+    4.221653853565916e-07
+ 2.54e+10    
+    4.218004438078867e-07
+      1.6225445223365e-07
+    4.176746667893101e-07
+    5.594825069129262e-08
+     1.03930121631291e-07
+    4.176188158506052e-07
+    3.389403176242158e-08
+    5.594758847856834e-08
+    1.623036104020134e-07
+    4.222475918882618e-07
+ 2.55e+10    
+    4.218827755627886e-07
+    1.623234615483458e-07
+    4.177433365604386e-07
+    5.599147181716305e-08
+    1.039856921150831e-07
+    4.176875412389689e-07
+    3.392295967636255e-08
+    5.599085289502499e-08
+     1.62372663523573e-07
+    4.223299408496816e-07
+ 2.56e+10    
+     4.21965251568228e-07
+     1.62392523977427e-07
+    4.178120914763792e-07
+    5.603456872243815e-08
+    1.040412517349652e-07
+    4.177563524808124e-07
+     3.39516665852699e-08
+      5.6033993528928e-08
+    1.624417700790023e-07
+    4.224124330633965e-07
+ 2.57e+10    
+    4.220478726355346e-07
+    1.624616402454297e-07
+    4.178809324098293e-07
+    5.607754174949183e-08
+    1.040968011015177e-07
+    4.178252504440926e-07
+     3.39801527470231e-08
+    5.607701072357599e-08
+    1.625109307940252e-07
+    4.224950693451797e-07
+ 2.58e+10    
+    4.221306395689878e-07
+    1.625308110653478e-07
+    4.179498602241371e-07
+    5.612039123698789e-08
+    1.041523408089798e-07
+    4.178942359865563e-07
+    3.400841842317408e-08
+    5.611990481856641e-08
+    1.625801463827058e-07
+     4.22577850503956e-07
+ 2.59e+10    
+    4.222135531657543e-07
+    1.626000371386579e-07
+    4.180188757731971e-07
+    5.616311751980579e-08
+    1.042078714354989e-07
+    4.179633099556654e-07
+    3.403646387877042e-08
+    5.616267614972115e-08
+    1.626494175474773e-07
+    4.226607773417315e-07
+ 2.6e+10     
+    4.222966142158299e-07
+    1.626693191553496e-07
+    4.180879799013521e-07
+    5.620572092897114e-08
+    1.042633935433789e-07
+    4.180324731885188e-07
+    3.406428938218306e-08
+     5.62053250490157e-08
+    1.627187449791744e-07
+    4.227438506535285e-07
+ 2.61e+10    
+    4.223798235019893e-07
+    1.627386577939612e-07
+    4.181571734432985e-07
+    5.624820179158967e-08
+    1.043189076793298e-07
+    4.181017265117842e-07
+    3.409189520493803e-08
+    5.624785184451268e-08
+    1.627881293570709e-07
+    4.228270712273272e-07
+ 2.62e+10    
+    4.224631817997395e-07
+    1.628080537216175e-07
+    4.182264572239925e-07
+    5.629056043078532e-08
+     1.04374414374715e-07
+    4.181710707416323e-07
+    3.411928162155219e-08
+     5.62902568602992e-08
+    1.628575713489219e-07
+    4.229104398440131e-07
+ 2.63e+10    
+    4.225466898772789e-07
+    1.628775075940736e-07
+    4.182958320585598e-07
+    5.633279716564166e-08
+     1.04429914145798e-07
+    4.182405066836725e-07
+    3.414644890937273e-08
+    5.633254041642737e-08
+     1.62927071611009e-07
+    4.229939572773261e-07
+ 2.64e+10    
+    4.226303484954613e-07
+     1.62947020055761e-07
+    4.183652987522126e-07
+    5.637491231114729e-08
+    1.044854074939885e-07
+    4.183100351328982e-07
+     3.41733973484209e-08
+    5.637470282885897e-08
+    1.629966307881905e-07
+    4.230776242938196e-07
+ 2.65e+10    
+    4.227141584077653e-07
+     1.63016591739838e-07
+     4.18434858100163e-07
+    5.641690617814422e-08
+     1.04540894906087e-07
+    4.183796568736315e-07
+    3.420012722123915e-08
+    5.641674440941284e-08
+    1.630662495139544e-07
+    4.231614416528216e-07
+ 2.66e+10    
+    4.227981203602653e-07
+    1.630862232682424e-07
+    4.185045108875447e-07
+    5.645877907327999e-08
+    1.045963768545277e-07
+    4.184493726794747e-07
+    3.422663881274228e-08
+     5.64586654657161e-08
+    1.631359284104754e-07
+    4.232454101063988e-07
+ 2.67e+10    
+    4.228822350916123e-07
+    1.631559152517494e-07
+    4.185742578893388e-07
+     5.65005312989626e-08
+    1.046518537976199e-07
+    4.185191833132644e-07
+    3.425293241007202e-08
+    5.650046630115845e-08
+    1.632056680886748e-07
+    4.233295303993305e-07
+ 2.68e+10    
+    4.229665033330111e-07
+    1.632256682900296e-07
+    4.186440998702984e-07
+    5.654216315331895e-08
+    1.047073261797885e-07
+     4.18589089527032e-07
+    3.427900830245528e-08
+      5.6542147214849e-08
+    1.632754691482834e-07
+    4.234138032690808e-07
+ 2.69e+10    
+    4.230509258082109e-07
+    1.632954829717123e-07
+    4.187140375848813e-07
+    5.658367493015569e-08
+    1.047627944318111e-07
+    4.186590920619657e-07
+    3.430486678106588e-08
+      5.6583708501577e-08
+    1.633453321779077e-07
+    4.234982294457772e-07
+ 2.7e+10     
+    4.231355032334901e-07
+    1.633653598744496e-07
+    4.187840717771828e-07
+     5.66250669189237e-08
+    1.048182589710547e-07
+    4.187291916483781e-07
+    3.433050813888977e-08
+    5.662515045177443e-08
+    1.634152577550982e-07
+    4.235828096521946e-07
+ 2.71e+10    
+    4.232202363176509e-07
+    1.634352995649845e-07
+     4.18854203180877e-07
+    5.666633940468455e-08
+    1.048737202017096e-07
+    4.187993890056792e-07
+    3.435593267059348e-08
+    5.666647335148232e-08
+    1.634852464464208e-07
+    4.236675446037422e-07
+ 2.72e+10    
+     4.23305125762018e-07
+    1.635053025992198e-07
+    4.189244325191561e-07
+    5.670749266808042e-08
+    1.049291785150214e-07
+    4.188696848423506e-07
+    3.438114067239605e-08
+    5.670767748231886e-08
+    1.635552988075298e-07
+    4.237524350084509e-07
+ 2.73e+10    
+    4.233901722604328e-07
+    1.635753695222905e-07
+    4.189947605046788e-07
+    5.674852698530597e-08
+    1.049846342895205e-07
+    4.189400798559254e-07
+    3.440613244194403e-08
+    5.674876312145079e-08
+    1.636254153832442e-07
+    4.238374815669694e-07
+ 2.74e+10    
+    4.234753764992631e-07
+    1.636455008686371e-07
+    4.190651878395186e-07
+    5.678944262808318e-08
+      1.0504008789125e-07
+    4.190105747329759e-07
+    3.443090827818984e-08
+    5.678973054156697e-08
+    1.636955967076252e-07
+    4.239226849725596e-07
+ 2.75e+10    
+    4.235607391574028e-07
+    1.637156971620819e-07
+    4.191357152151193e-07
+    5.683023986363835e-08
+    1.050955396739907e-07
+    4.190811701490968e-07
+    3.445546848127299e-08
+    5.683058001085425e-08
+    1.637658433040561e-07
+    4.240080459110964e-07
+ 2.76e+10    
+    4.236462609062833e-07
+     1.63785958915906e-07
+    4.192063433122512e-07
+    5.687091895468161e-08
+    1.051509899794837e-07
+    4.191518667689015e-07
+     3.44798133524047e-08
+    5.687131179297612e-08
+    1.638361556853231e-07
+    4.240935650610712e-07
+ 2.77e+10    
+    4.237319424098873e-07
+    1.638562866329288e-07
+    4.192770728009769e-07
+    5.691148015938862e-08
+    1.052064391376515e-07
+    4.192226652460178e-07
+    3.450394319375523e-08
+    5.691192614705319e-08
+    1.639065343536996e-07
+    4.241792430935967e-07
+ 2.78e+10    
+    4.238177843247581e-07
+    1.639266808055889e-07
+    4.193479043406154e-07
+    5.695192373138439e-08
+    1.052618874668152e-07
+    4.192935662230887e-07
+    3.452785830834425e-08
+    5.695242332764607e-08
+    1.639769798010304e-07
+    4.242650806724165e-07
+ 2.79e+10    
+    4.239037873000199e-07
+    1.639971419160256e-07
+    4.194188385797136e-07
+    5.699224991972951e-08
+    1.053173352739107e-07
+    4.193645703317782e-07
+    3.455155899993415e-08
+    5.699280358474041e-08
+    1.640474925088177e-07
+    4.243510784539147e-07
+ 2.8e+10     
+    4.239899519773951e-07
+    1.640676704361633e-07
+    4.194898761560229e-07
+    5.703245896890795e-08
+    1.053727828547015e-07
+    4.194356781927801e-07
+    3.457504557292607e-08
+    5.703306716373383e-08
+    1.641180729483095e-07
+    4.244372370871309e-07
+ 2.81e+10    
+    4.240762789912266e-07
+    1.641382668277958e-07
+    4.195610176964782e-07
+    5.707255111881729e-08
+    1.054282304939889e-07
+     4.19506890415831e-07
+    3.459831833225886e-08
+    5.707321430542502e-08
+    1.641887215805871e-07
+    4.245235572137751e-07
+ 2.82e+10    
+    4.241627689685003e-07
+    1.642089315426724e-07
+    4.196322638171825e-07
+    5.711252660476059e-08
+    1.054836784658202e-07
+    4.195782075997288e-07
+    3.462137758331063e-08
+    5.711324524600474e-08
+    1.642594388566562e-07
+    4.246100394682474e-07
+ 2.83e+10    
+    4.242494225288711e-07
+    1.642796650225849e-07
+    4.197036151233957e-07
+    5.715238565744032e-08
+    1.055391270336946e-07
+    4.196496303323538e-07
+    3.464422363180296e-08
+    5.715316021704826e-08
+    1.643302252175371e-07
+     4.24696684477656e-07
+ 2.84e+10    
+    4.243362402846895e-07
+    1.643504676994556e-07
+    4.197750722095296e-07
+    5.719212850295388e-08
+    1.055945764507655e-07
+    4.197211591906955e-07
+    3.466685678370793e-08
+    5.719295944551049e-08
+    1.644010810943569e-07
+    4.247834928618426e-07
+ 2.85e+10    
+    4.244232228410336e-07
+    1.644213399954261e-07
+    4.198466356591428e-07
+    5.723175536279065e-08
+    1.056500269600406e-07
+    4.197927947408799e-07
+    3.468927734515742e-08
+    5.723264315372195e-08
+    1.644720069084422e-07
+    4.248704652334038e-07
+ 2.86e+10    
+    4.245103707957358e-07
+    1.644922823229475e-07
+     4.19918306044948e-07
+    5.727126645383155e-08
+    1.057054787945808e-07
+    4.198645375382063e-07
+    3.471148562235523e-08
+    5.727221155938694e-08
+    1.645430030714127e-07
+    4.249576021977201e-07
+ 2.87e+10    
+     4.24597684739419e-07
+      1.6456329508487e-07
+    4.199900839288158e-07
+    5.731066198834909e-08
+    1.057609321776942e-07
+    4.199363881271829e-07
+    3.473348192149148e-08
+    5.731166487558321e-08
+    1.646140699852749e-07
+    4.250449043529828e-07
+ 2.88e+10    
+    4.246851652555296e-07
+    1.646343786745352e-07
+    4.200619698617887e-07
+    5.734994217400975e-08
+    1.058163873231294e-07
+      4.2000834704157e-07
+     3.47552665486595e-08
+    5.735100331076312e-08
+    1.646852080425174e-07
+    4.251323722902232e-07
+ 2.89e+10    
+    4.247728129203736e-07
+    1.647055334758672e-07
+     4.20133964384097e-07
+    5.738910721387759e-08
+    1.058718444352658e-07
+    4.200804148044239e-07
+    3.477683980977518e-08
+    5.739022706875657e-08
+    1.647564176262063e-07
+    4.252200065933459e-07
+ 2.9e+10     
+    4.248606283031526e-07
+     1.64776759863465e-07
+    4.202060680251811e-07
+    5.742815730641933e-08
+    1.059273037093007e-07
+    4.201525919281482e-07
+     3.47982020104984e-08
+    5.742933634877505e-08
+    1.648276991100802e-07
+    4.253078078391585e-07
+ 2.91e+10    
+    4.249486119660035e-07
+    1.648480582026954e-07
+    4.202782813037182e-07
+    5.746709264551099e-08
+    1.059827653314351e-07
+     4.20224878914546e-07
+    3.481935345615722e-08
+    5.746833134541764e-08
+    1.648990528586476e-07
+    4.253957765974113e-07
+ 2.92e+10    
+     4.25036764464039e-07
+    1.649194288497865e-07
+    4.203506047276503e-07
+    5.750591342044535e-08
+    1.060382294790553e-07
+    4.202972762548768e-07
+     3.48402944516738e-08
+    5.750721224867766e-08
+    1.649704792272822e-07
+    4.254839134308269e-07
+ 2.93e+10    
+    4.251250863453866e-07
+    1.649908721519209e-07
+    4.204230387942241e-07
+    5.754461981594148e-08
+    1.060936963209143e-07
+     4.20369784429917e-07
+    3.486102530149282e-08
+    5.754597924395147e-08
+    1.650419785623205e-07
+    4.255722188951413e-07
+ 2.94e+10    
+    4.252135781512317e-07
+    1.650623884473305e-07
+    4.204955839900273e-07
+    5.758321201215504e-08
+    1.061491660173086e-07
+    4.204424039100259e-07
+    3.488154630951213e-08
+    5.758463251204793e-08
+    1.651135512011584e-07
+    4.256606935391408e-07
+ 2.95e+10    
+    4.253022404158606e-07
+    1.651339780653893e-07
+    4.205682407910346e-07
+    5.762169018468981e-08
+    1.062046387202533e-07
+      4.2051513515521e-07
+     3.49018577790153e-08
+    5.762317222919949e-08
+    1.651851974723488e-07
+    4.257493379047024e-07
+ 2.96e+10    
+    4.253910736667052e-07
+    1.652056413267092e-07
+    4.206410096626566e-07
+    5.766005450461055e-08
+    1.062601145736559e-07
+    4.205879786151982e-07
+    3.492196001260637e-08
+    5.766159856707419e-08
+    1.652569176956983e-07
+    4.258381525268323e-07
+ 2.97e+10    
+     4.25480078424386e-07
+    1.652773785432342e-07
+    4.207138910597957e-07
+    5.769830513845688e-08
+    1.063155937134854e-07
+    4.206609347295131e-07
+    3.494185331214672e-08
+    5.769991169278927e-08
+    1.653287121823646e-07
+    4.259271379337101e-07
+ 2.98e+10    
+    4.255692552027613e-07
+    1.653491900183349e-07
+    4.207868854268993e-07
+    5.773644224825845e-08
+    1.063710762679412e-07
+    4.207340039275511e-07
+    3.496153797869384e-08
+    5.773811176892537e-08
+    1.654005812349541e-07
+    4.260162946467288e-07
+ 2.99e+10    
+    4.256586045089695e-07
+    1.654210760469031e-07
+    4.208599931980261e-07
+    5.777446599155064e-08
+    1.064265623576184e-07
+    4.208071866286617e-07
+    3.498101431244202e-08
+    5.777619895354211e-08
+    1.654725251476192e-07
+    4.261056231805403e-07
+ 3e+10       
+    4.257481268434799e-07
+    1.654930369154476e-07
+    4.209332147969124e-07
+    5.781237652139211e-08
+    1.064820520956712e-07
+    4.208804832422342e-07
+    3.500028261266523e-08
+    5.781417340019499e-08
+    1.655445442061549e-07
+    4.261951240430981e-07
+ 3.01e+10    
+    4.258378227001411e-07
+    1.655650729021879e-07
+    4.210065506370407e-07
+    5.785017398638242e-08
+    1.065375455879734e-07
+    4.209538941677823e-07
+     3.50193431776616e-08
+    5.785203525795258e-08
+    1.656166386880961e-07
+    4.262847977357036e-07
+ 3.02e+10    
+    4.259276925662262e-07
+    1.656371842771496e-07
+    4.210800011217164e-07
+    5.788785853068122e-08
+    1.065930429332777e-07
+    4.210274197950362e-07
+    3.503819630469995e-08
+    5.788978467141544e-08
+    1.656888088628146e-07
+    4.263746447530506e-07
+ 3.03e+10    
+    4.260177369224856e-07
+    1.657093713022592e-07
+    4.211535666441472e-07
+     5.79254302940282e-08
+    1.066485442233718e-07
+    4.211010605040349e-07
+    3.505684228996802e-08
+    5.792742178073552e-08
+    1.657610549916155e-07
+    4.264646655832732e-07
+ 3.04e+10    
+    4.261079562431952e-07
+    1.657816342314376e-07
+    4.212272475875223e-07
+     5.79628894117636e-08
+    1.067040495432322e-07
+    4.211748166652223e-07
+    3.507528142852267e-08
+    5.796494672163671e-08
+    1.658333773278337e-07
+    4.265548607079922e-07
+ 3.05e+10    
+    4.261983509962067e-07
+    1.658539733106959e-07
+    4.213010443251047e-07
+    5.800023601485009e-08
+    1.067595589711765e-07
+    4.212486886395456e-07
+    3.509351401424157e-08
+    5.800235962543599e-08
+    1.659057761169291e-07
+    4.266452306023621e-07
+ 3.06e+10    
+    4.262889216430001e-07
+    1.659263887782289e-07
+    4.213749572203164e-07
+    5.803747022989494e-08
+    1.068150725790129e-07
+    4.213226767785565e-07
+    3.511154033977706e-08
+    5.803966061906595e-08
+     1.65978251596584e-07
+    4.267357757351223e-07
+ 3.07e+10    
+    4.263796686387331e-07
+    1.659988808645086e-07
+    4.214489866268353e-07
+    5.807459217917325e-08
+    1.068705904321877e-07
+    4.213967814245148e-07
+    3.512936069651106e-08
+    5.807684982509752e-08
+    1.660508039967967e-07
+    4.268264965686412e-07
+ 3.08e+10    
+     4.26470592432292e-07
+    1.660714497923787e-07
+    4.215231328886917e-07
+    5.811160198065191e-08
+    1.069261125899303e-07
+    4.214710029104931e-07
+    3.514697537451227e-08
+    5.811392736176371e-08
+    1.661234335399774e-07
+    4.269173935589699e-07
+ 3.09e+10    
+    4.265616934663481e-07
+    1.661440957771474e-07
+    4.215973963403684e-07
+    5.814849974801419e-08
+     1.06981639105397e-07
+    4.215453415604877e-07
+     3.51643846624947e-08
+     5.81508933429844e-08
+    1.661961404410425e-07
+    4.270084671558901e-07
+ 3.1e+10     
+    4.266529721774035e-07
+    1.662168190266808e-07
+    4.216717773069063e-07
+    5.818528559068501e-08
+    1.070371700258114e-07
+    4.216197976895254e-07
+    3.518158884777771e-08
+     5.81877478783913e-08
+    1.662689249075082e-07
+     4.27099717802963e-07
+ 3.11e+10    
+    4.267444289958495e-07
+    1.662896197414951e-07
+    4.217462761040097e-07
+    5.822195961385695e-08
+    1.070927053926035e-07
+    4.216943716037776e-07
+    3.519858821624792e-08
+    5.822449107335421e-08
+    1.663417871395852e-07
+    4.271911459375829e-07
+ 3.12e+10    
+    4.268360643460152e-07
+     1.66362498114849e-07
+    4.218208930381568e-07
+    5.825852191851663e-08
+    1.071482452415468e-07
+    4.217690636006735e-07
+    3.521538305232235e-08
+    5.826112302900736e-08
+      1.6641472733027e-07
+    4.272827519910243e-07
+ 3.13e+10    
+    4.269278786462235e-07
+    1.664354543328361e-07
+    4.218956284067135e-07
+    5.829497260147232e-08
+    1.072037896028925e-07
+    4.218438739690179e-07
+    3.523197363891331e-08
+    5.829764384227682e-08
+    1.664877456654388e-07
+    4.273745363884961e-07
+ 3.14e+10    
+    4.270198723088414e-07
+    1.665084885744753e-07
+    4.219704824980479e-07
+    5.833131175538119e-08
+     1.07259338501503e-07
+    4.219188029891062e-07
+    3.524836025739467e-08
+    5.833405360590832e-08
+    1.665608423239389e-07
+     4.27466499549191e-07
+ 3.15e+10    
+    4.271120457403366e-07
+    1.665816010118031e-07
+     4.22045455591649e-07
+    5.836753946877799e-08
+    1.073148919569818e-07
+    4.219938509328447e-07
+    3.526454318756953e-08
+    5.837035240849569e-08
+    1.666340174776799e-07
+    4.275586418863371e-07
+ 3.16e+10    
+     4.27204399341327e-07
+    1.666547918099626e-07
+    4.221205479582467e-07
+     5.84036558261037e-08
+    1.073704499838029e-07
+    4.220690180638714e-07
+     3.52805227076395e-08
+    5.840654033450997e-08
+    1.667072712917249e-07
+    4.276509638072515e-07
+ 3.17e+10    
+    4.272969335066379e-07
+     1.66728061127294e-07
+    4.221957598599349e-07
+    5.843966090773492e-08
+    1.074260125914371e-07
+    4.221443046376777e-07
+    3.529629909417519e-08
+    5.844261746432883e-08
+    1.667806039243797e-07
+    4.277434657133902e-07
+ 3.18e+10    
+    4.273896486253528e-07
+    1.668014091154245e-07
+    4.222710915502972e-07
+    5.847555479001358e-08
+    1.074815797844767e-07
+    4.222197109017305e-07
+    3.531187262208819e-08
+    5.847858387426676e-08
+     1.66854015527283e-07
+    4.278361480004004e-07
+ 3.19e+10    
+     4.27482545080869e-07
+    1.668748359193559e-07
+    4.223465432745314e-07
+    5.851133754527745e-08
+    1.075371515627589e-07
+    4.222952370955981e-07
+    3.532724356460437e-08
+    5.851443963660549e-08
+     1.66927506245495e-07
+    4.279290110581739e-07
+ 3.2e+10     
+    4.275756232509492e-07
+    1.669483416775539e-07
+    4.224221152695806e-07
+    5.854700924189047e-08
+    1.075927279214858e-07
+     4.22370883451074e-07
+    3.534241219323853e-08
+    5.855018481962512e-08
+    1.670010762175852e-07
+    4.280220552708987e-07
+ 3.21e+10    
+    4.276688835077766e-07
+    1.670219265220349e-07
+    4.224978077642631e-07
+    5.858256994427413e-08
+    1.076483088513443e-07
+    4.224466501923029e-07
+    3.535737877777024e-08
+    5.858581948763538e-08
+    1.670747255757194e-07
+    4.281152810171097e-07
+ 3.22e+10    
+    4.277623262180081e-07
+    1.670955905784536e-07
+    4.225736209794036e-07
+    5.861801971293901e-08
+    1.077038943386229e-07
+      4.2252253753591e-07
+    3.537214358622126e-08
+    5.862134370100795e-08
+    1.671484544457475e-07
+    4.282086886697442e-07
+ 3.23e+10    
+    4.278559517428281e-07
+    1.671693339661888e-07
+     4.22649555127967e-07
+    5.865335860451636e-08
+    1.077594843653263e-07
+    4.225985456911235e-07
+    3.538670688483373e-08
+    5.865675751620821e-08
+    1.672222629472879e-07
+    4.283022785961922e-07
+ 3.24e+10    
+    4.279497604380006e-07
+    1.672431567984288e-07
+    4.227256104151928e-07
+     5.86885866717906e-08
+    1.078150789092897e-07
+    4.226746748599076e-07
+    3.540106893805007e-08
+    5.869206098582815e-08
+    1.672961511938137e-07
+    4.283960511583482e-07
+ 3.25e+10    
+    4.280437526539248e-07
+    1.673170591822572e-07
+    4.228017870387309e-07
+    5.872370396373179e-08
+      1.0787067794429e-07
+    4.227509252370894e-07
+    3.541523000849383e-08
+    5.872725415861945e-08
+    1.673701192927366e-07
+    4.284900067126663e-07
+ 3.26e+10    
+    4.281379287356854e-07
+    1.673910412187362e-07
+    4.228780851887793e-07
+    5.875871052552839e-08
+    1.079262814401555e-07
+    4.228272970104848e-07
+    3.542919035695167e-08
+    5.876233707952668e-08
+      1.6744416734549e-07
+    4.285841456102089e-07
+ 3.27e+10    
+    4.282322890231084e-07
+    1.674651030029906e-07
+    4.229545050482196e-07
+    5.879360639862062e-08
+    1.079818893628738e-07
+    4.229037903610323e-07
+    3.544295024235682e-08
+    5.879730978972109e-08
+    1.675182954476129e-07
+    4.286784681967024e-07
+ 3.28e+10    
+    4.283268338508127e-07
+    1.675392446242901e-07
+     4.23031046792756e-07
+    5.882839162073369e-08
+    1.080375016746981e-07
+    4.229804054629192e-07
+    3.545650992177321e-08
+     5.88321723266344e-08
+    1.675925036888307e-07
+    4.287729748125867e-07
+ 3.29e+10    
+    4.284215635482645e-07
+    1.676134661661325e-07
+    4.231077105910556e-07
+    5.886306622591178e-08
+    1.080931183342516e-07
+    4.230571424837105e-07
+    3.546986965038128e-08
+    5.886692472399329e-08
+    1.676667921531368e-07
+    4.288676657930689e-07
+ 3.3e+10     
+    4.285164784398273e-07
+     1.67687767706323e-07
+    4.231844966048848e-07
+    5.889763024455172e-08
+    1.081487392966301e-07
+    4.231340015844799e-07
+    3.548302968146429e-08
+    5.890156701185369e-08
+    1.677411609188729e-07
+    4.289625414681747e-07
+ 3.31e+10    
+    4.286115788448162e-07
+     1.67762149317056e-07
+    4.232614049892509e-07
+    5.893208370343734e-08
+    1.082043645135029e-07
+    4.232109829199374e-07
+    3.549599026639624e-08
+    5.893609921663574e-08
+    1.678156100588083e-07
+    4.290576021628006e-07
+ 3.32e+10    
+    4.287068650775509e-07
+    1.678366110649947e-07
+    4.233384358925412e-07
+    5.896642662577385e-08
+    1.082599939332122e-07
+    4.232880866385583e-07
+    3.550875165463048e-08
+    5.897052136115862e-08
+    1.678901396402188e-07
+     4.29152848196765e-07
+ 3.33e+10    
+    4.288023374474055e-07
+    1.679111530113491e-07
+    4.234155894566612e-07
+    5.900065903122234e-08
+    1.083156275008703e-07
+    4.233653128827114e-07
+    3.552131409368956e-08
+     5.90048334646758e-08
+    1.679647497249642e-07
+    4.292482798848604e-07
+ 3.34e+10    
+    4.288979962588627e-07
+    1.679857752119555e-07
+    4.234928658171771e-07
+    5.903478093593481e-08
+    1.083712651584561e-07
+     4.23442661788788e-07
+    3.553367782915609e-08
+    5.903903554291058e-08
+    1.680394403695653e-07
+    4.293438975369047e-07
+ 3.35e+10    
+    4.289938418115636e-07
+    1.680604777173516e-07
+    4.235702651034515e-07
+    5.906879235258875e-08
+    1.084269068449083e-07
+    4.235201334873275e-07
+    3.554584310466433e-08
+    5.907312760809142e-08
+    1.681142116252796e-07
+     4.29439701457792e-07
+ 3.36e+10    
+    4.290898744003607e-07
+    1.681352605728549e-07
+    4.236477874387852e-07
+    5.910269329042271e-08
+    1.084825524962189e-07
+    4.235977281031461e-07
+    3.555781016189326e-08
+    5.910710966898791e-08
+    1.681890635381769e-07
+    4.295356919475439e-07
+ 3.37e+10    
+    4.291860943153688e-07
+    1.682101238186372e-07
+    4.237254329405545e-07
+    5.913648375527125e-08
+    1.085382020455237e-07
+    4.236754457554611e-07
+    3.556957924056016e-08
+    5.914098173094655e-08
+    1.682639961492137e-07
+    4.296318693013609e-07
+ 3.38e+10    
+    4.292825018420141e-07
+     1.68285067489799e-07
+    4.238032017203497e-07
+    5.917016374960034e-08
+    1.085938554231915e-07
+    4.237532865580185e-07
+    3.558115057841531e-08
+    5.917474379592691e-08
+    1.683390094943061e-07
+    4.297282338096732e-07
+ 3.39e+10    
+    4.293790972610871e-07
+    1.683600916164443e-07
+    4.238810938841114e-07
+    5.920373327254312e-08
+    1.086495125569119e-07
+    4.238312506192148e-07
+    3.559252441123767e-08
+    5.920839586253771e-08
+    1.684141036044022e-07
+    4.298247857581882e-07
+ 3.4e+10     
+    4.294758808487921e-07
+    1.684351962237525e-07
+    4.239591095322688e-07
+    5.923719231993537e-08
+    1.087051733717819e-07
+    4.239093380422242e-07
+    3.560370097283145e-08
+    5.924193792607326e-08
+    1.684892785055547e-07
+    4.299215254279458e-07
+ 3.41e+10    
+    4.295728528767978e-07
+    1.685103813320513e-07
+    4.240372487598734e-07
+    5.927054088435122e-08
+    1.087608377903898e-07
+    4.239875489251176e-07
+    3.561468049502344e-08
+     5.92753699785496e-08
+    1.685645342189908e-07
+    4.300184530953643e-07
+ 3.42e+10    
+    4.296700136122853e-07
+    1.685856469568871e-07
+     4.24115511656735e-07
+    5.930377895513906e-08
+    1.088165057328983e-07
+    4.240658833609864e-07
+    3.562546320766133e-08
+     5.93086920087411e-08
+    1.686398707611818e-07
+    4.301155690322908e-07
+ 3.43e+10    
+    4.297673633180006e-07
+    1.686609931090959e-07
+    4.241938983075549e-07
+     5.93369065184573e-08
+    1.088721771171268e-07
+    4.241443414380636e-07
+    3.563604933861296e-08
+    5.934190400221724e-08
+    1.687152881439133e-07
+    4.302128735060527e-07
+ 3.44e+10    
+    4.298649022523017e-07
+    1.687364197948729e-07
+    4.242724087920601e-07
+     5.93699235573107e-08
+    1.089278518586304e-07
+    4.242229232398422e-07
+     3.56464391137663e-08
+    5.937500594137894e-08
+    1.687907863743521e-07
+    4.303103667795046e-07
+ 3.45e+10    
+    4.299626306692078e-07
+    1.688119270158399e-07
+    4.243510431851307e-07
+    5.940283005158578e-08
+    1.089835298707788e-07
+    4.243016288451924e-07
+    3.565663275703017e-08
+    5.940799780549527e-08
+    1.688663654551136e-07
+    4.304080491110788e-07
+ 3.46e+10    
+    4.300605488184482e-07
+    1.688875147691143e-07
+    4.244298015569347e-07
+    5.943562597808752e-08
+    1.090392110648337e-07
+    4.243804583284812e-07
+    3.566663049033612e-08
+    5.944087957074046e-08
+    1.689420253843289e-07
+    4.305059207548332e-07
+ 3.47e+10    
+    4.301586569455114e-07
+    1.689631830473751e-07
+    4.245086839730534e-07
+    5.946831131057509e-08
+    1.090948953500239e-07
+    4.244594117596861e-07
+    3.567643253364063e-08
+    5.947365121023028e-08
+    1.690177661557087e-07
+    4.306039819604994e-07
+ 3.48e+10    
+    4.302569552916909e-07
+    1.690389318389287e-07
+    4.245876904946092e-07
+    5.950088601979817e-08
+    1.091505826336192e-07
+    4.245384892045102e-07
+    3.568603910492854e-08
+    5.950631269405914e-08
+    1.690935877586093e-07
+    4.307022329735318e-07
+ 3.49e+10    
+    4.303554440941358e-07
+    1.691147611277743e-07
+    4.246668211783929e-07
+    5.953335007353302e-08
+    1.092062728210041e-07
+    4.246176907244952e-07
+    3.569545042021691e-08
+    5.953886398933674e-08
+    1.691694901780955e-07
+    4.308006740351543e-07
+ 3.5e+10     
+    4.304541235858954e-07
+    1.691906708936673e-07
+    4.247460760769855e-07
+     5.95657034366187e-08
+    1.092619658157478e-07
+    4.246970163771321e-07
+    3.570466669355988e-08
+    5.957130506022495e-08
+    1.692454733950033e-07
+    4.308993053824099e-07
+ 3.51e+10    
+    4.305529939959679e-07
+    1.692666611121831e-07
+     4.24825455238883e-07
+    5.959794607099331e-08
+    1.093176615196751e-07
+    4.247764662159721e-07
+    3.571368813705406e-08
+    5.960363586797463e-08
+     1.69321537386002e-07
+    4.309981272482048e-07
+ 3.52e+10    
+    4.306520555493467e-07
+    1.693427317547793e-07
+     4.24904958708616e-07
+    5.963007793573021e-08
+    1.093733598329344e-07
+    4.248560402907352e-07
+    3.572251496084483e-08
+    5.963585637096239e-08
+    1.693976821236549e-07
+    4.310971398613575e-07
+ 3.53e+10    
+    4.307513084670664e-07
+    1.694188827888566e-07
+    4.249845865268688e-07
+      5.9662098987074e-08
+     1.09429060654065e-07
+    4.249357386474159e-07
+    3.573114737313324e-08
+    5.966796652472749e-08
+    1.694739075764799e-07
+    4.311963434466458e-07
+ 3.54e+10    
+    4.308507529662486e-07
+    1.694951141778196e-07
+     4.25064338730597e-07
+    5.969400917847693e-08
+     1.09484763880063e-07
+    4.250155613283901e-07
+    3.573958558018362e-08
+    5.969996628200855e-08
+     1.69550213709008e-07
+    4.312957382248509e-07
+ 3.55e+10    
+    4.309503892601484e-07
+    1.695714258811365e-07
+    4.251442153531431e-07
+    5.972580846063501e-08
+    1.095404694064458e-07
+    4.250955083725181e-07
+    3.574782978633188e-08
+    5.973185559278028e-08
+    1.696266004818424e-07
+    4.313953244128052e-07
+ 3.56e+10    
+    4.310502175581994e-07
+    1.696478178543975e-07
+    4.252242164243507e-07
+    5.975749678152405e-08
+    1.095961771273149e-07
+    4.251755798152467e-07
+    3.575588019399455e-08
+    5.976363440429019e-08
+    1.697030678517153e-07
+    4.314951022234381e-07
+ 3.57e+10    
+    4.311502380660575e-07
+     1.69724290049373e-07
+     4.25304341970675e-07
+    5.978907408643571e-08
+    1.096518869354184e-07
+    4.252557756887095e-07
+    3.576373700367835e-08
+    5.979530266109541e-08
+    1.697796157715454e-07
+    4.315950718658202e-07
+ 3.58e+10    
+    4.312504509856482e-07
+    1.698008424140703e-07
+    4.253845920152935e-07
+     5.98205403180139e-08
+    1.097075987222111e-07
+    4.253360960218272e-07
+    3.577140041399055e-08
+    5.982686030509898e-08
+     1.69856244190493e-07
+    4.316952335452083e-07
+ 3.59e+10    
+    4.313508565152069e-07
+    1.698774748927897e-07
+    4.254649665782147e-07
+    5.985189541629034e-08
+    1.097633123779143e-07
+    4.254165408404027e-07
+    3.577887062164978e-08
+    5.985830727558681e-08
+    1.699329530540151e-07
+    4.317955874630918e-07
+ 3.6e+10     
+     4.31451454849327e-07
+    1.699541874261798e-07
+     4.25545465676382e-07
+    5.988313931872086e-08
+    1.098190277915737e-07
+    4.254971101672169e-07
+    3.578614782149773e-08
+    5.988964350926393e-08
+    1.700097423039194e-07
+    4.318961338172351e-07
+ 3.61e+10    
+    4.315522461789999e-07
+    1.700309799512917e-07
+    4.256260893237793e-07
+     5.99142719602212e-08
+    1.098747448511162e-07
+    4.255778040221252e-07
+    3.579323220651114e-08
+    5.992086894029097e-08
+    1.700866118784185e-07
+    4.319968728017228e-07
+ 3.62e+10    
+    4.316532306916612e-07
+    1.701078524016328e-07
+    4.257068375315323e-07
+    5.994529327320287e-08
+    1.099304634434059e-07
+    4.256586224221449e-07
+    3.580012396781464e-08
+    5.995198350032056e-08
+    1.701635617121807e-07
+    4.320978046070027e-07
+ 3.63e+10    
+    4.317544085712318e-07
+     1.70184804707219e-07
+     4.25787710308009e-07
+      5.9976203187609e-08
+    1.099861834542985e-07
+    4.257395653815492e-07
+    3.580682329469412e-08
+    5.998298711853368e-08
+    1.702405917363833e-07
+    4.321989294199299e-07
+ 3.64e+10    
+    4.318557799981594e-07
+    1.702618367946269e-07
+    4.258687076589166e-07
+    6.000700163095004e-08
+    1.100419047686946e-07
+    4.258206329119541e-07
+    3.581333037461054e-08
+    6.001387972167579e-08
+    1.703177018787624e-07
+    4.323002474238094e-07
+ 3.65e+10    
+    4.319573451494638e-07
+    1.703389485870448e-07
+    4.259498295873981e-07
+    6.003768852833947e-08
+     1.10097627270592e-07
+     4.25901825022406e-07
+    3.581964539321447e-08
+    6.004466123409299e-08
+    1.703948920636633e-07
+    4.324017587984389e-07
+ 3.66e+10    
+     4.32059104198775e-07
+    1.704161400043221e-07
+    4.260310760941252e-07
+     6.00682638025293e-08
+    1.101533508431367e-07
+    4.259831417194648e-07
+    3.582576853436109e-08
+    6.007533157776812e-08
+    1.704721622120895e-07
+    4.325034637201506e-07
+ 3.67e+10    
+    4.321610573163779e-07
+    1.704934109630197e-07
+    4.261124471773919e-07
+    6.009872737394578e-08
+    1.102090753686729e-07
+    4.260645830072903e-07
+    3.583169998012585e-08
+    6.010589067235671e-08
+    1.705495122417516e-07
+    4.326053623618552e-07
+ 3.68e+10    
+     4.32263204669251e-07
+    1.705707613764576e-07
+    4.261939428332005e-07
+    6.012907916072456e-08
+    1.102648007287918e-07
+    4.261461488877209e-07
+    3.583743991082039e-08
+     6.01363384352226e-08
+    1.706269420671143e-07
+    4.327074548930798e-07
+ 3.69e+10    
+    4.323655464211087e-07
+    1.706481911547631e-07
+     4.26275563055354e-07
+    6.015931907874644e-08
+    1.103205268043797e-07
+    4.262278393603556e-07
+    3.584298850500937e-08
+    6.016667478147429e-08
+     1.70704451599444e-07
+    4.328097414800135e-07
+ 3.7e+10     
+    4.324680827324404e-07
+    1.707257002049176e-07
+    4.263573078355378e-07
+    6.018944704167225e-08
+    1.103762534756643e-07
+     4.26309654422631e-07
+    3.584834593952746e-08
+    6.019689962399991e-08
+    1.707820407468543e-07
+    4.329122222855463e-07
+ 3.71e+10    
+    4.325708137605515e-07
+    1.708032884308022e-07
+    4.264391771634041e-07
+    6.021946296097824e-08
+    1.104319806222605e-07
+    4.263915940698967e-07
+    3.585351238949702e-08
+    6.022701287350329e-08
+    1.708597094143518e-07
+    4.330148974693087e-07
+ 3.72e+10    
+    4.326737396596023e-07
+    1.708809557332441e-07
+     4.26521171026655e-07
+    6.024936674599118e-08
+    1.104877081232152e-07
+    4.264736582954913e-07
+    3.585848802834627e-08
+    6.025701443853919e-08
+    1.709374575038804e-07
+    4.331177671877144e-07
+ 3.73e+10    
+    4.327768605806472e-07
+    1.709587020100599e-07
+    4.266032894111198e-07
+    6.027915830392331e-08
+     1.10543435857051e-07
+    4.265558470908168e-07
+     3.58632730278278e-08
+    6.028690422554879e-08
+    1.710152849143655e-07
+    4.332208315939989e-07
+ 3.74e+10    
+    4.328801766716759e-07
+    1.710365271561004e-07
+     4.26685532300833e-07
+    6.030883753990728e-08
+    1.105991637018084e-07
+    4.266381604454062e-07
+    3.586786755803778e-08
+    6.031668213889475e-08
+    1.710931915417573e-07
+    4.333240908382597e-07
+ 3.75e+10    
+     4.32983688077648e-07
+     1.71114431063293e-07
+     4.26767899678111e-07
+    6.033840435703093e-08
+     1.10654891535088e-07
+    4.267205983469954e-07
+    3.587227178743533e-08
+    6.034634808089645e-08
+    1.711711772790719e-07
+    4.334275450674931e-07
+ 3.76e+10    
+     4.33087394940534e-07
+    1.711924136206842e-07
+    4.268503915236235e-07
+    6.036785865637196e-08
+    1.107106192340908e-07
+    4.268031607815906e-07
+    3.587648588286272e-08
+    6.037590195186514e-08
+    1.712492420164355e-07
+    4.335311944256392e-07
+ 3.77e+10    
+    4.331912973993536e-07
+    1.712704747144812e-07
+    4.269330078164663e-07
+    6.039720033703275e-08
+    1.107663466756583e-07
+    4.268858477335346e-07
+    3.588051000956563e-08
+    6.040534365013853e-08
+    1.713273856411229e-07
+    4.336350390536138e-07
+ 3.78e+10    
+     4.33295395590211e-07
+    1.713486142280924e-07
+    4.270157485342306e-07
+    6.042642929617449e-08
+     1.10822073736311e-07
+    4.269686591855714e-07
+    3.588434433121408e-08
+    6.043467307211582e-08
+    1.714056080375994e-07
+    4.337390790893498e-07
+ 3.79e+10    
+    4.333996896463341e-07
+    1.714268320421682e-07
+    4.270986136530707e-07
+    6.045554542905199e-08
+    1.108778002922868e-07
+    4.270515951189084e-07
+     3.58879890099238e-08
+    6.046389011229236e-08
+    1.714839090875599e-07
+    4.338433146678366e-07
+ 3.8e+10     
+    4.335041796981111e-07
+    1.715051280346399e-07
+    4.271816031477678e-07
+    6.048454862904772e-08
+    1.109335262195775e-07
+    4.271346555132795e-07
+    3.589144420627781e-08
+    6.049299466329391e-08
+    1.715622886699679e-07
+    4.339477459211541e-07
+ 3.81e+10    
+    4.336088658731252e-07
+    1.715835020807581e-07
+     4.27264716991798e-07
+    6.051343878770596e-08
+    1.109892513939654e-07
+    4.272178403470022e-07
+    3.589471007934869e-08
+    6.052198661591158e-08
+    1.716407466610942e-07
+    4.340523729785137e-07
+ 3.82e+10    
+     4.33713748296193e-07
+    1.716619540531313e-07
+    4.273479551573898e-07
+    6.054221579476704e-08
+    1.110449756910582e-07
+    4.273011495970391e-07
+    3.589778678672085e-08
+    6.055086585913552e-08
+    1.717192829345536e-07
+    4.341571959662911e-07
+ 3.83e+10    
+    4.338188270893996e-07
+    1.717404838217633e-07
+    4.274313176155865e-07
+    6.057087953820138e-08
+    1.111006989863241e-07
+    4.273845832390511e-07
+    3.590067448451384e-08
+    6.057963228018962e-08
+    1.717978973613432e-07
+    4.342622150080674e-07
+ 3.84e+10    
+    4.339241023721331e-07
+    1.718190912540893e-07
+    4.275148043363045e-07
+    6.059942990424298e-08
+    1.111564211551245e-07
+    4.274681412474552e-07
+     3.59033733274053e-08
+    6.060828576456523e-08
+    1.718765898098778e-07
+    4.343674302246629e-07
+ 3.85e+10    
+    4.340295742611213e-07
+    1.718977762150124e-07
+    4.275984152883903e-07
+    6.062786677742343e-08
+     1.11212142072748e-07
+    4.275518235954764e-07
+    3.590588346865471e-08
+     6.06368261960553e-08
+    1.719553601460263e-07
+    4.344728417341727e-07
+ 3.86e+10    
+    4.341352428704664e-07
+    1.719765385669389e-07
+    4.276821504396723e-07
+    6.065619004060562e-08
+    1.112678616144412e-07
+     4.27635630255201e-07
+    3.590820506012756e-08
+     6.06652534567879e-08
+    1.720342082331458e-07
+    4.345784496520029e-07
+ 3.87e+10    
+    4.342411083116776e-07
+    1.720553781698126e-07
+    4.277660097570174e-07
+    6.068439957501697e-08
+    1.113235796554407e-07
+    4.277195611976258e-07
+    3.591033825231954e-08
+    6.069356742726021e-08
+    1.721131339321177e-07
+    4.346842540909069e-07
+ 3.88e+10    
+     4.34347170693708e-07
+    1.721342948811496e-07
+    4.278499932063817e-07
+    6.071249526028309e-08
+    1.113792960710036e-07
+    4.278036163927097e-07
+    3.591228319438151e-08
+    6.072176798637194e-08
+    1.721921371013805e-07
+    4.347902551610192e-07
+ 3.89e+10    
+    4.344534301229859e-07
+    1.722132885560719e-07
+    4.279341007528592e-07
+    6.074047697446092e-08
+     1.11435010736437e-07
+    4.278877958094186e-07
+    3.591404003414441e-08
+    6.074985501145868e-08
+    1.722712175969633e-07
+      4.3489645296989e-07
+ 3.9e+10     
+    4.345598867034505e-07
+    1.722923590473391e-07
+      4.2801833236073e-07
+    6.076834459407194e-08
+     1.11490723527127e-07
+    4.279720994157746e-07
+    3.591560891814475e-08
+    6.077782837832523e-08
+    1.723503752725189e-07
+    4.350028476225196e-07
+ 3.91e+10    
+    4.346665405365833e-07
+    1.723715062053818e-07
+    4.281026879935074e-07
+    6.079609799413513e-08
+    1.115464343185671e-07
+    4.280565271788982e-07
+    3.591698999165033e-08
+     6.08056879612788e-08
+    1.724296099793557e-07
+    4.351094392213928e-07
+ 3.92e+10    
+    4.347733917214426e-07
+    1.724507298783335e-07
+    4.281871676139831e-07
+    6.082373704820009e-08
+    1.116021429863856e-07
+    4.281410790650546e-07
+    3.591818339868642e-08
+    6.083343363316206e-08
+    1.725089215664696e-07
+    4.352162278665138e-07
+ 3.93e+10    
+    4.348804403546932e-07
+    1.725300299120609e-07
+    4.282717711842712e-07
+    6.085126162837969e-08
+     1.11657849406373e-07
+    4.282257550396953e-07
+    3.591918928206199e-08
+    6.086106526538595e-08
+    1.725883098805749e-07
+    4.353232136554356e-07
+ 3.94e+10    
+    4.349876865306433e-07
+    1.726094061501948e-07
+     4.28356498665847e-07
+     6.08786716053828e-08
+    1.117135534545074e-07
+    4.283105550674973e-07
+    3.592000778339654e-08
+    6.088858272796251e-08
+    1.726677747661348e-07
+    4.354303966832974e-07
+ 3.95e+10    
+    4.350951303412721e-07
+    1.726888584341605e-07
+    4.284413500195916e-07
+    6.090596684854692e-08
+    1.117692550069807e-07
+    4.283954791124069e-07
+    3.592063904314697e-08
+    6.091598588953752e-08
+    1.727473160653918e-07
+    4.355377770428551e-07
+ 3.96e+10    
+    4.352027718762629e-07
+     1.72768386603207e-07
+    4.285263252058286e-07
+    6.093314722587052e-08
+    1.118249539402235e-07
+    4.284805271376738e-07
+    3.592108320063501e-08
+    6.094327461742307e-08
+    1.728269336183967e-07
+    4.356453548245139e-07
+ 3.97e+10    
+    4.353106112230351e-07
+    1.728479904944357e-07
+    4.286114241843626e-07
+    6.096021260404554e-08
+    1.118806501309291e-07
+    4.285656991058923e-07
+    3.592134039407462e-08
+    6.097044877762987e-08
+     1.72906627263038e-07
+    4.357531301163606e-07
+ 3.98e+10    
+    4.354186484667749e-07
+    1.729276699428297e-07
+    4.286966469145147e-07
+    6.098716284848945e-08
+    1.119363434560771e-07
+    4.286509949790347e-07
+    3.592141076059998e-08
+     6.09975082348995e-08
+      1.7298639683507e-07
+    4.358611030041961e-07
+ 3.99e+10    
+    4.355268836904648e-07
+    1.730074247812808e-07
+    4.287819933551593e-07
+    6.101399782337748e-08
+    1.119920337929569e-07
+    4.287364147184887e-07
+    3.592129443629354e-08
+    6.102445285273668e-08
+    1.730662421681413e-07
+    4.359692735715649e-07
+ 4e+10       
+    4.356353169749146e-07
+     1.73087254840617e-07
+    4.288674634647542e-07
+    6.104071739167439e-08
+    1.120477210191898e-07
+    4.288219582850884e-07
+    3.592099155621433e-08
+    6.105128249344097e-08
+    1.731461630938217e-07
+    4.360776418997881e-07
+ 4.01e+10    
+    4.357439483987927e-07
+    1.731671599496303e-07
+    4.289530572013783e-07
+    6.106732141516658e-08
+     1.12103405012751e-07
+    4.289076256391507e-07
+    3.592050225442679e-08
+    6.107799701813909e-08
+    1.732261594416299e-07
+    4.361862080679946e-07
+ 4.02e+10    
+    4.358527780386537e-07
+    1.732471399351022e-07
+     4.29038774522757e-07
+    6.109380975449368e-08
+    1.121590856519911e-07
+    4.289934167405042e-07
+    3.591982666402948e-08
+    6.110459628681624e-08
+    1.733062310390594e-07
+    4.362949721531496e-07
+ 4.03e+10    
+    4.359618059689704e-07
+    1.733271946218305e-07
+    4.291246153862973e-07
+    6.112018226918014e-08
+    1.122147628156564e-07
+    4.290793315485207e-07
+    3.591896491718436e-08
+    6.113108015834796e-08
+     1.73386377711605e-07
+    4.364039342300869e-07
+ 4.04e+10    
+    4.360710322621599e-07
+    1.734073238326535e-07
+    4.292105797491129e-07
+    6.114643881766682e-08
+    1.122704363829097e-07
+     4.29165370022145e-07
+    3.591791714514599e-08
+    6.115744849053141e-08
+    1.734665992827883e-07
+    4.365130943715368e-07
+ 4.05e+10    
+    4.361804569886149e-07
+     1.73487527388477e-07
+    4.292966675680546e-07
+    6.117257925734225e-08
+    1.123261062333498e-07
+    4.292515321199232e-07
+    3.591668347829129e-08
+    6.118370114011712e-08
+    1.735468955741829e-07
+    4.366224526481583e-07
+ 4.06e+10    
+    4.362900802167316e-07
+     1.73567805108297e-07
+    4.293828787997336e-07
+      6.1198603444574e-08
+    1.123817722470304e-07
+    4.293378178000309e-07
+    3.591526404614937e-08
+    6.120983796283975e-08
+    1.736272664054396e-07
+     4.36732009128567e-07
+ 4.07e+10    
+    4.363999020129376e-07
+    1.736481568092248e-07
+    4.294692134005512e-07
+    6.122451123473969e-08
+    1.124374343044793e-07
+    4.294242270202998e-07
+    3.591365897743147e-08
+    6.123585881344942e-08
+      1.7370771159431e-07
+    4.368417638793632e-07
+ 4.08e+10    
+    4.365099224417198e-07
+     1.73728582306511e-07
+    4.295556713267197e-07
+     6.12503024822581e-08
+    1.124930922867164e-07
+    4.295107597382417e-07
+    3.591186840006128e-08
+    6.126176354574273e-08
+    1.737882309566708e-07
+     4.36951716965163e-07
+ 4.09e+10    
+    4.366201415656532e-07
+    1.738090814135681e-07
+    4.296422525342874e-07
+    6.127597704061996e-08
+     1.12548746075271e-07
+    4.295974159110759e-07
+    3.590989244120548e-08
+    6.128755201259353e-08
+    1.738688243065475e-07
+    4.370618684486253e-07
+ 4.1e+10     
+    4.367305594454278e-07
+    1.738896539419939e-07
+    4.297289569791617e-07
+    6.130153476241887e-08
+    1.126043955521999e-07
+    4.296841954957518e-07
+    3.590773122730434e-08
+    6.131322406598367e-08
+    1.739494914561374e-07
+    4.371722183904803e-07
+ 4.11e+10    
+    4.368411761398735e-07
+    1.739702997015937e-07
+    4.298157846171284e-07
+    6.132697549938175e-08
+    1.126600406001034e-07
+    4.297710984489723e-07
+    3.590538488410258e-08
+    6.133877955703357e-08
+    1.740302322158321e-07
+    4.372827668495577e-07
+ 4.12e+10    
+    4.369519917059925e-07
+    1.740510185004028e-07
+    4.299027354038745e-07
+    6.135229910239946e-08
+    1.127156811021423e-07
+    4.298581247272142e-07
+    3.590285353668048e-08
+    6.136421833603266e-08
+      1.7411104639424e-07
+    4.373935138828134e-07
+ 4.13e+10    
+    4.370630061989792e-07
+     1.74131810144708e-07
+     4.29989809295008e-07
+    6.137750542155726e-08
+    1.127713169420531e-07
+    4.299452742867533e-07
+    3.590013730948512e-08
+    6.138954025246985e-08
+    1.741919337982086e-07
+    4.375044595453591e-07
+ 4.14e+10    
+    4.371742196722508e-07
+    1.742126744390685e-07
+    4.300770062460735e-07
+    6.140259430616494e-08
+    1.128269480041644e-07
+    4.300325470836817e-07
+    3.589723632636175e-08
+    6.141474515506366e-08
+    1.742728942328453e-07
+    4.376156038904865e-07
+ 4.15e+10    
+    4.372856321774728e-07
+    1.742936111863379e-07
+    4.301643262125743e-07
+    6.142756560478722e-08
+     1.12882574173411e-07
+    4.301199430739295e-07
+    3.589415071058543e-08
+    6.143983289179214e-08
+    1.743539275015395e-07
+    4.377269469696961e-07
+ 4.16e+10    
+    4.373972437645844e-07
+    1.743746201876839e-07
+    4.302517691499872e-07
+    6.145241916527353e-08
+    1.129381953353494e-07
+    4.302074622132827e-07
+     3.58908805848928e-08
+    6.146480330992326e-08
+    1.744350334059829e-07
+    4.378384888327238e-07
+ 4.17e+10    
+    4.375090544818228e-07
+    1.744557012426089e-07
+    4.303393350137787e-07
+    6.147715483478808e-08
+    1.129938113761716e-07
+    4.302951044574026e-07
+    3.588742607151392e-08
+     6.14896562560443e-08
+    1.745162117461902e-07
+    4.379502295275653e-07
+ 4.18e+10    
+    4.376210643757504e-07
+    1.745368541489702e-07
+    4.304270237594238e-07
+    6.150177245983963e-08
+    1.130494221827191e-07
+    4.303828697618424e-07
+    3.588378729220446e-08
+    6.151439157609193e-08
+    1.745974623205192e-07
+    4.380621691005049e-07
+ 4.19e+10    
+    4.377332734912783e-07
+    1.746180787029989e-07
+    4.305148353424144e-07
+    6.152627188631112e-08
+    1.131050276424966e-07
+    4.304707580820651e-07
+    3.587996436827783e-08
+    6.153900911538142e-08
+    1.746787849256909e-07
+    4.381743075961377e-07
+ 4.2e+10     
+    4.378456818716928e-07
+      1.7469937469932e-07
+    4.306027697182819e-07
+    6.155065295948938e-08
+    1.131606276436848e-07
+    4.305587693734596e-07
+    3.587595742063763e-08
+    6.156350871863659e-08
+    1.747601793568089e-07
+    4.382866450573997e-07
+ 4.21e+10    
+    4.379582895586779e-07
+    1.747807419309704e-07
+    4.306908268426034e-07
+    6.157491552409437e-08
+    1.132162220751538e-07
+     4.30646903591356e-07
+    3.587176656981006e-08
+    6.158789023001867e-08
+    1.748416454073782e-07
+     4.38399181525588e-07
+ 4.22e+10    
+    4.380710965923398e-07
+    1.748621801894182e-07
+    4.307790066710187e-07
+    6.159905942430859e-08
+    1.132718108264747e-07
+    4.307351606910411e-07
+    3.586739193597664e-08
+    6.161215349315584e-08
+     1.74923182869325e-07
+    4.385119170403895e-07
+ 4.23e+10    
+    4.381841030112326e-07
+    1.749436892645807e-07
+    4.308673091592412e-07
+    6.162308450380626e-08
+    1.133273937879325e-07
+     4.30823540627772e-07
+    3.586283363900693e-08
+    6.163629835117215e-08
+     1.75004791533014e-07
+    4.386248516399044e-07
+ 4.24e+10    
+    4.382973088523806e-07
+    1.750252689448428e-07
+    4.309557342630692e-07
+    6.164699060578247e-08
+    1.133829708505376e-07
+    4.309120433567912e-07
+    3.585809179849152e-08
+    6.166032464671665e-08
+    1.750864711872681e-07
+    4.387379853606693e-07
+ 4.25e+10    
+    4.384107141513003e-07
+    1.751069190170738e-07
+    4.310442819383985e-07
+    6.167077757298201e-08
+    1.134385419060371e-07
+    4.310006688333391e-07
+    3.585316653377487e-08
+    6.168423222199216e-08
+    1.751682216193853e-07
+     4.38851318237684e-07
+ 4.26e+10    
+    4.385243189420281e-07
+     1.75188639266646e-07
+    4.311329521412312e-07
+    6.169444524772828e-08
+    1.134941068469261e-07
+    4.310894170126662e-07
+    3.584805796398856e-08
+    6.170802091878383e-08
+    1.752500426151565e-07
+    4.389648503044326e-07
+ 4.27e+10    
+    4.386381232571385e-07
+    1.752704294774504e-07
+    4.312217448276849e-07
+    6.171799347195189e-08
+    1.135496655664585e-07
+    4.311782878500465e-07
+    3.584276620808448e-08
+    6.173169057848807e-08
+     1.75331933958884e-07
+    4.390785815929101e-07
+ 4.28e+10    
+    4.387521271277695e-07
+    1.753522894319151e-07
+    4.313106599540048e-07
+    6.174142208721958e-08
+    1.136052179586579e-07
+    4.312672813007893e-07
+    3.583729138486817e-08
+    6.175524104214076e-08
+     1.75413895433397e-07
+    4.391925121336427e-07
+ 4.29e+10    
+    4.388663305836438e-07
+    1.754342189110206e-07
+    4.313996974765705e-07
+    6.176473093476213e-08
+    1.136607639183273e-07
+    4.313563973202485e-07
+    3.583163361303215e-08
+    6.177867215044572e-08
+    1.754959268200698e-07
+    4.393066419557136e-07
+ 4.3e+10     
+    4.389807336530919e-07
+     1.75516217694317e-07
+    4.314888573519058e-07
+    6.178791985550332e-08
+    1.137163033410593e-07
+    4.314456358638349e-07
+    3.582579301118961e-08
+    6.180198374380296e-08
+    1.755780278988376e-07
+    4.394209710867856e-07
+ 4.31e+10    
+    4.390953363630747e-07
+    1.755982855599395e-07
+    4.315781395366844e-07
+    6.181098869008775e-08
+    1.137718361232461e-07
+    4.315349968870277e-07
+    3.581976969790786e-08
+    6.182517566233668e-08
+    1.756601984482132e-07
+     4.39535499553121e-07
+ 4.32e+10    
+    4.392101387392035e-07
+    1.756804222846243e-07
+    4.316675439877396e-07
+    6.183393727890896e-08
+    1.138273621620884e-07
+    4.316244803453796e-07
+    3.581356379174205e-08
+    6.184824774592343e-08
+    1.757424382453031e-07
+    4.396502273796083e-07
+ 4.33e+10    
+    4.393251408057621e-07
+    1.757626276437246e-07
+     4.31757070662071e-07
+    6.185676546213774e-08
+     1.13882881355605e-07
+    4.317140861945328e-07
+    3.580717541126896e-08
+    6.187119983421974e-08
+    1.758247470658231e-07
+    4.397651545897808e-07
+ 4.34e+10    
+    4.394403425857297e-07
+    1.758449014112251e-07
+    4.318467195168504e-07
+    6.187947307974957e-08
+    1.139383936026417e-07
+    4.318038143902222e-07
+    3.580060467512082e-08
+    6.189403176669017e-08
+    1.759071246841143e-07
+    4.398802812058412e-07
+ 4.35e+10    
+    4.395557441008003e-07
+     1.75927243359758e-07
+    4.319364905094267e-07
+    6.190205997155272e-08
+    1.139938988028796e-07
+    4.318936648882871e-07
+    3.579385170201914e-08
+    6.191674338263455e-08
+    1.759895708731576e-07
+    4.399956072486811e-07
+ 4.36e+10    
+    4.396713453714027e-07
+    1.760096532606168e-07
+    4.320263835973368e-07
+    6.192452597721563e-08
+     1.14049396856844e-07
+    4.319836376446788e-07
+    3.578691661080874e-08
+    6.193933452121581e-08
+    1.760720854045901e-07
+     4.40111132737904e-07
+ 4.37e+10    
+    4.397871464167251e-07
+    1.760921308837722e-07
+    4.321163987383048e-07
+    6.194687093629445e-08
+    1.141048876659124e-07
+    4.320737326154671e-07
+    3.577979952049171e-08
+    6.196180502148723e-08
+    1.761546680487192e-07
+    4.402268576918476e-07
+ 4.38e+10    
+    4.399031472547303e-07
+    1.761746759978854e-07
+    4.322065358902522e-07
+    6.196909468826061e-08
+    1.141603711323225e-07
+      4.3216394975685e-07
+    3.577250055026151e-08
+     6.19841547224196e-08
+    1.762373185745368e-07
+    4.403427821276011e-07
+ 4.39e+10    
+    4.400193479021804e-07
+    1.762572883703228e-07
+    4.322967950112989e-07
+    6.199119707252783e-08
+    1.142158471591799e-07
+      4.3225428902516e-07
+    3.576501981953702e-08
+    6.200638346292851e-08
+    1.763200367497353e-07
+    4.404589060610301e-07
+ 4.4e+10     
+    4.401357483746529e-07
+    1.763399677671696e-07
+    4.323871760597707e-07
+     6.20131779284793e-08
+    1.142713156504657e-07
+    4.323447503768686e-07
+    3.575735744799671e-08
+    6.202849108190115e-08
+    1.764028223407199e-07
+    4.405752295067949e-07
+ 4.41e+10    
+    4.402523486865657e-07
+    1.764227139532446e-07
+    4.324776789942027e-07
+    6.203503709549487e-08
+    1.143267765110439e-07
+     4.32435333768597e-07
+    3.574951355561287e-08
+    6.205047741822344e-08
+    1.764856751126244e-07
+    4.406917524783712e-07
+ 4.42e+10    
+    4.403691488511889e-07
+    1.765055266921125e-07
+    4.325683037733421e-07
+    6.205677441297764e-08
+    1.143822296466683e-07
+    4.325260391571185e-07
+    3.574148826268573e-08
+    6.207234231080659e-08
+     1.76568594829324e-07
+    4.408084749880707e-07
+ 4.43e+10    
+    4.404861488806727e-07
+    1.765884057460978e-07
+     4.32659050356153e-07
+    6.207838972038101e-08
+    1.144376749639896e-07
+    4.326168664993657e-07
+     3.57332816898778e-08
+    6.209408559861377e-08
+    1.766515812534489e-07
+    4.409253970470613e-07
+ 4.44e+10    
+    4.406033487860599e-07
+    1.766713508762981e-07
+    4.327499187018195e-07
+    6.209988285723514e-08
+    1.144931123705624e-07
+    4.327078157524381e-07
+    3.572489395824802e-08
+    6.211570712068669e-08
+    1.767346341463986e-07
+    4.410425186653861e-07
+ 4.45e+10    
+    4.407207485773074e-07
+    1.767543618425971e-07
+    4.328409087697499e-07
+    6.212125366317343e-08
+    1.145485417748511e-07
+    4.327988868736027e-07
+    3.571632518928612e-08
+    6.213720671617198e-08
+    1.768177532683541e-07
+    4.411598398519831e-07
+ 4.46e+10    
+    4.408383482633071e-07
+    1.768374384036773e-07
+    4.329320205195771e-07
+    6.214250197795918e-08
+    1.146039630862369e-07
+    4.328900798203051e-07
+    3.570757550494686e-08
+    6.215858422434728e-08
+    1.769009383782916e-07
+    4.412773606147039e-07
+ 4.47e+10    
+    4.409561478518996e-07
+    1.769205803170325e-07
+    4.330232539111642e-07
+    6.216362764151153e-08
+    1.146593762150237e-07
+    4.329813945501685e-07
+     3.56986450276844e-08
+    6.217983948464757e-08
+    1.769841892339952e-07
+    4.413950809603343e-07
+ 4.48e+10    
+    4.410741473498963e-07
+    1.770037873389805e-07
+    4.331146089046052e-07
+    6.218463049393177e-08
+     1.14714781072444e-07
+    4.330728310210022e-07
+    3.568953388048648e-08
+    6.220097233669114e-08
+    1.770675055920698e-07
+    4.415130008946128e-07
+ 4.49e+10    
+    4.411923467630962e-07
+    1.770870592246757e-07
+     4.33206085460228e-07
+    6.220551037552935e-08
+     1.14770177570665e-07
+    4.331643891908044e-07
+    3.568024218690883e-08
+    6.222198262030542e-08
+    1.771508872079531e-07
+    4.416311204222475e-07
+ 4.5e+10     
+    4.413107460963032e-07
+    1.771703957281204e-07
+    4.332976835385971e-07
+    6.222626712684772e-08
+    1.148255656227942e-07
+    4.332560690177662e-07
+    3.567077007110937e-08
+    6.224287017555282e-08
+    1.772343338359283e-07
+    4.417494395469368e-07
+ 4.51e+10    
+    4.414293453533455e-07
+    1.772537966021774e-07
+    4.333894031005133e-07
+    6.224690058869018e-08
+    1.148809451428848e-07
+     4.33347870460277e-07
+    3.566111765788255e-08
+    6.226363484275616e-08
+    1.773178452291367e-07
+    4.418679582713855e-07
+ 4.52e+10    
+    4.415481445370909e-07
+    1.773372615985815e-07
+    4.334812441070182e-07
+    6.226741060214536e-08
+    1.149363160459414e-07
+    4.334397934769256e-07
+    3.565128507269355e-08
+    6.228427646252448e-08
+    1.774014211395888e-07
+    4.419866765973254e-07
+ 4.53e+10    
+    4.416671436494665e-07
+    1.774207904679517e-07
+    4.335732065193949e-07
+    6.228779700861294e-08
+    1.149916782479247e-07
+    4.335318380265061e-07
+    3.564127244171261e-08
+    6.230479487577824e-08
+    1.774850613181768e-07
+    4.421055945255309e-07
+ 4.54e+10    
+    4.417863426914729e-07
+    1.775043829598018e-07
+    4.336652902991689e-07
+    6.230805964982889e-08
+    1.150470316657574e-07
+    4.336240040680208e-07
+    3.563107989184914e-08
+    6.232518992377459e-08
+    1.775687655146864e-07
+    4.422247120558381e-07
+ 4.55e+10    
+    4.419057416632043e-07
+    1.775880388225524e-07
+    4.337574954081088e-07
+    6.232819836789063e-08
+    1.151023762173278e-07
+    4.337162915606815e-07
+    3.562070755078593e-08
+    6.234546144813241e-08
+    1.776525334778076e-07
+    4.423440291871605e-07
+ 4.56e+10    
+    4.420253405638637e-07
+    1.776717578035422e-07
+    4.338498218082305e-07
+    6.234821300528255e-08
+     1.15157711821496e-07
+    4.338087004639151e-07
+    3.561015554701336e-08
+    6.236560929085759e-08
+    1.777363649551471e-07
+    4.424635459175088e-07
+ 4.57e+10    
+    4.421451393917782e-07
+    1.777555396490385e-07
+    4.339422694617946e-07
+    6.236810340490059e-08
+    1.152130383980981e-07
+    4.339012307373658e-07
+    3.559942400986347e-08
+    6.238563329436758e-08
+    1.778202596932391e-07
+    4.425832622440063e-07
+ 4.58e+10    
+    4.422651381444185e-07
+    1.778393841042489e-07
+      4.3403483833131e-07
+    6.238786941007729e-08
+      1.1526835586795e-07
+    4.339938823408954e-07
+    3.558851306954397e-08
+    6.240553330151637e-08
+    1.779042174375558e-07
+     4.42703178162905e-07
+ 4.59e+10    
+    4.423853368184112e-07
+    1.779232909133311e-07
+    4.341275283795335e-07
+    6.240751086460648e-08
+     1.15323664152853e-07
+    4.340866552345895e-07
+    3.557742285717231e-08
+    6.242530915561889e-08
+    1.779882379325194e-07
+    4.428232936696037e-07
+ 4.6e+10     
+    4.425057354095585e-07
+    1.780072598194045e-07
+    4.342203395694703e-07
+    6.242702761276805e-08
+     1.15378963175597e-07
+    4.341795493787575e-07
+    3.556615350480964e-08
+    6.244496070047571e-08
+    1.780723209215123e-07
+    4.429436087586649e-07
+ 4.61e+10    
+    4.426263339128514e-07
+    1.780912905645603e-07
+    4.343132718643761e-07
+    6.244641949935221e-08
+    1.154342528599656e-07
+    4.342725647339351e-07
+    3.555470514549472e-08
+    6.246448778039723e-08
+    1.781564661468883e-07
+    4.430641234238292e-07
+ 4.62e+10    
+    4.427471323224872e-07
+    1.781753828898719e-07
+    4.344063252277568e-07
+    6.246568636968391e-08
+    1.154895331307392e-07
+    4.343657012608881e-07
+    3.554307791327774e-08
+    6.248389024022802e-08
+    1.782406733499826e-07
+    4.431848376580334e-07
+ 4.63e+10    
+    4.428681306318821e-07
+    1.782595365354049e-07
+    4.344994996233671e-07
+    6.248482806964708e-08
+    1.155448039136997e-07
+    4.344589589206112e-07
+    3.553127194325405e-08
+    6.250316792537077e-08
+    1.783249422711224e-07
+    4.433057514534252e-07
+ 4.64e+10    
+     4.42989328833691e-07
+    1.783437512402284e-07
+    4.345927950152162e-07
+    6.250384444570895e-08
+    1.156000651356342e-07
+    4.345523376743349e-07
+    3.551928737159799e-08
+    6.252232068181045e-08
+    1.784092726496374e-07
+    4.434268648013781e-07
+ 4.65e+10    
+    4.431107269198186e-07
+    1.784280267424235e-07
+    4.346862113675614e-07
+    6.252273534494352e-08
+    1.156553167243382e-07
+    4.346458374835216e-07
+    3.550712433559635e-08
+    6.254134835613791e-08
+      1.7849366422387e-07
+    4.435481776925093e-07
+ 4.66e+10    
+    4.432323248814356e-07
+    1.785123627790945e-07
+    4.347797486449131e-07
+    6.254150061505568e-08
+    1.157105586086196e-07
+    4.347394583098714e-07
+    3.549478297368207e-08
+    6.256025079557381e-08
+    1.785781167311853e-07
+    4.436696901166943e-07
+ 4.67e+10    
+    4.433541227089939e-07
+    1.785967590863777e-07
+    4.348734068120335e-07
+    6.256014010440491e-08
+    1.157657907183022e-07
+    4.348332001153228e-07
+    3.548226342546758e-08
+    6.257902784799193e-08
+    1.786626299079807e-07
+    4.437914020630806e-07
+ 4.68e+10    
+    4.434761203922411e-07
+     1.78681215399452e-07
+    4.349671858339368e-07
+    6.257865366202879e-08
+    1.158210129842292e-07
+    4.349270628620528e-07
+    3.546956583177823e-08
+    6.259767936194283e-08
+    1.787472034896966e-07
+    4.439133135201036e-07
+ 4.69e+10    
+    4.435983179202348e-07
+    1.787657314525482e-07
+    4.350610856758896e-07
+    6.259704113766639e-08
+    1.158762253382662e-07
+    4.350210465124803e-07
+    3.545669033468558e-08
+    6.261620518667701e-08
+     1.78831837210825e-07
+    4.440354244755025e-07
+ 4.7e+10     
+    4.437207152813566e-07
+    1.788503069789578e-07
+    4.351551063034094e-07
+    6.261530238178146e-08
+    1.159314277133045e-07
+    4.351151510292666e-07
+    3.544363707754053e-08
+     6.26346051721681e-08
+    1.789165308049201e-07
+    4.441577349163338e-07
+ 4.71e+10    
+     4.43843312463326e-07
+    1.789349417110436e-07
+    4.352492476822684e-07
+    6.263343724558582e-08
+    1.159866200432645e-07
+    4.352093763753162e-07
+    3.543040620500644e-08
+    6.265287916913595e-08
+    1.790012840046075e-07
+    4.442802448289863e-07
+ 4.72e+10    
+    4.439661094532152e-07
+    1.790196353802482e-07
+    4.353435097784883e-07
+    6.265144558106218e-08
+    1.160418022630985e-07
+    4.353037225137793e-07
+    3.541699786309202e-08
+    6.267102702906931e-08
+    1.790860965415931e-07
+    4.444029541991949e-07
+ 4.73e+10    
+    4.440891062374627e-07
+    1.791043877171033e-07
+    4.354378925583452e-07
+    6.266932724098696e-08
+    1.160969743087935e-07
+    4.353981894080515e-07
+    3.540341219918434e-08
+    6.268904860424893e-08
+    1.791709681466733e-07
+     4.44525863012055e-07
+ 4.74e+10    
+    4.442123028018854e-07
+    1.791891984512388e-07
+    4.355323959883652e-07
+    6.268708207895324e-08
+    1.161521361173745e-07
+    4.354927770217762e-07
+    3.538964936208134e-08
+    6.270694374776968e-08
+    1.792558985497432e-07
+    4.446489712520364e-07
+ 4.75e+10    
+    4.443356991316941e-07
+    1.792740673113921e-07
+    4.356270200353287e-07
+    6.270470994939325e-08
+    1.162072876269069e-07
+    4.355874853188448e-07
+    3.537570950202469e-08
+    6.272471231356363e-08
+    1.793408874798067e-07
+    4.447722789029984e-07
+ 4.76e+10    
+    4.444592952115063e-07
+    1.793589940254166e-07
+    4.357217646662655e-07
+    6.272221070760058e-08
+    1.162624287764993e-07
+    4.356823142633977e-07
+    3.536159277073213e-08
+    6.274235415642186e-08
+    1.794259346649848e-07
+    4.448957859482008e-07
+ 4.77e+10    
+    4.445830910253572e-07
+    1.794439783202906e-07
+    4.358166298484589e-07
+    6.273958420975297e-08
+    1.163175595063063e-07
+    4.357772638198261e-07
+    3.534729932142986e-08
+     6.27598691320169e-08
+    1.795110398325246e-07
+    4.450194923703205e-07
+ 4.78e+10    
+    4.447070865567163e-07
+    1.795290199221265e-07
+    4.359116155494425e-07
+    6.275683031293408e-08
+    1.163726797575307e-07
+     4.35872333952772e-07
+     3.53328293088848e-08
+    6.277725709692474e-08
+    1.795962027088083e-07
+    4.451433981514617e-07
+ 4.79e+10    
+    4.448312817884964e-07
+    1.796141185561784e-07
+    4.360067217370023e-07
+    6.277394887515569e-08
+    1.164277894724265e-07
+    4.359675246271292e-07
+    3.531818288943666e-08
+    6.279451790864674e-08
+    1.796814230193619e-07
+    4.452675032731722e-07
+ 4.8e+10     
+    4.449556767030708e-07
+    1.796992739468523e-07
+    4.361019483791753e-07
+    6.279093975537963e-08
+    1.164828885943008e-07
+    4.360628358080447e-07
+    3.530336022102998e-08
+    6.281165142563157e-08
+    1.797667004888639e-07
+    4.453918077164539e-07
+ 4.81e+10    
+    4.450802712822799e-07
+    1.797844858177126e-07
+    4.361972954442494e-07
+    6.280780281353925e-08
+    1.165379770675164e-07
+    4.361582674609189e-07
+    3.528836146324568e-08
+     6.28286575072964e-08
+    1.798520348411536e-07
+    4.455163114617769e-07
+ 4.82e+10    
+    4.452050655074486e-07
+    1.798697538914921e-07
+    4.362927629007619e-07
+    6.282453791056149e-08
+     1.16593054837494e-07
+     4.36253819551406e-07
+    3.527318677733307e-08
+    6.284553601404884e-08
+    1.799374257992398e-07
+    4.456410144890918e-07
+ 4.83e+10    
+    4.453300593593965e-07
+    1.799550778900993e-07
+    4.363883507175031e-07
+    6.284114490838785e-08
+    1.166481218507144e-07
+    4.363494920454154e-07
+    3.525783632624103e-08
+    6.286228680730807e-08
+    1.800228730853086e-07
+    4.457659167778422e-07
+ 4.84e+10    
+    4.454552528184505e-07
+    1.800404575346276e-07
+    4.364840588635121e-07
+    6.285762366999601e-08
+    1.167031780547207e-07
+    4.364452849091126e-07
+    3.524231027464958e-08
+    6.287890974952613e-08
+    1.801083764207328e-07
+    4.458910183069777e-07
+ 4.85e+10    
+    4.455806458644557e-07
+    1.801258925453624e-07
+    4.365798873080785e-07
+    6.287397405942089e-08
+    1.167582233981205e-07
+    4.365411981089188e-07
+    3.522660878900088e-08
+    6.289540470420877e-08
+    1.801939355260791e-07
+    4.460163190549655e-07
+ 4.86e+10    
+    4.457062384767875e-07
+    1.802113826417894e-07
+    4.366758360207422e-07
+    6.289019594177564e-08
+    1.168132578305873e-07
+    4.366372316115125e-07
+    3.521073203753032e-08
+    6.291177153593668e-08
+    1.802795501211168e-07
+    4.461418189998022e-07
+ 4.87e+10    
+    4.458320306343649e-07
+    1.802969275426039e-07
+    4.367719049712923e-07
+     6.29062891832726e-08
+    1.168682813028634e-07
+    4.367333853838292e-07
+     3.51946801902974e-08
+    6.292801011038592e-08
+    1.803652199248253e-07
+    4.462675181190268e-07
+ 4.88e+10    
+     4.45958022315659e-07
+    1.803825269657169e-07
+     4.36868094129769e-07
+    6.292225365124384e-08
+     1.16923293766761e-07
+    4.368296593930628e-07
+    3.517845341921625e-08
+     6.29441202943488e-08
+    1.804509446554028e-07
+    4.463934163897312e-07
+ 4.89e+10    
+     4.46084213498707e-07
+    1.804681806282639e-07
+    4.369644034664594e-07
+    6.293808921416195e-08
+    1.169782951751647e-07
+    4.369260536066659e-07
+    3.516205189808626e-08
+    6.296010195575411e-08
+    1.805367240302739e-07
+    4.465195137885736e-07
+ 4.9e+10     
+    4.462106041611218e-07
+    1.805538882466127e-07
+     4.37060832951902e-07
+    6.295379574166029e-08
+    1.170332854820325e-07
+    4.370225679923498e-07
+    3.514547580262225e-08
+    6.297595496368769e-08
+    1.806225577660969e-07
+    4.466458102917873e-07
+ 4.91e+10    
+    4.463371942801039e-07
+     1.80639649536371e-07
+    4.371573825568834e-07
+    6.296937310455342e-08
+    1.170882646423984e-07
+    4.371192025180865e-07
+     3.51287253104846e-08
+    6.299167918841222e-08
+    1.807084455787725e-07
+    4.467723058751949e-07
+ 4.92e+10    
+    4.464639838324515e-07
+    1.807254642123941e-07
+    4.372540522524401e-07
+    6.298482117485699e-08
+    1.171432326123733e-07
+     4.37215957152107e-07
+    3.511180060130927e-08
+    6.300727450138776e-08
+    1.807943871834508e-07
+    4.468990005142175e-07
+ 4.93e+10    
+    4.465909727945732e-07
+    1.808113319887927e-07
+    4.373508420098566e-07
+    6.300013982580798e-08
+    1.171981893491475e-07
+    4.373128318629036e-07
+    3.509470185673734e-08
+    6.302274077529105e-08
+    1.808803822945393e-07
+    4.470258941838868e-07
+ 4.94e+10    
+    4.467181611424941e-07
+    1.808972525789397e-07
+    4.374477518006667e-07
+    6.301532893188421e-08
+    1.172531348109915e-07
+    4.374098266192298e-07
+    3.507742926044461e-08
+    6.303807788403563e-08
+    1.809664306257103e-07
+    4.471529868588557e-07
+ 4.95e+10    
+    4.468455488518733e-07
+    1.809832256954786e-07
+     4.37544781596652e-07
+    6.303038836882424e-08
+    1.173080689572576e-07
+    4.375069413901014e-07
+    3.505998299817091e-08
+    6.305328570279119e-08
+    1.810525318899081e-07
+    4.472802785134084e-07
+ 4.96e+10    
+     4.46973135898007e-07
+    1.810692510503303e-07
+    4.376419313698437e-07
+    6.304531801364678e-08
+    1.173629917483821e-07
+    4.376041761447946e-07
+    3.504236325774916e-08
+      6.3068364108003e-08
+    1.811386857993571e-07
+    4.474077691214723e-07
+ 4.97e+10    
+    4.471009222558437e-07
+    1.811553283547006e-07
+    4.377392010925209e-07
+    6.306011774467001e-08
+    1.174179031458858e-07
+    4.377015308528496e-07
+    3.502457022913429e-08
+    6.308331297741125e-08
+    1.812248920655687e-07
+    4.475354586566275e-07
+ 4.98e+10    
+     4.47228907899993e-07
+    1.812414573190881e-07
+    4.378365907372114e-07
+    6.307478744153084e-08
+    1.174728031123764e-07
+    4.377990054840698e-07
+    3.500660410443189e-08
+    6.309813219007003e-08
+    1.813111503993485e-07
+    4.476633470921181e-07
+ 4.99e+10    
+    4.473570928047344e-07
+      1.8132763765329e-07
+    4.379341002766918e-07
+    6.308932698520393e-08
+    1.175276916115488e-07
+    4.378966000085219e-07
+    3.498846507792663e-08
+    6.311282162636626e-08
+    1.813974605108041e-07
+    4.477914344008612e-07
+ 5e+10       
+    4.474854769440287e-07
+     1.81413869066411e-07
+    4.380317296839861e-07
+     6.31037362580204e-08
+    1.175825686081871e-07
+     4.37994314396536e-07
+    3.497015334611045e-08
+    6.312738116803858e-08
+    1.814838221093514e-07
+    4.479197205554576e-07
+ 5.01e+10    
+    4.476140602915257e-07
+    1.815001512668691e-07
+    4.381294789323677e-07
+    6.311801514368683e-08
+    1.176374340681659e-07
+    4.380921486187077e-07
+    3.495166910771069e-08
+     6.31418106981959e-08
+    1.815702349037228e-07
+    4.480482055282021e-07
+ 5.02e+10    
+     4.47742842820577e-07
+    1.815864839624029e-07
+    4.382273479953584e-07
+    6.313216352730356e-08
+    1.176922879584511e-07
+    4.381901026458969e-07
+    3.493301256371757e-08
+    6.315611010133575e-08
+    1.816566986019732e-07
+    4.481768892910926e-07
+ 5.03e+10    
+    4.478718245042421e-07
+    1.816728668600796e-07
+    4.383253368467281e-07
+    6.314618129538328e-08
+    1.177471302471014e-07
+    4.382881764492294e-07
+    3.491418391741205e-08
+    6.317027926336284e-08
+    1.817432129114878e-07
+    4.483057718158408e-07
+ 5.04e+10    
+    4.480010053152997e-07
+    1.817592996663005e-07
+    4.384234454604949e-07
+    6.316006833586909e-08
+    1.178019609032692e-07
+    4.383863700000963e-07
+    3.489518337439281e-08
+    6.318431807160692e-08
+    1.818297775389888e-07
+    4.484348530738801e-07
+ 5.05e+10    
+    4.481303852262561e-07
+    1.818457820868092e-07
+    4.385216738109281e-07
+    6.317382453815278e-08
+    1.178567798972022e-07
+    4.384846832701559e-07
+    3.487601114260341e-08
+    6.319822641484097e-08
+    1.819163921905418e-07
+    4.485641330363769e-07
+ 5.06e+10    
+    4.482599642093547e-07
+    1.819323138266976e-07
+    4.386200218725425e-07
+    6.318744979309243e-08
+    1.179115872002438e-07
+     4.38583116231332e-07
+    3.485666743235905e-08
+    6.321200418329881e-08
+    1.820030565715635e-07
+    4.486936116742387e-07
+ 5.07e+10    
+    4.483897422365857e-07
+    1.820188945904128e-07
+    4.387184896201043e-07
+    6.320094399303059e-08
+    1.179663827848348e-07
+     4.38681668855818e-07
+    3.483715245637313e-08
+    6.322565126869306e-08
+    1.820897703868283e-07
+    4.488232889581234e-07
+ 5.08e+10    
+    4.485197192796931e-07
+    1.821055240817646e-07
+    4.388170770286281e-07
+    6.321430703181142e-08
+    1.180211666245139e-07
+    4.387803411160725e-07
+    3.481746642978339e-08
+    6.323916756423223e-08
+    1.821765333404742e-07
+    4.489531648584489e-07
+ 5.09e+10    
+    4.486498953101835e-07
+    1.821922020039312e-07
+    4.389157840733783e-07
+    6.322753880479826e-08
+    1.180759386939188e-07
+    4.388791329848241e-07
+    3.479760957017806e-08
+    6.325255296463845e-08
+    1.822633451360105e-07
+    4.490832393454017e-07
+ 5.1e+10     
+    4.487802702993383e-07
+    1.822789280594665e-07
+    4.390146107298679e-07
+    6.324063920889117e-08
+    1.181306989687874e-07
+    4.389780444350699e-07
+    3.477758209762157e-08
+    6.326580736616428e-08
+    1.823502054763242e-07
+    4.492135123889452e-07
+ 5.11e+10    
+    4.489108442182169e-07
+    1.823657019503064e-07
+    4.391135569738608e-07
+    6.325360814254351e-08
+    1.181854474259582e-07
+    4.390770754400761e-07
+     3.47573842346799e-08
+    6.327893066660994e-08
+     1.82437114063686e-07
+    4.493439839588289e-07
+ 5.12e+10    
+    4.490416170376694e-07
+    1.824525233777758e-07
+    4.392126227813705e-07
+    6.326644550577921e-08
+    1.182401840433718e-07
+    4.391762259733788e-07
+    3.473701620644598e-08
+    6.329192276534002e-08
+    1.825240705997575e-07
+    4.494746540245976e-07
+ 5.13e+10    
+    4.491725887283417e-07
+    1.825393920425947e-07
+    4.393118081286616e-07
+    6.327915120020944e-08
+    1.182949088000711e-07
+    4.392754960087842e-07
+    3.471647824056444e-08
+    6.330478356330029e-08
+    1.826110747855979e-07
+     4.49605522555598e-07
+ 5.14e+10    
+    4.493037592606862e-07
+    1.826263076448847e-07
+    4.394111129922486e-07
+    6.329172512904909e-08
+    1.183496216762023e-07
+    4.393748855203701e-07
+    3.469577056725636e-08
+    6.331751296303386e-08
+    1.826981263216692e-07
+    4.497365895209891e-07
+ 5.15e+10    
+    4.494351286049674e-07
+    1.827132698841757e-07
+    4.395105373488977e-07
+    6.330416719713329e-08
+    1.184043226530162e-07
+    4.394743944824855e-07
+    3.467489341934359e-08
+    6.333011086869789e-08
+    1.827852249078442e-07
+    4.498678548897491e-07
+ 5.16e+10    
+    4.495666967312727e-07
+    1.828002784594124e-07
+    4.396100811756263e-07
+    6.331647731093358e-08
+     1.18459011712868e-07
+    4.395740228697498e-07
+     3.46538470322728e-08
+    6.334257718607952e-08
+    1.828723702434117e-07
+    4.499993186306833e-07
+ 5.17e+10    
+    4.496984636095172e-07
+    1.828873330689598e-07
+    4.397097444497036e-07
+    6.332865537857398e-08
+    1.185136888392188e-07
+    4.396737706570578e-07
+    3.463263164413933e-08
+    6.335491182261188e-08
+    1.829595620270833e-07
+    4.501309807124332e-07
+ 5.18e+10    
+    4.498304292094526e-07
+    1.829744334106106e-07
+    4.398095271486509e-07
+    6.334070130984697e-08
+    1.185683540166358e-07
+     4.39773637819575e-07
+    3.461124749571064e-08
+    6.336711468738993e-08
+    1.830467999569997e-07
+    4.502628411034833e-07
+ 5.19e+10    
+    4.499625935006768e-07
+     1.83061579181591e-07
+     4.39909429250243e-07
+    6.335261501622908e-08
+    1.186230072307932e-07
+     4.39873624332742e-07
+    3.458969483044953e-08
+    6.337918569118608e-08
+    1.831340837307368e-07
+     4.50394899772169e-07
+ 5.2e+10     
+    4.500949564526375e-07
+    1.831487700785669e-07
+    4.400094507325065e-07
+    6.336439641089648e-08
+    1.186776484684729e-07
+    4.399737301722728e-07
+    3.456797389453695e-08
+    6.339112474646568e-08
+    1.832214130453118e-07
+    4.505271566866856e-07
+ 5.21e+10    
+     4.50227518034642e-07
+    1.832360057976499e-07
+    4.401095915737235e-07
+    6.337604540874048e-08
+    1.187322777175646e-07
+    4.400739553141566e-07
+    3.454608493689472e-08
+    6.340293176740234e-08
+    1.833087875971895e-07
+    4.506596118150931e-07
+ 5.22e+10    
+    4.503602782158643e-07
+    1.833232860344037e-07
+    4.402098517524273e-07
+    6.338756192638235e-08
+    1.187868949670668e-07
+    4.401742997346575e-07
+    3.452402820920764e-08
+    6.341460666989276e-08
+    1.833962070822883e-07
+     4.50792265125326e-07
+ 5.23e+10    
+    4.504932369653518e-07
+    1.834106104838509e-07
+      4.4031023124741e-07
+    6.339894588218899e-08
+    1.188415002070876e-07
+    4.402747634103176e-07
+    3.450180396594565e-08
+    6.342614937157224e-08
+    1.834836711959867e-07
+    4.509251165851993e-07
+ 5.24e+10    
+    4.506263942520325e-07
+    1.834979788404771e-07
+    4.404107300377144e-07
+    6.341019719628702e-08
+    1.188960934288444e-07
+    4.403753463179533e-07
+     3.44794124643854e-08
+    6.343755979182892e-08
+    1.835711796331289e-07
+     4.51058166162417e-07
+ 5.25e+10    
+    4.507597500447217e-07
+    1.835853907982397e-07
+    4.405113481026428e-07
+    6.342131579057803e-08
+    1.189506746246652e-07
+    4.404760484346597e-07
+    3.445685396463143e-08
+    6.344883785181852e-08
+      1.8365873208803e-07
+    4.511914138245762e-07
+ 5.26e+10    
+    4.508933043121292e-07
+    1.836728460505711e-07
+    4.406120854217513e-07
+    6.343230158875274e-08
+    1.190052437879883e-07
+    4.405768697378098e-07
+    3.443412872963753e-08
+    6.345998347447892e-08
+    1.837463282544842e-07
+    4.513248595391784e-07
+ 5.27e+10    
+    4.510270570228656e-07
+     1.83760344290387e-07
+     4.40712941974855e-07
+     6.34431545163055e-08
+    1.190598009133634e-07
+     4.40677810205055e-07
+    3.441123702522707e-08
+    6.347099658454417e-08
+    1.838339678257683e-07
+    4.514585032736325e-07
+ 5.28e+10    
+    4.511610081454492e-07
+    1.838478852100909e-07
+    4.408139177420251e-07
+    6.345387450054824e-08
+    1.191143459964518e-07
+    4.407788698143261e-07
+    3.438817912011361e-08
+    6.348187710855871e-08
+    1.839216504946492e-07
+    4.515923449952644e-07
+ 5.29e+10    
+    4.512951576483126e-07
+    1.839354685015802e-07
+    4.409150127035913e-07
+    6.346446147062458e-08
+    1.191688790340265e-07
+    4.408800485438344e-07
+     3.43649552859208e-08
+    6.349262497489109e-08
+    1.840093759533889e-07
+    4.517263846713202e-07
+ 5.3e+10     
+    4.514295054998086e-07
+     1.84023093856253e-07
+    4.410162268401434e-07
+    6.347491535752353e-08
+    1.192234000239729e-07
+    4.409813463720714e-07
+    3.434156579720213e-08
+    6.350324011374781e-08
+    1.840971438937508e-07
+    4.518606222689772e-07
+ 5.31e+10    
+    4.515640516682179e-07
+    1.841107609650126e-07
+    4.411175601325294e-07
+    6.348523609409308e-08
+    1.192779089652891e-07
+    4.410827632778103e-07
+     3.43180109314603e-08
+    6.351372245718671e-08
+    1.841849540070049e-07
+    4.519950577553463e-07
+ 5.32e+10    
+    4.516987961217529e-07
+    1.841984695182743e-07
+    4.412190125618587e-07
+    6.349542361505351e-08
+    1.193324058580858e-07
+    4.411842992401066e-07
+     3.42942909691662e-08
+    6.352407193913046e-08
+    1.842728059839343e-07
+    4.521296910974805e-07
+ 5.33e+10    
+    4.518337388285664e-07
+    1.842862192059707e-07
+    4.413205841095014e-07
+    6.350547785701086e-08
+    1.193868907035874e-07
+    4.412859542382991e-07
+    3.427040619377759e-08
+    6.353428849537951e-08
+    1.843606995148404e-07
+    4.522645222623812e-07
+ 5.34e+10    
+    4.519688797567554e-07
+    1.843740097175576e-07
+    4.414222747570894e-07
+    6.351539875846967e-08
+    1.194413635041314e-07
+    4.413877282520083e-07
+    3.424635689175752e-08
+    6.354437206362521e-08
+    1.844486342895485e-07
+     4.52399551217003e-07
+ 5.35e+10    
+    4.521042188743695e-07
+    1.844618407420195e-07
+    4.415240844865172e-07
+    6.352518625984608e-08
+     1.19495824263169e-07
+    4.414896212611419e-07
+    3.422214335259216e-08
+    6.355432258346253e-08
+    1.845366099974139e-07
+     4.52534777928261e-07
+ 5.36e+10    
+    4.522397561494139e-07
+    1.845497119678759e-07
+    4.416260132799432e-07
+    6.353484030348028e-08
+    1.195502729852655e-07
+    4.415916332458913e-07
+    3.419776586880854e-08
+    6.356413999640267e-08
+    1.846246263273273e-07
+    4.526702023630354e-07
+ 5.37e+10    
+    4.523754915498576e-07
+     1.84637623083186e-07
+    4.417280611197895e-07
+     6.35443608336492e-08
+    1.196047096761003e-07
+    4.416937641867334e-07
+    3.417322473599183e-08
+    6.357382424588553e-08
+    1.847126829677199e-07
+    4.528058244881788e-07
+ 5.38e+10    
+    4.525114250436373e-07
+    1.847255737755547e-07
+    4.418302279887439e-07
+    6.355374779657867e-08
+    1.196591343424669e-07
+    4.417960140644323e-07
+    3.414852025280215e-08
+    6.358337527729183e-08
+    1.848007796065699e-07
+    4.529416442705218e-07
+ 5.39e+10    
+    4.526475565986636e-07
+     1.84813563732139e-07
+    4.419325138697596e-07
+    6.356300114045557e-08
+    1.197135469922735e-07
+    4.418983828600408e-07
+    3.412365272099125e-08
+    6.359279303795518e-08
+    1.848889159314073e-07
+    4.530776616768767e-07
+ 5.4e+10     
+    4.527838861828278e-07
+    1.849015926396522e-07
+    4.420349187460568e-07
+     6.35721208154398e-08
+    1.197679476345428e-07
+    4.420008705548986e-07
+    3.409862244541866e-08
+     6.36020774771741e-08
+    1.849770916293196e-07
+    4.532138766740458e-07
+ 5.41e+10    
+    4.529204137640048e-07
+    1.849896601843704e-07
+    4.421374426011236e-07
+    6.358110677367597e-08
+    1.198223362794119e-07
+     4.42103477130635e-07
+    3.407342973406746e-08
+    6.361122854622346e-08
+    1.850653063869572e-07
+    4.533502892288246e-07
+ 5.42e+10    
+    4.530571393100595e-07
+    1.850777660521374e-07
+    4.422400854187169e-07
+    6.358995896930478e-08
+    1.198767129381331e-07
+     4.42206202569169e-07
+    3.404807489805986e-08
+    6.362024619836615e-08
+     1.85153559890539e-07
+    4.534868993080085e-07
+ 5.43e+10    
+    4.531940627888531e-07
+    1.851659099283707e-07
+    4.423428471828618e-07
+    6.359867735847484e-08
+    1.199310776230731e-07
+    4.423090468527113e-07
+    3.402255825167211e-08
+    6.362913038886416e-08
+    1.852418518258579e-07
+    4.536237068783978e-07
+ 5.44e+10    
+    4.533311841682463e-07
+    1.852540914980666e-07
+    4.424457278778557e-07
+    6.360726189935329e-08
+    1.199854303477135e-07
+    4.424120099637632e-07
+    3.399688011234948e-08
+    6.363788107498997e-08
+    1.853301818782857e-07
+    4.537607119068023e-07
+ 5.45e+10    
+    4.534685034161056e-07
+    1.853423104458055e-07
+    4.425487274882655e-07
+    6.361571255213716e-08
+    1.200397711266511e-07
+    4.425150918851199e-07
+    3.397104080072026e-08
+    6.364649821603724e-08
+    1.854185497327787e-07
+     4.53897914360047e-07
+ 5.46e+10    
+    4.536060205003078e-07
+    1.854305664557581e-07
+    4.426518459989322e-07
+    6.362402927906403e-08
+    1.200940999755973e-07
+    4.426182925998687e-07
+    3.394504064061006e-08
+    6.365498177333168e-08
+    1.855069550738834e-07
+    4.540353142049773e-07
+ 5.47e+10    
+    4.537437353887443e-07
+    1.855188592116895e-07
+    4.427550833949694e-07
+    6.363221204442258e-08
+    1.201484169113783e-07
+    4.427216120913921e-07
+     3.39188799590551e-08
+    6.366333171024142e-08
+     1.85595397585741e-07
+    4.541729114084622e-07
+ 5.48e+10    
+    4.538816480493275e-07
+    1.856071883969655e-07
+    4.428584396617648e-07
+    6.364026081456309e-08
+    1.202027219519351e-07
+     4.42825050343367e-07
+    3.389255908631567e-08
+    6.367154799218758e-08
+    1.856838769520937e-07
+    4.543107059374026e-07
+ 5.49e+10    
+    4.540197584499942e-07
+    1.856955536945576e-07
+    4.429619147849813e-07
+    6.364817555790764e-08
+    1.202570151163238e-07
+    4.429286073397679e-07
+    3.386607835588869e-08
+     6.36796305866543e-08
+     1.85772392856289e-07
+    4.544486977587313e-07
+ 5.5e+10     
+     4.54158066558709e-07
+    1.857839547870483e-07
+    4.430655087505588e-07
+    6.365595624495997e-08
+    1.203112964247145e-07
+    4.430322830648642e-07
+     3.38394381045203e-08
+    6.368757946319862e-08
+    1.858609449812851e-07
+    4.545868868394223e-07
+ 5.51e+10    
+    4.542965723434723e-07
+    1.858723913566365e-07
+    4.431692215447144e-07
+    6.366360284831564e-08
+    1.203655658983923e-07
+    4.431360775032249e-07
+    3.381263867221788e-08
+    6.369539459346049e-08
+     1.85949533009657e-07
+    4.547252731464924e-07
+ 5.52e+10    
+    4.544352757723219e-07
+    1.859608630851426e-07
+    4.432730531539436e-07
+    6.367111534267134e-08
+    1.204198235597567e-07
+    4.432399906397172e-07
+    3.378568040226158e-08
+    6.370307595117212e-08
+    1.860381566236002e-07
+    4.548638566470067e-07
+ 5.53e+10    
+    4.545741768133366e-07
+    1.860493696540132e-07
+     4.43377003565021e-07
+    6.367849370483448e-08
+    1.204740694323211e-07
+    4.433440224595077e-07
+    3.375856364121567e-08
+    6.371062351216751e-08
+    1.861268155049371e-07
+    4.550026373080826e-07
+ 5.54e+10    
+    4.547132754346443e-07
+    1.861379107443278e-07
+    4.434810727650026e-07
+    6.368573791373248e-08
+    1.205283035407134e-07
+     4.43448172948065e-07
+    3.373128873893942e-08
+    6.371803725439163e-08
+    1.862155093351215e-07
+     4.55141615096895e-07
+ 5.55e+10    
+    4.548525716044229e-07
+    1.862264860368022e-07
+    4.435852607412254e-07
+    6.369284795042172e-08
+    1.205825259106752e-07
+    4.435524420911581e-07
+    3.370385604859742e-08
+    6.372531715790933e-08
+    1.863042377952438e-07
+    4.552807899806792e-07
+ 5.56e+10    
+    4.549920652909051e-07
+    1.863150952117947e-07
+    4.436895674813084e-07
+    6.369982379809643e-08
+    1.206367365690617e-07
+    4.436568298748589e-07
+    3.367626592666971e-08
+    6.373246320491419e-08
+    1.863930005660362e-07
+    4.554201619267361e-07
+ 5.57e+10    
+    4.551317564623827e-07
+    1.864037379493112e-07
+    4.437939929731564e-07
+     6.37066654420974e-08
+    1.206909355438417e-07
+    4.437613362855434e-07
+    3.364851873296152e-08
+     6.37394753797373e-08
+    1.864817973278776e-07
+    4.555597309024364e-07
+ 5.58e+10    
+    4.552716450872112e-07
+    1.864924139290096e-07
+    4.438985372049578e-07
+    6.371337286992045e-08
+    1.207451228640971e-07
+    4.438659613098916e-07
+    3.362061483061231e-08
+    6.374635366885539e-08
+    1.865706277607986e-07
+     4.55699496875223e-07
+ 5.59e+10    
+    4.554117311338129e-07
+     1.86581122830206e-07
+    4.440032001651871e-07
+    6.371994607122466e-08
+    1.207992985600231e-07
+      4.4397070493489e-07
+    3.359255458610482e-08
+    6.375309806089931e-08
+    1.866594915444869e-07
+    4.558394598126168e-07
+ 5.6e+10     
+    4.555520145706795e-07
+    1.866698643318785e-07
+    4.441079818426074e-07
+    6.372638503784045e-08
+    1.208534626629271e-07
+    4.440755671478305e-07
+    3.356433836927334e-08
+     6.37597085466619e-08
+    1.867483883582919e-07
+    4.559796196822202e-07
+ 5.61e+10    
+    4.556924953663796e-07
+    1.867586381126731e-07
+    4.442128822262679e-07
+    6.373268976377747e-08
+    1.209076152052291e-07
+    4.441805479363132e-07
+    3.353596655331186e-08
+    6.376618511910587e-08
+    1.868373178812294e-07
+    4.561199764517191e-07
+ 5.62e+10    
+    4.558331734895583e-07
+    1.868474438509087e-07
+     4.44317901305509e-07
+    6.373886024523227e-08
+    1.209617562204609e-07
+    4.442856472882465e-07
+    3.350743951478165e-08
+    6.377252777337147e-08
+    1.869262797919876e-07
+    4.562605300888895e-07
+ 5.63e+10    
+    4.559740489089426e-07
+    1.869362812245816e-07
+    4.444230390699614e-07
+      6.3744896480596e-08
+    1.210158857432663e-07
+    4.443908651918492e-07
+    3.347875763361839e-08
+    6.377873650678394e-08
+    1.870152737689309e-07
+    4.564012805615986e-07
+ 5.64e+10    
+    4.561151215933452e-07
+    1.870251499113707e-07
+    4.445282955095481e-07
+    6.375079847046114e-08
+    1.210700038094002e-07
+    4.444962016356492e-07
+    3.344992129313907e-08
+    6.378481131886067e-08
+    1.871042994901052e-07
+    4.565422278378095e-07
+ 5.65e+10    
+    4.562563915116674e-07
+    1.871140495886428e-07
+    4.446336706144837e-07
+    6.375656621762925e-08
+    1.211241104557282e-07
+    4.446016566084866e-07
+    3.342093088004828e-08
+    6.379075221131835e-08
+    1.871933566332431e-07
+    4.566833718855844e-07
+ 5.66e+10    
+    4.563978586329025e-07
+    1.872029799334571e-07
+    4.447391643752793e-07
+    6.376219972711761e-08
+    1.211782057202269e-07
+    4.447072300995154e-07
+    3.339178678444424e-08
+     6.37965591880798e-08
+    1.872824448757685e-07
+    4.568247126730883e-07
+ 5.67e+10    
+    4.565395229261389e-07
+    1.872919406225702e-07
+    4.448447767827392e-07
+     6.37676990061657e-08
+    1.212322896419827e-07
+    4.448129220982015e-07
+     3.33624893998243e-08
+    6.380223225528052e-08
+    1.873715638948013e-07
+    4.569662501685919e-07
+ 5.68e+10    
+    4.566813843605642e-07
+    1.873809313324412e-07
+    4.449505078279656e-07
+    6.377306406424198e-08
+    1.212863622611916e-07
+    4.449187325943268e-07
+    3.333303912309003e-08
+    6.380777142127537e-08
+    1.874607133671626e-07
+    4.571079843404749e-07
+ 5.69e+10    
+    4.568234429054671e-07
+    1.874699517392364e-07
+    4.450563575023588e-07
+     6.37782949130501e-08
+    1.213404236191588e-07
+    4.450246615779877e-07
+    3.330343635455205e-08
+    6.381317669664462e-08
+    1.875498929693789e-07
+    4.572499151572296e-07
+ 5.7e+10     
+    4.569656985302419e-07
+    1.875590015188342e-07
+    4.451623257976171e-07
+    6.378339156653503e-08
+    1.213944737582984e-07
+    4.451307090395989e-07
+    3.327368149793417e-08
+     6.38184480942001e-08
+    1.876391023776878e-07
+    4.573920425874638e-07
+ 5.71e+10    
+    4.571081512043904e-07
+    1.876480803468302e-07
+     4.45268412705741e-07
+    6.378835404088896e-08
+    1.214485127221325e-07
+    4.452368749698921e-07
+    3.324377496037735e-08
+    6.382358562899119e-08
+    1.877283412680422e-07
+    4.575343665999029e-07
+ 5.72e+10    
+    4.572508008975255e-07
+    1.877371878985413e-07
+    4.453746182190298e-07
+    6.379318235455679e-08
+    1.215025405552906e-07
+    4.453431593599179e-07
+    3.321371715244305e-08
+    6.382858931831011e-08
+    1.878176093161148e-07
+    4.576768871633955e-07
+ 5.73e+10    
+    4.573936475793733e-07
+    1.878263238490114e-07
+    4.454809423300881e-07
+    6.379787652824221e-08
+    1.215565573035099e-07
+    4.454495622010478e-07
+    3.318350848811634e-08
+    6.383345918169792e-08
+    1.879069061973035e-07
+    4.578196042469126e-07
+ 5.74e+10    
+     4.57536691219778e-07
+    1.879154878730158e-07
+    4.455873850318227e-07
+     6.38024365849123e-08
+    1.216105630136336e-07
+    4.455560834849726e-07
+    3.315314938480849e-08
+     6.38381952409494e-08
+    1.879962315867358e-07
+    4.579625178195544e-07
+ 5.75e+10    
+     4.57679931788702e-07
+     1.88004679645066e-07
+    4.456939463174485e-07
+    6.380686254980317e-08
+    1.216645577336113e-07
+    4.456627232037076e-07
+    3.312264026335901e-08
+    6.384279752011828e-08
+    1.880855851592731e-07
+     4.58105627850549e-07
+ 5.76e+10    
+    4.578233692562289e-07
+    1.880938988394141e-07
+    4.458006261804833e-07
+     6.38111544504246e-08
+    1.217185415124976e-07
+    4.457694813495897e-07
+    3.309198154803752e-08
+    6.384726604552213e-08
+    1.881749665895165e-07
+    4.582489343092589e-07
+ 5.77e+10    
+    4.579670035925703e-07
+    1.881831451300582e-07
+    4.459074246147549e-07
+    6.381531231656494e-08
+    1.217725144004521e-07
+     4.45876357915281e-07
+    3.306117366654504e-08
+    6.385160084574691e-08
+    1.882643755518104e-07
+    4.583924371651816e-07
+ 5.78e+10    
+    4.581108347680617e-07
+    1.882724181907471e-07
+    4.460143416144008e-07
+    6.381933618029538e-08
+    1.218264764487385e-07
+    4.459833528937683e-07
+    3.303021705001483e-08
+    6.385580195165169e-08
+    1.883538117202475e-07
+    4.585361363879518e-07
+ 5.79e+10    
+     4.58254862753171e-07
+    1.883617176949838e-07
+    4.461213771738664e-07
+    6.382322607597457e-08
+    1.218804277097238e-07
+    4.460904662783661e-07
+    3.299911213301285e-08
+    6.385986939637269e-08
+    1.884432747686734e-07
+    4.586800319473451e-07
+ 5.8e+10     
+    4.583990875184967e-07
+    1.884510433160322e-07
+    4.462285312879111e-07
+    6.382698204025246e-08
+    1.219343682368779e-07
+    4.461976980627152e-07
+    3.296785935353789e-08
+    6.386380321532755e-08
+     1.88532764370692e-07
+    4.588241238132816e-07
+ 5.81e+10    
+    4.585435090347736e-07
+    1.885403947269202e-07
+    4.463358039516066e-07
+    6.383060411207444e-08
+    1.219882980847726e-07
+     4.46305048240786e-07
+    3.293645915302103e-08
+    6.386760344621912e-08
+    1.886222801996687e-07
+    4.589684119558241e-07
+ 5.82e+10    
+    4.586881272728727e-07
+    1.886297716004447e-07
+    4.464431951603382e-07
+    6.383409233268485e-08
+    1.220422173090813e-07
+    4.464125168068783e-07
+    3.290491197632488e-08
+    6.387127012903919e-08
+     1.88711821928736e-07
+    4.591128963451854e-07
+ 5.83e+10    
+     4.58832942203805e-07
+    1.887191736091768e-07
+     4.46550704909807e-07
+    6.383744674563076e-08
+    1.220961259665778e-07
+    4.465201037556239e-07
+    3.287321827174239e-08
+    6.387480330607199e-08
+    1.888013892307981e-07
+    4.592575769517277e-07
+ 5.84e+10    
+    4.589779537987229e-07
+    1.888086004254661e-07
+     4.46658333196031e-07
+    6.384066739676509e-08
+    1.221500241151359e-07
+     4.46627809081986e-07
+    3.284137849099501e-08
+    6.387820302189746e-08
+    1.888909817785349e-07
+    4.594024537459642e-07
+ 5.85e+10    
+    4.591231620289236e-07
+    1.888980517214452e-07
+    4.467660800153475e-07
+    6.384375433424977e-08
+    1.222039118137284e-07
+    4.467356327812599e-07
+    3.280939308923073e-08
+    6.388146932339445e-08
+    1.889805992444069e-07
+    4.595475266985649e-07
+ 5.86e+10    
+    4.592685668658481e-07
+     1.88987527169034e-07
+    4.468739453644105e-07
+    6.384670760855871e-08
+    1.222577891224263e-07
+    4.468435748490777e-07
+    3.277726252502143e-08
+    6.388460225974345e-08
+    1.890702413006599e-07
+    4.596927957803549e-07
+ 5.87e+10    
+    4.594141682810885e-07
+    1.890770264399453e-07
+    4.469819292401966e-07
+    6.384952727248054e-08
+    1.223116561023981e-07
+    4.469516352814047e-07
+    3.274498726035996e-08
+    6.388760188242944e-08
+    1.891599076193295e-07
+    4.598382609623182e-07
+ 5.88e+10    
+    4.595599662463853e-07
+    1.891665492056891e-07
+     4.47090031640005e-07
+    6.385221338112116e-08
+    1.223655128159093e-07
+    4.470598140745439e-07
+    3.271256776065672e-08
+    6.389046824524442e-08
+    1.892495978722449e-07
+    4.599839222155996e-07
+ 5.89e+10    
+     4.59705960733631e-07
+     1.89256095137576e-07
+    4.471982525614575e-07
+    6.385476599190592e-08
+    1.224193593263208e-07
+    4.471681112251356e-07
+    3.268000449473582e-08
+    6.389320140428956e-08
+    1.893393117310347e-07
+    4.601297795115066e-07
+ 5.9e+10     
+    4.598521517148734e-07
+    1.893456639067232e-07
+    4.473065920024991e-07
+     6.38571851645821e-08
+    1.224731956980882e-07
+    4.472765267301605e-07
+    3.264729793483083e-08
+    6.389580141797743e-08
+    1.894290488671304e-07
+    4.602758328215117e-07
+ 5.91e+10    
+    4.599985391623153e-07
+    1.894352551840584e-07
+    4.474150499614032e-07
+    6.385947096122036e-08
+    1.225270219967618e-07
+    4.473850605869369e-07
+    3.261444855658007e-08
+    6.389826834703399e-08
+     1.89518808951771e-07
+    4.604220821172529e-07
+ 5.92e+10    
+    4.601451230483173e-07
+    1.895248686403244e-07
+    4.475236264367689e-07
+    6.386162344621689e-08
+    1.225808382889842e-07
+    4.474937127931252e-07
+    3.258145683902153e-08
+    6.390060225450022e-08
+     1.89608591656008e-07
+    4.605685273705376e-07
+ 5.93e+10    
+    4.602919033454002e-07
+    1.896145039460837e-07
+    4.476323214275247e-07
+    6.386364268629497e-08
+    1.226346446424909e-07
+    4.476024833467294e-07
+    3.254832326458729e-08
+    6.390280320573361e-08
+    1.896983966507094e-07
+     4.60715168553342e-07
+ 5.94e+10    
+    4.604388800262454e-07
+     1.89704160771723e-07
+    4.477411349329286e-07
+    6.386552875050586e-08
+    1.226884411261081e-07
+    4.477113722460952e-07
+    3.251504831909752e-08
+    6.390487126840961e-08
+    1.897882236065642e-07
+    4.608620056378147e-07
+ 5.95e+10    
+     4.60586053063698e-07
+    1.897938387874577e-07
+      4.4785006695257e-07
+    6.386728171023052e-08
+    1.227422278097526e-07
+    4.478203794899135e-07
+    3.248163249175418e-08
+    6.390680651252272e-08
+    1.898780721940872e-07
+    4.610090385962786e-07
+ 5.96e+10    
+    4.607334224307665e-07
+    1.898835376633364e-07
+    4.479591174863715e-07
+    6.386890163918018e-08
+      1.2279600476443e-07
+    4.479295050772211e-07
+    3.244807627513404e-08
+    6.390860901038739e-08
+    1.899679420836229e-07
+    4.611562674012293e-07
+ 5.97e+10    
+    4.608809881006271e-07
+    1.899732570692451e-07
+    4.480682865345879e-07
+    6.387038861339738e-08
+    1.228497720622347e-07
+    4.480387490074021e-07
+    3.241438016518159e-08
+    6.391027883663887e-08
+    1.900578329453504e-07
+    4.613036920253411e-07
+ 5.98e+10    
+    4.610287500466232e-07
+    1.900629966749123e-07
+    4.481775740978116e-07
+    6.387174271125626e-08
+    1.229035297763478e-07
+    4.481481112801868e-07
+    3.238054466120119e-08
+    6.391181606823363e-08
+    1.901477444492873e-07
+    4.614513124414654e-07
+ 5.99e+10    
+    4.611767082422665e-07
+    1.901527561499131e-07
+    4.482869801769702e-07
+    6.387296401346325e-08
+     1.22957277981037e-07
+    4.482575918956576e-07
+    3.234657026584915e-08
+    6.391322078444995e-08
+    1.902376762652947e-07
+     4.61599128622634e-07
+ 6e+10       
+    4.613248626612407e-07
+    1.902425351636733e-07
+    4.483965047733286e-07
+    6.387405260305699e-08
+    1.230110167516549e-07
+    4.483671908542448e-07
+    3.231245748512503e-08
+     6.39144930668878e-08
+    1.903276280630814e-07
+    4.617471405420585e-07
+ 6.01e+10    
+    4.614732132774014e-07
+    1.903323333854743e-07
+    4.485061478884918e-07
+    6.387500856540835e-08
+    1.230647461646379e-07
+    4.484769081567313e-07
+    3.227820682836282e-08
+    6.391563299946901e-08
+    1.904175995122077e-07
+    4.618953481731339e-07
+ 6.02e+10    
+     4.61621760064777e-07
+    1.904221504844577e-07
+    4.486159095244064e-07
+    6.387583198822044e-08
+    1.231184662975057e-07
+    4.485867438042522e-07
+    3.224381880822148e-08
+    6.391664066843704e-08
+    1.905075902820907e-07
+    4.620437514894378e-07
+ 6.03e+10    
+    4.617705029975707e-07
+    1.905119861296293e-07
+    4.487257896833593e-07
+    6.387652296152795e-08
+    1.231721772288595e-07
+    4.486966977982969e-07
+    3.220929394067525e-08
+     6.39175161623566e-08
+    1.905976000420083e-07
+    4.621923504647351e-07
+ 6.04e+10    
+    4.619194420501634e-07
+    1.906018399898636e-07
+    4.488357883679808e-07
+     6.38770815776968e-08
+    1.232258790383812e-07
+    4.488067701407105e-07
+    3.217463274500333e-08
+    6.391825957211288e-08
+    1.906876284611033e-07
+    4.623411450729739e-07
+ 6.05e+10    
+     4.62068577197111e-07
+    1.906917117339083e-07
+    4.489459055812471e-07
+    6.387750793142311e-08
+    1.232795718068323e-07
+    4.489169608336925e-07
+    3.213983574377928e-08
+    6.391887099091097e-08
+    1.907776752083876e-07
+    4.624901352882926e-07
+ 6.06e+10    
+    4.622179084131502e-07
+    1.907816010303889e-07
+    4.490561413264794e-07
+    6.387780211973244e-08
+    1.233332556160523e-07
+    4.490272698798007e-07
+     3.21049034628601e-08
+    6.391935051427479e-08
+    1.908677399527479e-07
+    4.626393210850173e-07
+ 6.07e+10    
+    4.623674356731951e-07
+    1.908715075478124e-07
+    4.491664956073453e-07
+    6.387796424197851e-08
+     1.23386930548958e-07
+    4.491376972819525e-07
+    3.206983643137454e-08
+    6.391969824004589e-08
+     1.90957822362948e-07
+     4.62788702437663e-07
+ 6.08e+10    
+    4.625171589523427e-07
+    1.909614309545726e-07
+    4.492769684278632e-07
+     6.38779943998418e-08
+    1.234405966895417e-07
+    4.492482430434222e-07
+    3.203463518171146e-08
+    6.391991426838216e-08
+    1.910479221076347e-07
+     4.62938279320937e-07
+ 6.09e+10    
+     4.62667078225872e-07
+    1.910513709189539e-07
+    4.493875597923998e-07
+    6.387789269732829e-08
+    1.234942541228709e-07
+    4.493589071678482e-07
+    3.199930024950742e-08
+    6.391999870175626e-08
+    1.911380388553417e-07
+    4.630880517097381e-07
+ 6.1e+10     
+    4.628171934692427e-07
+    1.911413271091357e-07
+    4.494982697056731e-07
+    6.387765924076736e-08
+    1.235479029350859e-07
+    4.494696896592285e-07
+    3.196383217363395e-08
+     6.39199516449539e-08
+    1.912281722744933e-07
+    4.632380195791585e-07
+ 6.11e+10    
+    4.629675046581012e-07
+    1.912312991931969e-07
+    4.496090981727548e-07
+    6.387729413880998e-08
+    1.236015432133991e-07
+    4.495805905219253e-07
+    3.192823149618453e-08
+    6.391977320507185e-08
+    1.913183220334098e-07
+    4.633881829044838e-07
+ 6.12e+10    
+    4.631180117682777e-07
+    1.913212868391205e-07
+    4.497200451990702e-07
+    6.387679750242698e-08
+     1.23655175046094e-07
+    4.496916097606656e-07
+    3.189249876246113e-08
+    6.391946349151604e-08
+     1.91408487800311e-07
+    4.635385416611946e-07
+ 6.13e+10    
+     4.63268714775788e-07
+    1.914112897147972e-07
+    4.498311107903989e-07
+    6.387616944490604e-08
+    1.237087985225232e-07
+    4.498027473805403e-07
+    3.185663452096007e-08
+    6.391902261599888e-08
+    1.914986692433204e-07
+    4.636890958249684e-07
+ 6.14e+10    
+    4.634196136568352e-07
+    1.915013074880306e-07
+    4.499422949528785e-07
+    6.387541008184988e-08
+    1.237624137331075e-07
+    4.499140033870096e-07
+    3.182063932335794e-08
+    6.391845069253723e-08
+    1.915888660304706e-07
+    4.638398453716781e-07
+ 6.15e+10    
+    4.635707083878112e-07
+     1.91591339826541e-07
+    4.500535976930043e-07
+    6.387451953117326e-08
+    1.238160207693343e-07
+    4.500253777858991e-07
+    3.178451372449675e-08
+     6.39177478374494e-08
+    1.916790778297061e-07
+    4.639907902773963e-07
+ 6.16e+10    
+    4.637219989452956e-07
+    1.916813863979698e-07
+    4.501650190176302e-07
+    6.387349791310007e-08
+    1.238696197237565e-07
+    4.501368705834045e-07
+     3.17482582823688e-08
+    6.391691416935249e-08
+    1.917693043088885e-07
+    4.641419305183917e-07
+ 6.17e+10    
+    4.638734853060569e-07
+    1.917714468698842e-07
+    4.502765589339719e-07
+    6.387234535016069e-08
+    1.239232106899909e-07
+    4.502484817860928e-07
+    3.171187355810126e-08
+    6.391594980915933e-08
+    1.918595451358009e-07
+    4.642932660711339e-07
+ 6.18e+10    
+    4.640251674470554e-07
+     1.91861520909781e-07
+    4.503882174496064e-07
+    6.387106196718826e-08
+    1.239767937627167e-07
+    4.503602114009006e-07
+    3.167536011594008e-08
+    6.391485488007513e-08
+    1.919497999781516e-07
+    4.644447969122923e-07
+ 6.19e+10    
+    4.641770453454405e-07
+    1.919516081850911e-07
+    4.504999945724741e-07
+    6.386964789131557e-08
+    1.240303690376744e-07
+    4.504720594351383e-07
+    3.163871852323388e-08
+     6.39136295075943e-08
+    1.920400685035785e-07
+    4.645965230187362e-07
+ 6.2e+10     
+    4.643291189785553e-07
+     1.92041708363184e-07
+    4.506118903108799e-07
+    6.386810325197151e-08
+    1.240839366116637e-07
+    4.505840258964898e-07
+    3.160194935041708e-08
+    6.391227381949673e-08
+    1.921303503796538e-07
+    4.647484443675382e-07
+ 6.21e+10    
+    4.644813883239355e-07
+     1.92131821111372e-07
+    4.507239046734961e-07
+     6.38664281808772e-08
+    1.241374965825429e-07
+    4.506961107930135e-07
+    3.156505317099295e-08
+    6.391078794584408e-08
+    1.922206452738878e-07
+    4.649005609359709e-07
+ 6.22e+10    
+    4.646338533593079e-07
+    1.922219460969149e-07
+    4.508360376693614e-07
+    6.386462281204206e-08
+    1.241910490492269e-07
+    4.508083141331454e-07
+    3.152803056151594e-08
+    6.390917201897585e-08
+    1.923109528537333e-07
+    4.650528727015113e-07
+ 6.23e+10    
+    4.647865140625939e-07
+    1.923120829870224e-07
+    4.509482893078815e-07
+    6.386268728175963e-08
+    1.242445941116852e-07
+    4.509206359256972e-07
+      3.1490882101574e-08
+    6.390742617350516e-08
+    1.924012727865899e-07
+    4.652053796418387e-07
+ 6.24e+10    
+     4.64939370411911e-07
+    1.924022314488619e-07
+    4.510606595988365e-07
+    6.386062172860355e-08
+    1.242981318709415e-07
+    4.510330761798601e-07
+    3.145360837377035e-08
+    6.390555054631473e-08
+    1.924916047398083e-07
+     4.65358081734837e-07
+ 6.25e+10    
+    4.650924223855701e-07
+    1.924923911495591e-07
+    4.511731485523731e-07
+    6.385842629342264e-08
+    1.243516624290711e-07
+    4.511456349052047e-07
+    3.141620996370455e-08
+    6.390354527655204e-08
+    1.925819483806942e-07
+    4.655109789585945e-07
+ 6.26e+10    
+    4.652456699620779e-07
+     1.92582561756205e-07
+    4.512857561790142e-07
+    6.385610111933661e-08
+    1.244051858892001e-07
+    4.512583121116827e-07
+    3.137868745995395e-08
+    6.390141050562507e-08
+    1.926723033765136e-07
+    4.656640712914049e-07
+ 6.27e+10    
+    4.653991131201382e-07
+    1.926727429358589e-07
+    4.513984824896561e-07
+    6.385364635173113e-08
+    1.244587023555033e-07
+    4.513711078096283e-07
+    3.134104145405394e-08
+    6.389914637719724e-08
+    1.927626693944953e-07
+    4.658173587117675e-07
+ 6.28e+10    
+    4.655527518386503e-07
+    1.927629343555524e-07
+    4.515113274955684e-07
+     6.38510621382527e-08
+    1.245122119332026e-07
+    4.514840220097579e-07
+    3.130327254047838e-08
+    6.389675303718236e-08
+    1.928530461018368e-07
+     4.65970841198387e-07
+ 6.29e+10    
+    4.657065860967116e-07
+    1.928531356822949e-07
+     4.51624291208401e-07
+    6.384834862880356e-08
+    1.245657147285656e-07
+    4.515970547231731e-07
+    3.126538131661946e-08
+    6.389423063373977e-08
+    1.929434331657076e-07
+    4.661245187301755e-07
+ 6.3e+10     
+    4.658606158736168e-07
+    1.929433465830769e-07
+    4.517373736401783e-07
+    6.384550597553647e-08
+    1.246192108489041e-07
+    4.517102059613612e-07
+    3.122736838276719e-08
+    6.389157931726865e-08
+    1.930338302532536e-07
+    4.662783912862514e-07
+ 6.31e+10    
+    4.660148411488587e-07
+    1.930335667248745e-07
+     4.51850574803307e-07
+    6.384253433284886e-08
+    1.246727004025716e-07
+    4.518234757361962e-07
+    3.118923434208856e-08
+    6.388879924040278e-08
+    1.931242370316019e-07
+    4.664324588459414e-07
+ 6.32e+10    
+    4.661692619021301e-07
+    1.931237957746541e-07
+    4.519638947105732e-07
+    6.383943385737758e-08
+    1.247261834989631e-07
+    4.519368640599403e-07
+    3.115097980060632e-08
+    6.388589055800473e-08
+    1.932146531678639e-07
+     4.66586721388779e-07
+ 6.33e+10    
+      4.6632387811332e-07
+    1.932140333993758e-07
+    4.520773333751453e-07
+    6.383620470799254e-08
+    1.247796602485115e-07
+    4.520503709452443e-07
+    3.111260536717747e-08
+    6.388285342715997e-08
+     1.93305078329141e-07
+    4.667411788945071e-07
+ 6.34e+10    
+    4.664786897625196e-07
+    1.933042792659986e-07
+    4.521908908105748e-07
+    6.383284704579105e-08
+    1.248331307626875e-07
+    4.521639964051509e-07
+    3.107411165347125e-08
+    6.387968800717103e-08
+    1.933955121825274e-07
+    4.668958313430759e-07
+ 6.35e+10    
+    4.666336968300188e-07
+    1.933945330414844e-07
+     4.52304567030799e-07
+    6.382936103409159e-08
+    1.248865951539971e-07
+    4.522777404530932e-07
+      3.1035499273947e-08
+    6.387639445955114e-08
+    1.934859543951156e-07
+    4.670506787146458e-07
+ 6.36e+10    
+    4.667888992963066e-07
+    1.934847943928015e-07
+    4.524183620501406e-07
+      6.3825746838427e-08
+    1.249400535359796e-07
+    4.523916031028972e-07
+    3.099676884583138e-08
+    6.387297294801796e-08
+    1.935764046339995e-07
+    4.672057209895854e-07
+ 6.37e+10    
+    4.669442971420751e-07
+    1.935750629869302e-07
+    4.525322758833098e-07
+    6.382200462653869e-08
+    1.249935060232066e-07
+    4.525055843687829e-07
+    3.095792098909557e-08
+    6.386942363848711e-08
+    1.936668625662794e-07
+    4.673609581484736e-07
+ 6.38e+10    
+    4.670998903482155e-07
+    1.936653384908662e-07
+    4.526463085454052e-07
+    6.381813456836925e-08
+    1.250469527312794e-07
+    4.526196842653658e-07
+    3.091895632643181e-08
+    6.386574669906525e-08
+    1.937573278590659e-07
+    4.675163901720982e-07
+ 6.39e+10    
+    4.672556788958196e-07
+    1.937556205716247e-07
+    4.527604600519167e-07
+    6.381413683605598e-08
+    1.251003937768279e-07
+    4.527339028076582e-07
+    3.087987548322992e-08
+    6.386194230004375e-08
+    1.938478001794846e-07
+    4.676720170414587e-07
+ 6.4e+10     
+    4.674116627661826e-07
+    1.938459088962456e-07
+    4.528747304187248e-07
+    6.381001160392377e-08
+    1.251538292775079e-07
+    4.528482400110693e-07
+    3.084067908755316e-08
+    6.385801061389102e-08
+    1.939382791946797e-07
+    4.678278387377632e-07
+ 6.41e+10    
+    4.675678419407997e-07
+    1.939362031317966e-07
+    4.529891196621023e-07
+    6.380575904847782e-08
+    1.252072593520001e-07
+    4.529626958914071e-07
+    3.080136777011405e-08
+    6.385395181524592e-08
+    1.940287645718185e-07
+    4.679838552424318e-07
+ 6.42e+10    
+    4.677242164013692e-07
+    1.940265029453788e-07
+    4.531036277987178e-07
+    6.380137934839648e-08
+    1.252606841200078e-07
+    4.530772704648807e-07
+    3.076194216424966e-08
+    6.384976608091014e-08
+    1.941192559780958e-07
+    4.681400665370949e-07
+ 6.43e+10    
+    4.678807861297916e-07
+    1.941168080041297e-07
+     4.53218254845634e-07
+    6.379687268452359e-08
+    1.253141037022548e-07
+    4.531919637480981e-07
+    3.072240290589669e-08
+    6.384545358984077e-08
+    1.942097530807379e-07
+    4.682964726035937e-07
+ 6.44e+10    
+    4.680375511081693e-07
+    1.942071179752281e-07
+    4.533330008203102e-07
+    6.379223923986075e-08
+    1.253675182204839e-07
+    4.533067757580721e-07
+    3.068275063356612e-08
+    6.384101452314262e-08
+     1.94300255547007e-07
+    4.684530734239808e-07
+ 6.45e+10    
+    4.681945113188079e-07
+    1.942974325258983e-07
+    4.534478657406047e-07
+    6.378747919955978e-08
+    1.254209277974549e-07
+    4.534217065122182e-07
+    3.064298598831775e-08
+    6.383644906406064e-08
+    1.943907630442055e-07
+    4.686098689805204e-07
+ 6.46e+10    
+    4.683516667442166e-07
+    1.943877513234148e-07
+    4.535628496247744e-07
+    6.378259275091447e-08
+    1.254743325569422e-07
+     4.53536756028356e-07
+    3.060310961373413e-08
+    6.383175739797167e-08
+    1.944812752396801e-07
+    4.687668592556888e-07
+ 6.47e+10    
+    4.685090173671063e-07
+    1.944780740351055e-07
+    4.536779524914777e-07
+    6.377758008335258e-08
+    1.255277326237335e-07
+     4.53651924324712e-07
+    3.056312215589442e-08
+    6.382693971237656e-08
+    1.945717918008261e-07
+    4.689240442321732e-07
+ 6.48e+10    
+    4.686665631703927e-07
+    1.945684003283572e-07
+    4.537931743597756e-07
+    6.377244138842755e-08
+    1.255811281236273e-07
+    4.537672114199196e-07
+    3.052302426334783e-08
+    6.382199619689182e-08
+    1.946623123950916e-07
+    4.690814238928727e-07
+ 6.49e+10    
+    4.688243041371944e-07
+     1.94658729870619e-07
+    4.539085152491306e-07
+    6.376717685981002e-08
+    1.256345191834312e-07
+    4.538826173330206e-07
+    3.048281658708684e-08
+    6.381692704324119e-08
+    1.947528366899819e-07
+    4.692389982208995e-07
+ 6.5e+10     
+    4.689822402508334e-07
+    1.947490623294069e-07
+    4.540239751794114e-07
+    6.376178669327925e-08
+    1.256879059309596e-07
+    4.539981420834668e-07
+    3.044249978052004e-08
+    6.381173244524722e-08
+    1.948433643530637e-07
+    4.693967671995777e-07
+ 6.51e+10    
+     4.69140371494837e-07
+    1.948393973723084e-07
+    4.541395541708935e-07
+    6.375627108671445e-08
+    1.257412884950317e-07
+    4.541137856911196e-07
+    3.040207449944467e-08
+    6.380641259882239e-08
+    1.949338950519689e-07
+    4.695547308124425e-07
+ 6.52e+10    
+    4.692986978529352e-07
+    1.949297346669861e-07
+    4.542552522442576e-07
+    6.375063024008577e-08
+    1.257946670054698e-07
+    4.542295481762537e-07
+    3.036154140201894e-08
+    6.380096770196039e-08
+    1.950244284544001e-07
+    4.697128890432433e-07
+ 6.53e+10    
+    4.694572193090623e-07
+    1.950200738811825e-07
+    4.543710694205947e-07
+    6.374486435544541e-08
+    1.258480415930967e-07
+    4.543454295595561e-07
+    3.032090114873405e-08
+      6.3795397954727e-08
+    1.951149642281334e-07
+    4.698712418759411e-07
+ 6.54e+10    
+    4.696159358473581e-07
+    1.951104146827246e-07
+    4.544870057214066e-07
+    6.373897363691849e-08
+    1.259014123897342e-07
+    4.544614298621298e-07
+     3.02801544023859e-08
+     6.37897035592512e-08
+    1.952055020410237e-07
+    4.700297892947099e-07
+ 6.55e+10    
+     4.69774847452166e-07
+    1.952007567395271e-07
+    4.546030611686044e-07
+    6.373295829069339e-08
+    1.259547795282001e-07
+     4.54577549105491e-07
+    3.023930182804646e-08
+    6.378388471971548e-08
+    1.952960415610082e-07
+    4.701885312839362e-07
+ 6.56e+10    
+    4.699339541080339e-07
+    1.952910997195978e-07
+    4.547192357845135e-07
+    6.372681852501271e-08
+     1.26008143142307e-07
+    4.546937873115747e-07
+    3.019834409303504e-08
+    6.377794164234684e-08
+    1.953865824561118e-07
+    4.703474678282199e-07
+ 6.57e+10    
+     4.70093255799716e-07
+    1.953814432910414e-07
+    4.548355295918724e-07
+    6.372055455016348e-08
+    1.260615033668598e-07
+    4.548101445027335e-07
+    3.015728186688912e-08
+     6.37718745354069e-08
+      1.9547712439445e-07
+    4.705065989123728e-07
+ 6.58e+10    
+    4.702527525121685e-07
+    1.954717871220638e-07
+    4.549519426138369e-07
+    6.371416657846725e-08
+     1.26114860337653e-07
+    4.549266207017387e-07
+    3.011611582133495e-08
+    6.376568360918237e-08
+    1.955676670442343e-07
+    4.706659245214211e-07
+ 6.59e+10    
+    4.704124442305557e-07
+    1.955621308809766e-07
+    4.550684748739763e-07
+    6.370765482427058e-08
+    1.261682141914696e-07
+    4.550432159317828e-07
+    3.007484663025798e-08
+    6.375936907597512e-08
+    1.956582100737756e-07
+    4.708254446406029e-07
+ 6.6e+10     
+    4.705723309402458e-07
+    1.956524742362015e-07
+    4.551851263962811e-07
+     6.37010195039348e-08
+    1.262215650660778e-07
+    4.551599302164799e-07
+    3.003347496967301e-08
+    6.375293115009234e-08
+    1.957487531514897e-07
+    4.709851592553703e-07
+ 6.61e+10    
+    4.707324126268118e-07
+    1.957428168562742e-07
+    4.553018972051598e-07
+     6.36942608358257e-08
+    1.262749131002295e-07
+     4.55276763579866e-07
+    2.999200151769385e-08
+    6.374637004783619e-08
+    1.958392959459001e-07
+    4.711450683513881e-07
+ 6.62e+10    
+    4.708926892760323e-07
+    1.958331584098491e-07
+    4.554187873254415e-07
+    6.368737904030366e-08
+    1.263282584336579e-07
+    4.553937160464031e-07
+    2.995042695450318e-08
+    6.373968598749377e-08
+    1.959298381256437e-07
+    4.713051719145357e-07
+ 6.63e+10    
+    4.710531608738919e-07
+    1.959234985657033e-07
+    4.555357967823773e-07
+    6.368037433971284e-08
+    1.263816012070748e-07
+    4.555107876409771e-07
+    2.990875196232169e-08
+    6.373287918932656e-08
+    1.960203793594741e-07
+    4.714654699309036e-07
+ 6.64e+10    
+    4.712138274065803e-07
+    1.960138369927415e-07
+    4.556529256016421e-07
+    6.367324695837086e-08
+    1.264349415621693e-07
+    4.556279783889009e-07
+    2.986697722537738e-08
+    6.372594987556009e-08
+    1.961109193162664e-07
+    4.716259623867972e-07
+ 6.65e+10    
+     4.71374688860493e-07
+         1.9610417336e-07
+    4.557701738093359e-07
+    6.366599712255798e-08
+    1.264882796416044e-07
+    4.557452883159151e-07
+    2.982510342987432e-08
+    6.371889827037315e-08
+    1.962014576650215e-07
+    4.717866492687356e-07
+ 6.66e+10    
+    4.715357452222318e-07
+    1.961945073366508e-07
+    4.558875414319834e-07
+    6.365862506050633e-08
+    1.265416155890153e-07
+    4.558627174481897e-07
+    2.978313126396136e-08
+    6.371172459988705e-08
+    1.962919940748703e-07
+    4.719475305634507e-07
+ 6.67e+10    
+    4.716969964786027e-07
+    1.962848385920061e-07
+    4.560050284965381e-07
+    6.365113100238909e-08
+    1.265949495490072e-07
+    4.559802658123245e-07
+    2.974106141770055e-08
+    6.370442909215481e-08
+    1.963825282150782e-07
+    4.721086062578884e-07
+ 6.68e+10    
+    4.718584426166199e-07
+    1.963751667955233e-07
+    4.561226350303811e-07
+    6.364351518030926e-08
+    1.266482816671525e-07
+    4.560979334353512e-07
+    2.969889458303539e-08
+    6.369701197715005e-08
+    1.964730597550494e-07
+     4.72269876339209e-07
+ 6.69e+10    
+     4.72020083623502e-07
+    1.964654916168083e-07
+    4.562403610613244e-07
+    6.363577782828844e-08
+    1.267016120899888e-07
+    4.562157203447331e-07
+    2.965663145375868e-08
+    6.368947348675584e-08
+     1.96563588364331e-07
+    4.724313407947847e-07
+ 6.7e+10     
+     4.72181919486675e-07
+    1.965558127256206e-07
+    4.563582066176107e-07
+    6.362791918225591e-08
+    1.267549409650166e-07
+      4.5633362656837e-07
+    2.961427272548052e-08
+    6.368181385475352e-08
+    1.966541137126176e-07
+    4.725929996122031e-07
+ 6.71e+10    
+    4.723439501937704e-07
+    1.966461297918775e-07
+    4.564761717279158e-07
+     6.36199394800366e-08
+    1.268082684406962e-07
+    4.564516521345942e-07
+    2.957181909559563e-08
+    6.367403331681113e-08
+    1.967446354697559e-07
+     4.72754852779265e-07
+ 6.72e+10    
+    4.725061757326267e-07
+    1.967364424856587e-07
+    4.565942564213496e-07
+    6.361183896133999e-08
+    1.268615946664464e-07
+    4.565697970721749e-07
+    2.952927126325091e-08
+    6.366613211047225e-08
+    1.968351533057485e-07
+    4.729169002839859e-07
+ 6.73e+10    
+    4.726685960912887e-07
+    1.968267504772099e-07
+    4.567124607274569e-07
+    6.360361786774828e-08
+    1.269149197926412e-07
+    4.566880614103205e-07
+     2.94866299293125e-08
+    6.365811047514387e-08
+    1.969256668907587e-07
+    4.730791421145947e-07
+ 6.74e+10    
+    4.728312112580073e-07
+    1.969170534369481e-07
+    4.568307846762195e-07
+    6.359527644270462e-08
+    1.269682439706078e-07
+    4.568064451786765e-07
+    2.944389579633276e-08
+    6.364996865208517e-08
+    1.970161758951146e-07
+    4.732415782595335e-07
+ 6.75e+10    
+    4.729940212212409e-07
+    1.970073510354655e-07
+    4.569492282980575e-07
+    6.358681493150122e-08
+    1.270215673526239e-07
+    4.569249484073297e-07
+     2.94010695685171e-08
+    6.364170688439532e-08
+    1.971066799893141e-07
+    4.734042087074609e-07
+ 6.76e+10    
+    4.731570259696555e-07
+    1.970976429435348e-07
+    4.570677916238303e-07
+    6.357823358126727e-08
+    1.270748900919153e-07
+    4.570435711268066e-07
+    2.935815195169058e-08
+    6.363332541700161e-08
+     1.97197178844028e-07
+    4.735670334472472e-07
+ 6.77e+10    
+    4.733202254921215e-07
+    1.971879288321114e-07
+    4.571864746848366e-07
+    6.356953264095694e-08
+    1.271282123426538e-07
+    4.571623133680788e-07
+    2.931514365326415e-08
+    6.362482449664739e-08
+    1.972876721301063e-07
+    4.737300524679794e-07
+ 6.78e+10    
+      4.7348361977772e-07
+    1.972782083723408e-07
+    4.573052775128199e-07
+    6.356071236133712e-08
+     1.27181534259954e-07
+    4.572811751625599e-07
+    2.927204538220117e-08
+    6.361620437187991e-08
+    1.973781595185807e-07
+    4.738932657589565e-07
+ 6.79e+10    
+    4.736472088157362e-07
+    1.973684812355603e-07
+    4.574242001399646e-07
+    6.355177299497483e-08
+    1.272348559998713e-07
+    4.574001565421083e-07
+    2.922885784898327e-08
+     6.36074652930379e-08
+    1.974686406806704e-07
+    4.740566733096945e-07
+ 6.8e+10     
+    4.738109925956651e-07
+    1.974587470933059e-07
+    4.575432425989011e-07
+    6.354271479622525e-08
+    1.272881777193993e-07
+    4.575192575390308e-07
+    2.918558176557636e-08
+     6.35986075122393e-08
+    1.975591152877859e-07
+    4.742202751099223e-07
+ 6.81e+10    
+     4.73974971107208e-07
+    1.975490056173146e-07
+    4.576624049227058e-07
+    6.353353802121858e-08
+    1.273414995764669e-07
+    4.576384781860791e-07
+    2.914221784539627e-08
+    6.358963128336869e-08
+    1.976495830115333e-07
+    4.743840711495838e-07
+ 6.82e+10    
+    4.741391443402745e-07
+    1.976392564795301e-07
+    4.577816871449023e-07
+    6.352424292784792e-08
+    1.273948217299367e-07
+    4.577578185164562e-07
+    2.909876680327445e-08
+    6.358053686206471e-08
+    1.977400435237195e-07
+    4.745480614188389e-07
+ 6.83e+10    
+    4.743035122849817e-07
+    1.977294993521069e-07
+    4.579010892994619e-07
+    6.351482977575609e-08
+    1.274481443396009e-07
+    4.578772785638136e-07
+    2.905522935542328e-08
+    6.357132450570714e-08
+    1.978304964963556e-07
+    4.747122459080605e-07
+ 6.84e+10    
+    4.744680749316554e-07
+     1.97819733907415e-07
+    4.580206114208086e-07
+    6.350529882632307e-08
+    1.275014675661801e-07
+    4.579968583622546e-07
+    2.901160621940155e-08
+    6.356199447340451e-08
+    1.979209416016625e-07
+    4.748766246078395e-07
+ 6.85e+10    
+    4.746328322708289e-07
+    1.979099598180437e-07
+    4.581402535438154e-07
+    6.349565034265278e-08
+      1.2755479157132e-07
+    4.581165579463349e-07
+    2.896789811407938e-08
+    6.355254702598072e-08
+    1.980113785120742e-07
+    4.750411975089785e-07
+ 6.86e+10    
+    4.747977842932446e-07
+    1.980001767568071e-07
+    4.582600157038091e-07
+    6.348588458956015e-08
+    1.276081165175889e-07
+    4.582363773510641e-07
+    2.892410575960331e-08
+    6.354298242596232e-08
+    1.981018069002433e-07
+    4.752059646024986e-07
+ 6.87e+10    
+    4.749629309898539e-07
+    1.980903843967479e-07
+    4.583798979365705e-07
+    6.347600183355805e-08
+    1.276614425684755e-07
+    4.583563166119076e-07
+    2.888022987736132e-08
+    6.353330093756534e-08
+    1.981922264390449e-07
+    4.753709258796346e-07
+ 6.88e+10    
+    4.751282723518162e-07
+     1.98180582411142e-07
+    4.584999002783361e-07
+    6.346600234284384e-08
+    1.277147698883854e-07
+    4.584763757647864e-07
+    2.883627118994736e-08
+    6.352350282668204e-08
+    1.982826368015813e-07
+    4.755360813318385e-07
+ 6.89e+10    
+    4.752938083705004e-07
+    1.982707704735031e-07
+    4.586200227657991e-07
+    6.345588638728611e-08
+     1.27768098642639e-07
+    4.585965548460787e-07
+    2.879223042112609e-08
+    6.351358836086764e-08
+    1.983730376611864e-07
+     4.75701430950777e-07
+ 6.9e+10     
+     4.75459539037485e-07
+    1.983609482575872e-07
+    4.587402654361104e-07
+    6.344565423841128e-08
+    1.278214289974689e-07
+    4.587168538926237e-07
+     2.87481082957974e-08
+    6.350355780932684e-08
+    1.984634286914303e-07
+    4.758669747283329e-07
+ 6.91e+10    
+    4.756254643445567e-07
+     1.98451115437397e-07
+    4.588606283268813e-07
+    6.343530616938998e-08
+    1.278747611200171e-07
+    4.588372729417176e-07
+    2.870390553996075e-08
+    6.349341144290055e-08
+    1.985538095661237e-07
+    4.760327126566061e-07
+ 6.92e+10    
+    4.757915842837145e-07
+    1.985412716871869e-07
+    4.589811114761838e-07
+    6.342484245502357e-08
+    1.279280951783322e-07
+    4.589578120311213e-07
+    2.865962288067953e-08
+    6.348314953405217e-08
+    1.986441799593229e-07
+    4.761986447279131e-07
+ 6.93e+10    
+    4.759578988471655e-07
+    1.986314166814668e-07
+    4.591017149225511e-07
+     6.34142633717303e-08
+    1.279814313413664e-07
+    4.590784711990558e-07
+    2.861526104604519e-08
+    6.347277235685394e-08
+    1.987345395453336e-07
+     4.76364770934786e-07
+ 6.94e+10    
+    4.761244080273272e-07
+    1.987215500950075e-07
+    4.592224387049824e-07
+    6.340356919753159e-08
+    1.280347697789739e-07
+    4.591992504842081e-07
+    2.857082076514135e-08
+    6.346228018697331e-08
+    1.988248879987157e-07
+    4.765310912699751e-07
+ 6.95e+10    
+    4.762911118168292e-07
+    1.988116716028444e-07
+     4.59343282862939e-07
+    6.339276021203821e-08
+    1.280881106619065e-07
+    4.593201499257296e-07
+    2.852630276800783e-08
+    6.345167330165899e-08
+    1.989152249942885e-07
+     4.76697605726447e-07
+ 6.96e+10    
+    4.764580102085106e-07
+    1.989017808802826e-07
+    4.594642474363499e-07
+    6.338183669643609e-08
+    1.281414541618124e-07
+    4.594411695632375e-07
+    2.848170778560449e-08
+    6.344095197972713e-08
+    1.990055502071343e-07
+    4.768643142973867e-07
+ 6.97e+10    
+    4.766251031954218e-07
+    1.989918776029015e-07
+    4.595853324656123e-07
+     6.33707989334727e-08
+    1.281948004512325e-07
+    4.595623094368186e-07
+    2.843703654977513e-08
+    6.343011650154734e-08
+    1.990958633126037e-07
+    4.770312169761957e-07
+ 6.98e+10    
+    4.767923907708254e-07
+    1.990819614465592e-07
+    4.597065379915918e-07
+    6.335964720744253e-08
+    1.282481497035979e-07
+    4.596835695870271e-07
+    2.839228979321116e-08
+    6.341916714902856e-08
+    1.991861639863196e-07
+    4.771983137564942e-07
+ 6.99e+10    
+    4.769598729281957e-07
+    1.991720320873971e-07
+    4.598278640556243e-07
+     6.33483818041731e-08
+     1.28301502093227e-07
+     4.59804950054889e-07
+    2.834746824941541e-08
+    6.340810420560505e-08
+    1.992764519041824e-07
+    4.773656046321209e-07
+ 7e+10       
+    4.771275496612187e-07
+    1.992620892018445e-07
+    4.599493106995181e-07
+    6.333700301101069e-08
+    1.283548577953231e-07
+    4.599264508819013e-07
+    2.830257265266555e-08
+    6.339692795622215e-08
+    1.993667267423742e-07
+    4.775330895971331e-07
* NOTE: Solution at 1e+08 Hz used as DC point.

.model g_m4lines_HFSS_W_1 sp N=4 SPACING=nonuniform VALTYPE=real
+ INTERPOLATION=spline
+ DATA = 700
+ 0           
+    0.0008510784137774075
+   -0.0001574885068096611
+    0.0008545778793345019
+   -1.126766962080041e-06
+   -6.750040879516493e-05
+    0.0008550095139155642
+    1.916452937783147e-07
+   -1.124233049329695e-06
+   -0.0001577728606750277
+    0.0008493537729414312
+ 2e+08       
+     0.001771925943544663
+   -0.0003422192817968613
+     0.001783399601946027
+   -1.914479231735113e-06
+   -0.0001439836006190334
+     0.001784884906339565
+   -6.883795793363981e-07
+   -1.813070534314566e-06
+   -0.0003453609017088446
+     0.001767794398634545
+ 3e+08       
+     0.002589167663714148
+   -0.0004862325620218706
+     0.002602172368458493
+    -4.24264201150778e-06
+   -0.0002051949894804335
+     0.002603649703392652
+   -1.940403693732582e-07
+   -4.204261684875072e-06
+   -0.0004883451826726586
+     0.002583267608278901
+ 4e+08       
+     0.003410105892792772
+   -0.0006320826667550488
+     0.003424593582586204
+     -5.1603471438556e-06
+   -0.0002692968407564275
+     0.003426344206001315
+    5.596352698386012e-07
+   -5.145223856449713e-06
+   -0.0006336447058186832
+     0.003402965625411628
+ 5e+08       
+     0.004251253720891197
+   -0.0007859891797900177
+     0.004268388482517638
+   -5.531784450129825e-06
+   -0.0003363604182242495
+     0.004270538996314664
+    1.186565496963342e-06
+   -5.519217064341381e-06
+   -0.0007874793443164447
+     0.004242635950122304
+ 6e+08       
+     0.005100762312396182
+   -0.0009430014308700359
+     0.005121210927044995
+   -6.066091067623449e-06
+   -0.0004039347148926231
+     0.005123776599907521
+     1.67805249550687e-06
+   -6.051272278310955e-06
+   -0.0009446545702791783
+     0.005090428624025207
+ 7e+08       
+     0.005949399036259124
+     -0.00109962973832101
+     0.005973202478298719
+   -6.900387855348104e-06
+   -0.0004708633623819473
+     0.005976190203725119
+     2.12850066081404e-06
+   -6.883330585852565e-06
+    -0.001101564261166545
+     0.005937328260258257
+ 8e+08       
+     0.006794944394096883
+    -0.001255145629963329
+     0.006821879978445718
+   -7.853925401216596e-06
+   -0.0005371624762598283
+     0.006825307379807402
+    2.624896992374523e-06
+   -7.835220263012374e-06
+    -0.001257412333507148
+     0.006781220521678108
+ 9e+08       
+     0.007639961161126815
+    -0.001410465549404944
+     0.007669958032171864
+   -8.650914985511579e-06
+   -0.0006034038777395368
+     0.007673828728046199
+    3.223908515412809e-06
+   -8.630619741544247e-06
+    -0.001413048983927965
+     0.007624599633091086
+ 1e+09       
+     0.008489164179541578
+    -0.001567089680793842
+     0.008522596763779127
+    -9.03333658169665e-06
+   -0.0006702837516171617
+     0.008526868098619748
+    3.958713626491957e-06
+   -9.010999740784024e-06
+    -0.001569901800190448
+     0.008471994312932428
+ 1.1e+09     
+     0.009370647301407945
+    -0.001727787200074973
+     0.009366855562822688
+    2.415753765599126e-05
+   -0.0007731112902522894
+     0.009372232254302549
+    7.229876557251434e-06
+    2.376656699290953e-05
+     -0.00173176563934494
+     0.009354598768759034
+ 1.2e+09     
+       0.0102481223536672
+    -0.001893792607697756
+      0.01020599011969163
+    6.175949272137525e-05
+    -0.000875200365219594
+      0.01021245539685559
+    1.123096981270121e-05
+    6.088508263419267e-05
+    -0.001898791643576986
+       0.0102330163588807
+ 1.3e+09     
+      0.01112041975081529
+    -0.002063656109322664
+      0.01104263376733386
+     0.000102874446857622
+   -0.0009764142184808645
+      0.01105015451077592
+    1.591830416995091e-05
+    0.0001014511619776099
+    -0.002069527879584429
+      0.01110601519893433
+ 1.4e+09     
+      0.01198724065482033
+    -0.002236133562164627
+      0.01187865960779419
+    0.0001466380742092825
+    -0.001076632308078522
+      0.01188718920433201
+    2.124832611136886e-05
+    0.0001446069757917355
+    -0.002242734772765423
+      0.01197325234240678
+ 1.5e+09     
+      0.01284877041680372
+    -0.002410173362987844
+       0.0127152885567882
+    0.0001922162197794848
+    -0.001175714386274561
+      0.01272477074283052
+    2.718409444819653e-05
+     0.000189526522906921
+    -0.002417370281828081
+      0.01283488768183583
+ 1.6e+09     
+      0.01370543903549413
+    -0.002584896957589115
+      0.01355323305411264
+     0.000238799400336694
+    -0.001273489455692866
+      0.01356360581311114
+    3.369837973079664e-05
+    0.0002354100497845855
+    -0.002592568877574393
+      0.01369134270144969
+ 1.7e+09     
+      0.01455777874944024
+    -0.002759577593070296
+      0.01439283330006902
+    0.0002855979113489853
+    -0.001369756259910659
+      0.01440403231369711
+    4.077453484432626e-05
+    0.0002814791063353014
+    -0.002767618967939717
+      0.01454315515444611
+ 1.8e+09     
+      0.01540634302725012
+    -0.002933619714642403
+      0.01523417073709062
+    0.0003318390314702528
+     -0.00146428875876586
+      0.01524613217673532
+    4.840584160096333e-05
+    0.0003269736955020331
+    -0.002941941186973206
+      0.01539089469079203
+ 1.9e+09     
+      0.01625166303354024
+    -0.003106540153566941
+      0.01607715625213745
+    0.0003767671564605702
+    -0.001556843576729875
+      0.01608981886985449
+    5.659372497464395e-05
+    0.0003711523147648487
+    -0.003115068697747694
+      0.01623511603388296
+ 2e+09       
+      0.01709422627890081
+    -0.003277951577255939
+      0.01692159574232088
+    0.0004196472622141386
+    -0.001647168163274186
+      0.01693490231367333
+    6.534503743878899e-05
+      0.00041329525773653
+    -0.003286629969249832
+      0.01707633471927868
+ 2.1e+09     
+        0.017934468003719
+    -0.003447548313860495
+      0.01776723725470301
+    0.0004597717879266038
+    -0.001735009211229037
+      0.01778113546804745
+    7.466852545165344e-05
+    0.0004527112396934087
+    -0.003456334116939536
+      0.01791501608618398
+ 2.2e+09     
+      0.01877276960779892
+     -0.00361509447055591
+      0.01861380390581928
+    0.0004964707752278765
+     -0.00182012120071153
+      0.01862824680396661
+    8.457057299572797e-05
+    0.0004887471627429634
+    -0.003623958696506916
+      0.01875157186372533
+ 2.3e+09     
+      0.01960946077787977
+    -0.003780414157288139
+      0.01946101619099242
+    0.0005291248554867889
+    -0.001902275013119712
+      0.01947596226565441
+    9.505035203499285e-05
+    0.0005208006031701873
+    -0.003789339730602855
+      0.01958636096790648
+ 2.4e+09     
+      0.02044482338467004
+    -0.003943383565835744
+      0.02030860656018801
+    0.0005571804274668426
+    -0.001981266517371698
+      0.02032401958631233
+    0.0001060945791401594
+    0.0005483343675715219
+    -0.003952363687952576
+      0.02041969251081226
+ 2.5e+09     
+      0.02127909606650017
+    -0.004103924618200242
+      0.02115632845519693
+    0.0005801661137402342
+    -0.002056924936184155
+      0.02117217713686957
+    0.0001176721650096375
+    0.0005708922278218902
+    -0.004112961102613369
+      0.02125182985690808
+ 2.6e+09     
+       0.0221124789137657
+     -0.00426199987972247
+      0.02200396143633198
+     0.000597709347030693
+    -0.002129120693228044
+      0.02202021892167082
+    0.0001297291323772314
+    0.0005881147264947689
+    -0.004271101508156364
+      0.02208299505917611
+ 2.7e+09     
+      0.02294513795766312
+    -0.004417608427640809
+      0.02285131358366455
+    0.0006095517506740466
+    -0.002197772349593485
+      0.02286795689467205
+    0.0001421842499831509
+    0.0005997537752510265
+    -0.004426789362900149
+      0.02291337330497939
+ 2.8e+09     
+      0.02377720933319008
+     -0.00457078237465441
+      0.02369822202398833
+    0.0006155618814485248
+    -0.002262852181293944
+       0.0237152314391224
+    0.0001549258678697207
+    0.0006056846864074526
+    -0.004580060656719502
+      0.02374311717886512
+ 2.9e+09     
+       0.0246088030798157
+    -0.004721583770159432
+      0.02454455218965197
+    0.0006157439372094871
+    -0.002324389944978919
+      0.02456191061156775
+    0.0001678104263871977
+    0.0006059143179489863
+    -0.004730979917472486
+         0.02457235065453
+ 3e+09       
+      0.02544000659245026
+    -0.004870101639710163
+      0.02539019623904384
+    0.0006102412230531088
+    -0.002382474436732029
+      0.02540788857668361
+    0.0001806630374904203
+    0.0006005841988019397
+    -0.004879637375818873
+       0.0254011727884458
+ 3.1e+09     
+      0.02627088775706725
+    -0.005016448975080827
+      0.02623507094358997
+    0.0005993335231956621
+    -0.002437252570100854
+      0.02625308353543309
+    0.0001932804003838997
+    0.0005899678380341931
+    -0.005026146100141645
+      0.02622966111933483
+ 3.2e+09     
+      0.02710149780972174
+    -0.005160759550141085
+      0.02707911525878762
+    0.0005834280179734461
+    -0.002488925874893692
+      0.02709743536150087
+     0.000205436123405843
+    0.0005744618864403509
+    -0.005170638975630282
+      0.02705787479076393
+ 3.3e+09     
+      0.02793187395161908
+    -0.005303184506419809
+      0.02792228773627153
+    0.0005630439638953425
+    -0.002537744527639932
+      0.02794090309936488
+    0.0002168883002830655
+    0.0005545713628152256
+    -0.005313265468557956
+      0.02788585741538661
+ 3.4e+09     
+      0.02876204174144964
+    -0.005443888719776785
+      0.02876456389200632
+    0.0005387919448260688
+    -0.002583999239694218
+       0.0287834624339549
+    0.0002273889600042638
+    0.0005308897110293247
+    -0.005454188182058397
+      0.02871363969394558
+ 3.5e+09     
+      0.02959201727359843
+    -0.005583047018496853
+      0.02960593361630954
+    0.0005113490206740481
+    -0.002628011518390493
+      0.02962510321102079
+    0.0002366948074895692
+    0.0005040749407248069
+    -0.005593579266444441
+      0.02954124179422391
+ 3.6e+09     
+      0.03042180914026964
+      -0.0057208403666776
+      0.03044639869008598
+    0.0004814314710642994
+    -0.002670122952154642
+      0.03046582706509364
+    0.0002445785261507861
+    0.0004748234544459207
+    -0.005731616789244769
+      0.03036867548794295
+ 3.7e+09     
+      0.03125142016917327
+    -0.005857452150574937
+      0.03128597045530561
+    0.0004497670041635077
+    -0.002710684232779521
+      0.03130564519550107
+    0.0002508398438410798
+     0.000443843329658565
+    -0.005868481193652245
+      0.03119594603935744
+ 3.8e+09     
+      0.03208084892711605
+     -0.00599306470832225
+      0.03212466767437828
+    0.0004170682582863519
+    -0.002750044610666712
+      0.03214457631835928
+    0.0002553155785089251
+    0.0004118287892091217
+     -0.00600435197780593
+      0.03202305383904495
+ 3.9e+09     
+      0.03291009098331007
+    -0.006127856227173747
+      0.03296251460151633
+    0.0003840091857600784
+    -0.002788542388809657
+      0.03298264481253196
+    0.0002578879735385142
+    0.0003794373755870335
+    -0.006139404713114591
+      0.03284999578006012
+ 4e+09       
+      0.03373913993324316
+    -0.006261998101876382
+       0.0337995392789119
+    0.0003512055242523038
+    -0.002826496916853435
+      0.03381987906939121
+    0.0002584907884046528
+    0.0003472709878147909
+    -0.006273808491994882
+      0.03367676638025664
+ 4.1e+09     
+      0.03456798819276188
+     -0.00639565280921581
+      0.03463577206147291
+    0.0003192000970873611
+    -0.002864202372440208
+      0.03465631004935348
+     0.000257112804094033
+     0.000315861506174546
+    -0.006407723859719081
+      0.03450335866269059
+ 4.2e+09     
+      0.03539662758079039
+    -0.006528972313704695
+      0.03547124436607585
+    0.0002884532102741712
+    -0.002901923439030679
+      0.03549197004236003
+    0.0002537986091883906
+    0.0002856612835236969
+    -0.006541301247568349
+      0.03532976481402256
+ 4.3e+09     
+      0.03622504971632332
+    -0.006662096983301836
+      0.03630598763495973
+    0.0002593379890172339
+     -0.00293989282954634
+      0.03632689162464086
+    0.0002486467288062902
+    0.0002570383780261807
+    -0.006674679890353532
+      0.03615597664739791
+ 4.4e+09     
+      0.03705324626004568
+    -0.006795154965781257
+      0.03714003249813722
+    0.0002321401609126223
+    -0.002978310478765105
+      0.03716110680025468
+    0.0002418053277473301
+    0.0002302760794856962
+    -0.006807987184250396
+      0.03698198590054674
+ 4.5e+09     
+      0.03788120903279924
+    -0.006928261957739682
+      0.03797340811652306
+    0.0002070615661920185
+    -0.003017344141798576
+      0.03799464631304633
+    0.0002334658509830764
+    0.0002055760594897461
+    -0.006941338422637604
+      0.03780778440149136
+ 4.6e+09     
+      0.03870893004232793
+    -0.007061521289292571
+      0.03880614168578922
+    0.0001842265575227278
+     -0.00305713109138746
+      0.03882753911280925
+    0.0002238550551798787
+    0.0001830643558258739
+    -0.007074836838411634
+      0.03863336413343417
+ 4.7e+09     
+      0.03953640144685058
+    -0.007195024246979765
+      0.03963825808051636
+    0.0001636904292030031
+    -0.003097780598045354
+      0.03965981195851498
+    0.0002132259350821488
+    0.0001627993723517717
+    -0.007208573879996992
+      0.03945871722762944
+ 4.8e+09     
+      0.04036361547975068
+    -0.007328850563244681
+      0.04046977961876796
+    0.0001454490663398669
+    -0.003139376896069437
+      0.04049148914135626
+    0.0002018480621867326
+     0.000144781117068673
+    -0.007342629653146295
+      0.04028383590896492
+ 4.9e+09     
+      0.04119056435477896
+     -0.00746306901079105
+       0.0413007259284525
+    0.0001294491046020323
+    -0.003181982375954965
+      0.04132259231088921
+    0.0001899978355143665
+    0.0001289609912765656
+    -0.007477073469540401
+      0.04110871241429088
+ 5e+09       
+      0.04201724016626384
+    -0.007597738052047176
+      0.04213111389850598
+    0.0001155980179301121
+    -0.003225640791234438
+      0.04215314038856677
+    0.0001779491011949365
+    0.0001152515602866381
+    -0.007611964454170794
+      0.04193333889880217
+ 5.1e+09     
+      0.04284363479436769
+    -0.007732906506166455
+      0.04296095769976262
+    0.0001037736868291367
+    -0.003270380318194236
+      0.04298314955425043
+    0.0001659645347358784
+    0.0001035358637162609
+    -0.007747352174886688
+      0.04275770734145107
+ 5.2e+09     
+      0.04366973982169971
+    -0.007868614207256687
+      0.04379026886223096
+    9.383313020636526e-05
+    -0.003316216355195936
+      0.04381263329271918
+    0.0001542881027908355
+    9.367594790042318e-05
+     -0.00788327726813653
+      0.04358180945670434
+ 5.3e+09     
+      0.04449554646469148
+     -0.00800489263712823
+      0.04461905639721574
+    8.562020062872946e-05
+    -0.003363153991209084
+      0.04464160248863725
+    0.0001431388354362289
+    8.552041588150931e-05
+     -0.00801977204410281
+      0.04440563661707044
+ 5.4e+09     
+      0.04532104552106383
+     -0.00814176552347912
+      0.04544732695428011
+    7.897214182798839e-05
+    -0.003411190108983237
+      0.04547006555981802
+    0.0001327060507819213
+    7.891088704028602e-05
+    -0.008156861061785448
+        0.045229179788706
+ 5.5e+09     
+      0.04614622733333946
+    -0.008279249400077742
+      0.04627508500438419
+    7.372498674901377e-05
+    -0.003460315116567516
+      0.04629802861987575
+    0.0001231460864333892
+    7.368733683640427e-05
+    -0.008294561670091606
+      0.04605242948097246
+ 5.6e+09     
+      0.04697108176755842
+    -0.008417354129361938
+       0.0471023330416913
+    6.971783487570761e-05
+    -0.003510514321936216
+      0.04712549566248853
+    0.0001145805117526717
+    6.969234745396349e-05
+     -0.00843288451480349
+      0.04687537570992557
+ 5.7e+09     
+      0.04779559820596549
+    -0.008556083390248744
+      0.04792907179752124
+    6.679609066337071e-05
+    -0.003561768980076011
+      0.04795246876049225
+    0.0001070957252059972
+    6.677434374147357e-05
+    -0.008571834013683791
+       0.0476980079752281
+ 5.8e+09     
+      0.04861976555232193
+    -0.008695435135172689
+      0.04875530046078694
+    6.481377292872972e-05
+    -0.003614057051030589
+      0.04877894827391974
+    0.0001007437854812669
+    6.478991772826317e-05
+    -0.008711408803258866
+      0.04852031524975599
+ 5.9e+09     
+      0.04944357224852374
+    -0.008835402020773365
+      0.04958101690001128
+    6.363502051690782e-05
+    -0.003667353712127925
+      0.04960493306190198
+    9.554428537580744e-05
+    6.360536148842014e-05
+    -0.008851602161291456
+      0.04934228598109217
+ 6e+09       
+       0.0502670063013072
+    -0.008975971816510508
+       0.0504062178827185
+    6.313492497288047e-05
+    -0.003721631668935767
+      0.05043042069408202
+    9.148705418725799e-05
+    6.309753457876539e-05
+    -0.008992402408887741
+      0.05016390810410531
+ 6.1e+09     
+       0.0510900553179229
+    -0.009117127795022845
+      0.05123089928863848
+    6.319981863500061e-05
+    -0.003776861308293026
+      0.05125540765787887
+    8.853546667009519e-05
+    6.315419094948707e-05
+    -0.009133793295791979
+      0.05098516906381795
+ 6.2e+09     
+      0.05191270654973563
+    -0.009258849107430989
+      0.05205505631377821
+    6.372713865775571e-05
+    -0.003833010733814739
+      0.05207988955857452
+    8.663014264164728e-05
+    6.367388318426637e-05
+    -0.009275754371868224
+      0.05180605584776968
+ 6.3e+09     
+      0.05273494694275353
+    -0.009401111146131179
+      0.05287868366299585
+    6.462497581506877e-05
+    -0.003890045720199682
+      0.05290386130980098
+    8.569283835998642e-05
+    6.456555100581036e-05
+    -0.009418261347163693
+      0.05262655502705021
+ 6.4e+09     
+      0.05355676319409816
+    -0.009543885897001711
+      0.05370177572926522
+    6.581140309774083e-05
+    -0.003947929617986348
+      0.05372731731255915
+    8.563035578198347e-05
+    6.574788774400798e-05
+    -0.009561286442364276
+       0.0534466528051305
+ 6.5e+09     
+      0.05437814181342004
+    -0.009687142282390001
+      0.05452432675833167
+    6.721366437450208e-05
+    -0.004006623235495338
+      0.05455025162142136
+    8.633832562624996e-05
+    6.714856419612553e-05
+    -0.009704798730925612
+      0.05426633507355241
+ 6.6e+09     
+      0.05519906918824027
+    -0.009830846495776605
+      0.05534633099793359
+    6.876728873568723e-05
+    -0.004066084719853167
+      0.05537265809703259
+    8.770475194403186e-05
+    6.870337502009011e-05
+    -0.009848764473712345
+      0.05508558747347625
+ 6.7e+09     
+      0.05601953165218612
+    -0.009974962328626234
+        0.056167782831184
+    7.041518230312994e-05
+    -0.004126269454412951
+      0.05619453054443917
+    8.961323722684656e-05
+    7.035535923423592e-05
+    -0.009993147446603769
+      0.05590439546202857
+ 6.8e+09     
+       0.0568395155550816
+     -0.01011945148962717
+      0.05698867689408103
+    7.210673675857906e-05
+    -0.004187129985704166
+      0.05701586283713177
+    9.194583610480449e-05
+    7.205393406222371e-05
+      -0.0101379092612206
+      0.05672274438235515
+ 6.9e+09     
+      0.05765900733386645
+      -0.0102642739162764
+      0.05780900817742445
+    7.379698290149749e-05
+    -0.004248615989324207
+      0.05783664902698821
+    9.458551115924026e-05
+    7.375407054915906e-05
+     -0.01028300967868806
+      0.05754061953627353
+ 7e+09       
+      0.05847799358335177
+     -0.01040938807858097
+      0.05862877211367738
+    7.544580830715802e-05
+    -0.004310674280960753
+      0.05865688344054391
+    9.741818558776797e-05
+    7.541553022204781e-05
+       -0.010428406916161
+      0.05835800625842737
+ 7.1e+09     
+       0.0592964611258734
+     -0.01055475127450419
+       0.0594479646495128
+    7.701725060223474e-05
+    -0.004373248875996881
+      0.05947656076220834
+    0.0001003344041908337
+    7.700217456310969e-05
+     -0.01057405794569343
+      0.05917488999088438
+ 7.2e+09     
+      0.06011439707897451
+     -0.01070031991668015
+      0.06026658230493551
+    7.847887190992793e-05
+    -0.004436281098878922
+      0.06029567610518223
+    0.0001032306265293049
+    7.848135312272944e-05
+     -0.01071991878492601
+      0.05999125635717729
+ 7.3e+09     
+      0.06093178892033792
+     -0.01084604980984734
+      0.06108462221997773
+    7.980121546523702e-05
+    -0.004499709741575255
+        0.061114225070927
+    0.0001060101845270528
+    7.982337155420681e-05
+     -0.01086594477898825
+      0.06080709123486273
+ 7.4e+09     
+      0.06174862454928029
+      -0.0109918964184047
+      0.06190208219002505
+    8.095734208441851e-05
+    -0.004563471268980868
+      0.06193220379808818
+    0.0001085839417994975
+    8.100103752655763e-05
+     -0.01101209087296138
+      0.06162238082576305
+ 7.5e+09     
+      0.06256489234422634
+     -0.01113781512346969
+      0.06271896069086078
+    8.192244187231348e-05
+    -0.004627500067975601
+      0.06274960900180149
+    0.0001108706941945696
+     8.19892801584678e-05
+     -0.01115831187422128
+       0.0624371117231544
+ 7.6e+09     
+      0.06338058121568364
+     -0.01128376146881551
+      0.06353525689451184
+    8.267351508627426e-05
+    -0.004691728735980428
+      0.06356643800429919
+    0.0001127973510503745
+    8.276483712903009e-05
+      -0.0113045627039751
+      0.06325127097526799
+ 7.7e+09     
+      0.06419568065433982
+      -0.0114296913950779
+      0.06435097067695381
+    8.318911525155348e-05
+    -0.004756088404229038
+      0.06438268875771128
+    0.0001142989350789261
+    8.330600277655503e-05
+     -0.01145079863731865
+      0.06406484614457277
+ 7.8e+09     
+      0.06501018077400746
+     -0.01157556146165467
+      0.06516610261868466
+    8.344914729401767e-05
+    -0.004820509090547046
+      0.06519835985990741
+    0.0001153184360835669
+    8.359243014300667e-05
+     -0.01159697553117163
+       0.0648778253624134
+ 7.9e+09     
+      0.06582407234922885
+     -0.01172132905576496
+      0.06598065399911926
+    8.343471348116799e-05
+    -0.004884920076173317
+      0.06601345056417604
+    0.0001158065503320826
+    8.360497992468147e-05
+     -0.01174305003949484
+      0.06569019737867086
+ 8e+09       
+      0.06663734684744317
+     -0.01186695258819349
+      0.06679462678568493
+    8.312800023565245e-05
+    -0.004949250301039584
+       0.0668279607834657
+    0.0001157213336786256
+    8.332560954163546e-05
+     -0.01188897981525035
+      0.06650195160620648
+ 8.1e+09     
+      0.06744999645569237
+     -0.01201239167531202
+      0.06760802361842037
+     8.25121993204586e-05
+    -0.005013428771922453
+      0.06764189108985301
+     0.000115027792712279
+    8.273729595293603e-05
+     -0.01203472369863665
+      0.06731307815993343
+ 8.2e+09     
+      0.06826201410191134
+     -0.01215760730704517
+      0.06842084779080335
+    8.157145742544378e-05
+    -0.005077384977976215
+      0.06845524270982713
+    0.0001136974344979136
+    8.182398635645525e-05
+     -0.01218024189120881
+      0.06812356789043654
+ 8.3e+09     
+      0.06907339347090806
+     -0.01230256200053086
+       0.0692331032274504
+    8.029084876124646e-05
+    -0.005141049308330561
+      0.06926801751591356
+    0.0001117077919918818
+    8.057057147326354e-05
+     -0.01232549611557793
+      0.06893341241212894
+ 8.4e+09     
+      0.06988412901518755
+     -0.01244721993930725
+      0.07004479445925176
+    7.865636585167033e-05
+    -0.005204353466677565
+      0.07008021801509449
+    0.0001090419390415642
+    7.896287668804043e-05
+     -0.01247044976047426
+      0.06974260412599376
+ 8.5e+09     
+      0.07069421596081966
+      -0.0125915470979489
+       0.0708559265964316
+     7.66549242925983e-05
+    -0.005267230878068749
+      0.07089184733441832
+    0.0001056880060519979
+    7.698766687888733e-05
+     -0.01261506801104872
+      0.07055113623701272
+ 8.6e+09     
+       0.0715036503085807
+     -0.01273551135215817
+      0.07166650529994989
+    7.427437778823368e-05
+    -0.005329617083483782
+      0.07170290920413744
+    0.0001016387049398669
+    7.463266130347708e-05
+     -0.01275931796438039
+      0.07135900276642708
+ 8.7e+09     
+      0.07231242883063195
+     -0.01287908257440613
+      0.07247653675159808
+    7.150354028241846e-05
+    -0.005391450118106862
+      0.07251340793865671
+    9.689086988599795e-05
+    7.188655540747539e-05
+      -0.0129031687302474
+      0.07216619855901459
+ 8.8e+09     
+      0.07312054906301364
+     -0.01302223271529755
+      0.07328602762308116
+    6.833221246805205e-05
+    -0.005452670869650163
+      0.07332334841553549
+    9.144501862217618e-05
+    6.873904687468377e-05
+     -0.01304659151730643
+      0.07297271928559784
+ 8.9e+09     
+      0.07392800929425257
+     -0.01316493587091456
+      0.07409498504432396
+    6.475121037745866e-05
+    -0.005513223413485311
+      0.07413273605274134
+    8.530493751705381e-05
+    6.518086365615936e-05
+     -0.01318955970490946
+      0.07377856144102299
+ 9e+09       
+      0.07473480855038991
+     -0.01330716833646556
+      0.07490341657119427
+    6.075239413307645e-05
+    -0.005573055321776948
+       0.0749415767843235
+    7.847729252804343e-05
+    6.120379208253684e-05
+     -0.01333204890086552
+      0.07458372233787186
+ 9.1e+09     
+      0.07554094657674133
+     -0.01344890864663447
+      0.07571133015279748
+    5.632869527549312e-05
+    -0.005632117944253744
+      0.07574987703464645
+    7.097126712418277e-05
+    5.680070349855853e-05
+     -0.01347403698552648
+      0.07538820009617954
+ 9.2e+09     
+      0.07634642381670319
+     -0.01359013760308577
+      0.07651873409845922
+    5.147414138236781e-05
+    -0.005690366658689767
+      0.07655764369130259
+    6.279822752981896e-05
+    5.196557815042181e-05
+     -0.01361550414264266
+      0.07619199362944658
+ 9.3e+09     
+       0.0771512413879175
+     -0.01373083828963498
+      0.07732563704448983
+    4.618387695498437e-05
+    -0.005747761089603521
+      0.07736488407680467
+    5.397141505449239e-05
+    4.669352531928763e-05
+     -0.01375643287749264
+      0.07699510262723606
+ 9.4e+09     
+      0.07795540105610359
+     -0.01387099607564256
+      0.07813204792080115
+    4.045417978145539e-05
+    -0.005804265294103847
+      0.07817160591915054
+    4.450566483696307e-05
+    4.098079891801717e-05
+     -0.01389680802284254
+      0.07779752753465401
+ 9.5e+09     
+      0.07875890520685526
+     -0.01401059860822818
+      0.07893797591742954
+    3.428247218671633e-05
+    -0.005859847914218273
+      0.07897781732134339
+    3.441715001023071e-05
+    3.482480797379565e-05
+      -0.0140366167333357
+      0.07859926952900834
+ 9.6e+09     
+      0.07956175681569662
+      -0.0141496357939363
+      0.07974343045100651
+    2.766732675806341e-05
+    -0.005914482295426426
+      0.07978352672994329
+    2.372315007245123e-05
+    2.822412159033272e-05
+     -0.01417584846894824
+      0.07940033049394091
+ 9.7e+09     
+       0.0803639594166758
+     -0.01428809977051075
+      0.08054842113121496
+    2.060846628590282e-05
+    -0.005968146571484841
+      0.08058874290273435
+    1.244184210267207e-05
+    2.117846813792052e-05
+     -0.01431449496817849
+      0.08020071299132328
+ 9.8e+09     
+       0.0811655170697643
+     -0.01442598486945463
+      0.08135295772725755
+    1.310675779785906e-05
+    -0.006020823715967715
+      0.08139347487558041
+    5.921133757447704e-07
+    1.368872855113954e-05
+     -0.01445255021165742
+      0.08100042023119734
+ 9.9e+09     
+      0.08196643432731809
+      -0.0145632875700674
+      0.08215705013437155
+    5.164200672465183e-06
+    -0.006072501561257212
+      0.08219773192855788
+    -1.18066061048209e-05
+    5.756923727087433e-06
+     -0.01459001037688715
+       0.0817994560400383
+ 1e+10       
+      0.08276671619984004
+      -0.0147000064456568
+      0.08296070834041837
+   -3.216091076274673e-06
+    -0.006123172785997904
+      0.08300152355145053
+   -2.473449263825115e-05
+   -2.613803885043002e-06
+     -0.01472687378482095
+      0.08259782482760331
+ 1.01e+10    
+      0.08356636812127072
+     -0.01483614210262676
+      0.08376394239258232
+   -1.202991217560826e-05
+    -0.006172834872278019
+      0.08380485940870015
+   -3.817146087677862e-05
+   -1.141921432833582e-05
+     -0.01486314083900426
+      0.08339553155262137
+ 1.02e+10    
+      0.08436539591401813
+      -0.0149716971131393
+      0.08456676236421933
+   -2.127199488717059e-05
+      -0.0062214900340186
+      0.08460774930391393
+     -5.2097280302448e-05
+   -2.065399957644704e-05
+     -0.01499881395799409
+      0.08419258168756835
+ 1.03e+10    
+      0.08516380575392428
+     -0.01510667594204081
+      0.08536917832189828
+   -3.093604292283127e-05
+    -0.006269145118237253
+      0.08541020314403223
+   -6.649167747689025e-05
+   -3.031181806401268e-05
+     -0.01513389750176769
+      0.08498898118275607
+ 1.04e+10    
+      0.08596160413534769
+     -0.01524108486873209
+      0.08617120029268674
+    -4.10147701332133e-05
+    -0.006315811481009369
+      0.08621223090327078
+   -8.133442534183355e-05
+   -4.038533396398276e-05
+     -0.01526839769282052
+      0.08578473642995479
+ 1.05e+10    
+      0.08675879783653023
+     -0.01537493190464557
+      0.08697283823173804
+   -5.149994359075717e-05
+     -0.00636150484007285
+      0.08701384258695402
+   -9.660542077062238e-05
+   -5.086626082989815e-05
+     -0.01540232253263983
+      0.08657985422575426
+ 1.06e+10    
+      0.08755539388539914
+     -0.01550822670697573
+      0.08777410199024283
+   -6.238243065468069e-05
+    -0.006406245106120183
+      0.08781504819536058
+   -0.0001122847514951038
+    -6.17454091918811e-05
+     -0.01553568171421985
+      0.08737434173485299
+ 1.07e+10    
+      0.08835139952594125
+     -0.01564098048928602
+      0.08857500128381464
+   -7.365224959117933e-05
+    -0.006450056194887402
+      0.08861585768771089
+   -0.0001283527534515364
+   -7.301273767832848e-05
+       -0.015668486531266
+      0.08816820645345637
+ 1.08e+10    
+      0.08914682218527498
+     -0.01577320592959388
+      0.08937554566138387
+   -8.529862330254861e-05
+    -0.006492965822193944
+      0.08941628094642218
+   -0.0001447900595138991
+   -8.465740721888245e-05
+     -0.01580074978470856
+      0.08896145617294483
+ 1.09e+10    
+      0.08994166944152722
+     -0.01590491707650735
+      0.09017574447468016
+   -9.731003572090505e-05
+    -0.006535005284102367
+      0.09021632774176515
+   -0.0001615776405052144
+    -9.66678378825094e-05
+     -0.01593248568712341
+      0.08975409894396683
+ 1.1e+10     
+      0.09073594899261667
+     -0.01603612925396251
+      0.09097560684838657
+   -0.0001096742904123267
+    -0.006576209224365417
+      0.09101600769705509
+   -0.0001786968393079364
+   -0.0001090317678995117
+      -0.0160637097656268
+      0.09054614304109207
+ 1.11e+10    
+      0.09152966862602482
+     -0.01616685896507901
+      0.09177514165104972
+   -0.0001223785709509675
+     -0.00661661539129986
+      0.09181533025450685
+   -0.0001961293988232836
+   -0.0001217363144236012
+     -0.01619443876378364
+      0.09133759692815213
+ 1.12e+10    
+       0.0923228361896303
+     -0.01629712379562464
+      0.09257435746683719
+   -0.0001354095026218827
+    -0.006656264386186705
+      0.09261430464188658
+   -0.0002138574844665385
+   -0.0001347680355987648
+      -0.0163246905430377
+      0.09212846922437994
+ 1.13e+10    
+      0.09311545956366984
+     -0.01642694231754747
+      0.09337326256822823
+   -0.0001487532150327952
+    -0.006695199405236592
+      0.09341293984008875
+    -0.000231863701823196
+   -0.0001481129935056676
+     -0.01645448398414147
+      0.09291876867145106
+ 1.14e+10    
+      0.09390754663387586
+     -0.01655633399300463
+      0.09417186488972819
+   -0.0001623954052219034
+    -0.006733465977087122
+      0.09421124455176014
+   -0.0002501311100352051
+   -0.0001617568175810852
+     -0.01658383888903095
+      0.09370850410151314
+ 1.15e+10    
+      0.09469910526583512
+     -0.01668531907928595
+      0.09497017200269441
+   -0.0001763214008741659
+    -0.006771111697714323
+      0.09500922717109336
+   -0.0002686432314332739
+   -0.0001756847681187194
+     -0.01671277588356056
+      0.09449768440628491
+ 1.16e+10    
+      0.09549014328060032
+     -0.01681391853499905
+      0.09576819109135679
+    -0.000190516223274063
+    -0.006808185964544873
+      0.09580689575490244
+   -0.0002873840578824713
+   -0.0001898817994844299
+      -0.0168413163214798
+      0.09528631850729022
+ 1.17e+10    
+      0.09628066843158137
+     -0.01694215392785432
+      0.09656592893011871
+   -0.0002049646496485181
+    -0.006844739711454147
+      0.09660425799508945
+   -0.0003063380542635721
+   -0.0002043326226962442
+      -0.0169694821900029
+      0.09607441532728433
+ 1.18e+10    
+      0.09707068838273163
+     -0.01707004734435537
+      0.09736339186221456
+   -0.0002196512745735357
+     -0.00688082514622465
+      0.09740132119260075
+   -0.0003254901594712018
+   -0.0002190217670476717
+     -0.01709729601729171
+      0.09686198376292279
+ 1.19e+10    
+      0.09786021068803968
+     -0.01719762130167354
+      0.09816058577979656
+    -0.000234560570145862
+    -0.006916495491926243
+      0.09819809223296681
+    -0.000344825785271854
+    -0.000233933640472494
+     -0.01722478078214099
+      0.09764903265870831
+ 1.2e+10     
+      0.09864924277233009
+     -0.01732489866195541
+      0.09895751610552199
+   -0.0002496769446452246
+    -0.006951804733561326
+      0.09899457756350986
+   -0.0003643308133289501
+   -0.0002490525883811134
+     -0.01735195982612576
+      0.09843557078224896
+ 1.21e+10    
+      0.09943779191336999
+     -0.01745190254928416
+       0.0997541877756999
+   -0.0002649847994362088
+    -0.006986807371199782
+      0.09979078317229231
+   -0.0003839915906723181
+   -0.0002643629507157142
+     -0.01747885676844187
+      0.09922160680084782
+ 1.22e+10    
+       0.1002258652252732
+     -0.01757865626949005
+       0.1005506052250536
+   -0.0002804685838884326
+    -0.007021558180707656
+       0.1005867145688736
+   -0.0004037949238575966
+   -0.0002798491170047804
+     -0.01760549542364289
+       0.1000071492594407
+ 1.23e+10    
+        0.101013469643188
+     -0.01770518323297723
+       0.1013467723731456
+   -0.0002961128481146582
+    -0.007056111983054045
+       0.1013823767669306
+   -0.0004237280720369033
+   -0.0002954955792187465
+      -0.0177318997224487
+        0.100792206559889
+ 1.24e+10    
+       0.1018006119092505
+     -0.01783150688071203
+       0.1021426926125089
+   -0.0003119022933556529
+    -0.007090523423063029
+       0.1021777742687864
+   -0.0004437787391359982
+   -0.0003112869822540628
+     -0.01785809363577685
+       0.1015767869416297
+ 1.25e+10    
+       0.1025872985597828
+     -0.01795765061349141
+       0.1029383687985106
+   -0.0003278218198632054
+    -0.007124846758360549
+       0.1029729110518862
+    -0.000463935065311733
+   -0.0003272081718997226
+     -0.01798410110212233
+       0.1023608984636773
+ 1.26e+10    
+       0.1033735359137084
+     -0.01808363772459042
+       0.1037338032409788
+   -0.0003438565721556616
+    -0.007159135659154109
+       0.1037677905572425
+   -0.0004841856178440834
+   -0.0003432442401612532
+     -0.01810994595838733
+       0.1031445489879703
+ 1.27e+10    
+       0.1041593300621564
+     -0.01820949133586375
+       0.1045289976976039
+   -0.0003599919815467365
+    -0.007193443019373167
+       0.1045624156798685
+   -0.0005045193815970714
+   -0.0003593805678434748
+     -0.01823565187424241
+       0.1039277461640448
+ 1.28e+10    
+       0.1049446868592248
+     -0.01833523433735792
+       0.1053239533691245
+   -0.0003762138058671154
+    -0.007227820779593416
+       0.1053567887612048
+   -0.0005249257491681597
+   -0.0003756028643134351
+     -0.01836124229007711
+       0.1047104974150185
+ 1.29e+10    
+       0.1057296119138652
+     -0.01846088933047181
+       0.1061186708962955
+   -0.0003925081663217748
+    -0.007262319762068348
+       0.1061509115835352
+   -0.0005453945108296219
+   -0.0003918972043843293
+     -0.01848674035858078
+       0.1054928099248606
+ 1.3e+10     
+       0.1065141105828562
+     -0.01858647857468382
+       0.1069131503586319
+   -0.0004088615814446337
+    -0.007296989518094762
+       0.1069447853663791
+   -0.0005659158443514643
+   -0.0004082500622881111
+     -0.01861216888997393
+       0.1062746906269204
+ 1.31e+10    
+       0.1072981879648236
+     -0.01871202393784969
+       0.1077073912749077
+   -0.0004252609981321694
+    -0.007331878187850858
+       0.1077384107648386
+   -0.0005864803047842164
+   -0.0004246483427143089
+     -0.01873755030089477
+       0.1070561461936869
+ 1.32e+10    
+       0.1080818488952731
+     -0.01883754685005834
+       0.1085013926053894
+   -0.0004416938197553367
+    -0.007367032372759826
+       0.1085317878698692
+    -0.000607078814267806
+   -0.0004410794089169112
+     -0.01886290656692965
+       0.1078371830277439
+ 1.33e+10    
+       0.1088650979425892
+     -0.01896306826101932
+       0.1092951527557688
+     -0.00045814793136342
+    -0.007402497020354373
+       0.1093249162104356
+   -0.0006277026519232311
+   -0.0004575311079056156
+     -0.01898825917876003
+       0.1086178072538868
+ 1.34e+10    
+        0.109647939404963
+     -0.01908860860094248
+       0.1100886695827581
+   -0.0004746117220118777
+    -0.007438315321544499
+       0.1101177947575047
+   -0.0006483434438744884
+   -0.0004739917927513299
+     -0.01911362910188691
+       0.1093980247123619
+ 1.35e+10    
+       0.1104303773082043
+     -0.01921418774485843
+       0.1108819404012977
+   -0.0004910741042585021
+    -0.007474528620123786
+       0.1109104219298229
+   -0.0006689931534402884
+    -0.000490450342052794
+     -0.01923903673988107
+       0.1101778409531926
+ 1.36e+10    
+       0.1112124154043962
+     -0.01933982498031852
+       0.1116749619933291
+   -0.0005075245308841523
+    -0.007511176334290182
+       0.1117027956014165
+   -0.0006896440715277075
+   -0.0005068961766205894
+     -0.01936450190109448
+       0.1109572612315463
+ 1.37e+10    
+       0.1119940571713494
+     -0.01946553897840203
+       0.1124677306180706
+   -0.0005239530089071158
+    -0.007548295889900515
+       0.1124949131107485
+   -0.0007102888072534445
+   -0.0005233192734497259
+     -0.01949004376876144
+       0.1117362905041034
+ 1.38e+10    
+       0.1127753058128122
+     -0.01959134776795015
+       0.1132602420237332
+   -0.0005403501109712968
+    -0.007585922665129837
+       0.1132867712714575
+   -0.0007309202788127146
+   -0.0005397101770584275
+     -0.01961568087440576
+        0.112514933426385
+ 1.39e+10    
+       0.1135561642593942
+     -0.01971726871293968
+         0.11405249146061
+   -0.0005567069841930968
+    -0.007624089946163619
+       0.1140783663846046
+   -0.0007515317046106551
+   -0.0005560600082831577
+     -0.01974143107446483
+       0.1132931943509938
+ 1.4e+10     
+       0.1143366351701606
+     -0.01984331849290034
+       0.1148444736954627
+   -0.0005730153565664871
+    -0.007662828893511867
+       0.1148696942523427
+    -0.000772116594666473
+   -0.0005723604706256678
+     -0.01986731153003281
+       0.1140710773267251
+ 1.41e+10    
+       0.1151167209348552
+     -0.01996951308627642
+       0.1156361830271323
+   -0.0005892675410249825
+    -0.007702168518502887
+       0.1156607501929255
+   -0.0007926687422969252
+   -0.0005886038542545361
+     -0.01999333868962028
+       0.1148485860985022
+ 1.42e+10    
+       0.1158964236767096
+     -0.02009586775662591
+       0.1164276133032898
+   -0.0006054564372723219
+     -0.00774213566948549
+       0.1164515290569641
+    -0.000813182216081849
+   -0.0006047830377711528
+     -0.02011952827482135
+       0.1156257241080927
+ 1.43e+10    
+        0.116675745255799
+     -0.02022239704154857
+       0.1172187579382504
+   -0.0006215755314910396
+    -0.007782755027247889
+        0.117242025244845
+    -0.000833651352111634
+   -0.0006208914878528676
+     -0.02024589526877639
+       0.1164024944955592
+ 1.44e+10    
+       0.1174546872729024
+     -0.02034911474422853
+       0.1180096099317588
+   -0.0006376188940482779
+    -0.007824049109141761
+       0.1180322327252092
+   -0.0008540707465144385
+   -0.0006369232568893051
+     -0.02037245390731344
+       0.1171789001014015
+ 1.45e+10    
+       0.1182332510738287
+     -0.02047603392747638
+       0.1188001618886657
+   -0.0006535811753163457
+    -0.007866038281388031
+       0.1188221450544043
+   -0.0008744352482573988
+    -0.000652872978733351
+     -0.02049921767264989
+       0.1179549434693443
+ 1.46e+10    
+       0.1190114377541712
+     -0.02060316691015252
+        0.119590406039405
+   -0.0006694575997288487
+     -0.00790874077903116
+       0.1196117553968096
+    -0.000894739952216163
+   -0.0006687358626857355
+     -0.02062619928953326
+       0.1187306268497304
+ 1.47e+10    
+        0.119789248164451
+     -0.02073052526585273
+       0.1203803342611846
+   -0.0006852439581952534
+     -0.00795217273300344
+       0.1204010565459397
+   -0.0009149801925034773
+    -0.000684507685837909
+     -0.02075341072369834
+       0.1195059522034706
+ 1.48e+10    
+       0.1205666829156136
+     -0.02085811982373524
+        0.121169938099802
+   -0.0007009365989947996
+    -0.007996348203759602
+       0.1211900409462335
+    -0.000935151536047979
+    -0.000700184783893866
+     -0.02088086318251828
+       0.1202809212065145
+ 1.49e+10    
+       0.1213437423848441
+     -0.02098596067136988
+       0.1219592087919982
+   -0.0007165324172718141
+    -0.008041279220943101
+       0.1219787007154279
+   -0.0009552497764123962
+   -0.0007157640405936194
+     -0.02100856711772519
+        0.121055535254797
+ 1.5e+10     
+       0.1221204267216667
+     -0.02111405715948893
+        0.122748137288262
+   -0.0007320288432537522
+     -0.00808697582855104
+       0.1227670276674285
+   -0.0009752709278397992
+   -0.0007312428758588473
+     -0.02113653223007787
+        0.121829795469621
+ 1.51e+10    
+       0.1228967358542938
+     -0.02124241790852026
+       0.1235367142760004
+   -0.0007474238293091531
+    -0.008133446135071845
+       0.1235550133355822
+   -0.0009952112195160132
+   -0.0007466192327805054
+     -0.02126476747585394
+       0.1226037027034375
+ 1.52e+10    
+       0.1236726694961947
+     -0.02137105081678477
+       0.1243249302029902
+    -0.000762715835962096
+    -0.008180696368080515
+       0.1243426489962612
+    -0.001015067090036255
+    -0.000761891563563993
+     -0.02139328107504553
+       0.1233772575459862
+ 1.53e+10    
+       0.1244482271528542
+     -0.02149996307024201
+       0.1251127753010285
+   -0.0007779038169785201
+    -0.008228730932787637
+        0.125129925692672
+    -0.001034835182063112
+   -0.0007770588145462071
+     -0.02152208052113876
+       0.1241504603307563
+ 1.54e+10    
+       0.1252234081286887
+     -0.02162916115366889
+       0.1259002396097057
+   -0.0007929872036331843
+    -0.008277552474054393
+       0.1259168342588038
+    -0.001054512337163541
+   -0.0007921204103958869
+     -0.02165117259235944
+       0.1249233111417347
+ 1.55e+10    
+       0.1259982115340958
+     -0.02175865086315931
+       0.1266873130002172
+   -0.0008079658882644951
+    -0.008327161941400601
+       0.1267033653434329
+    -0.001074095590812432
+   -0.0008070762376036003
+     -0.02178056336427015
+       0.1256958098204077
+ 1.56e+10    
+       0.1267726362926079
+     -0.02188843731983514
+       0.1274739851991491
+   -0.0008228402072213274
+    -0.008377558656551423
+       0.1274895094341068
+    -0.001093582167550355
+   -0.0008219266273648473
+     -0.02191025822360606
+       0.1264679559729799
+ 1.57e+10    
+       0.1275466811481257
+     -0.02201852498466136
+       0.1282602458121583
+   -0.0008376109232986769
+    -0.008428740383087054
+       0.1282752568810293
+    -0.001112969476283732
+   -0.0008366723379556375
+     -0.02204026188323942
+       0.1272397489777817
+ 1.58e+10    
+       0.1283203446722075
+     -0.02214891767426087
+       0.1290460843474843
+   -0.0008522792077595985
+    -0.008480703397779257
+       0.1290605979207764
+    -0.001132255105715274
+   -0.0008513145366953077
+     -0.02217057839816623
+        0.128011187992834
+ 1.59e+10    
+       0.1290936252713925
+     -0.02227961857762933
+       0.1298314902392262
+   -0.0008668466220307942
+    -0.008533442563220771
+       0.1298455226997768
+    -0.001151436819893943
+   -0.0008658547815862299
+     -0.02230121118241248
+       0.1287822719635394
+ 1.6e+10     
+       0.1298665211945332
+     -0.02241063027365092
+       0.1306164528703257
+   -0.0008813150991584147
+    -0.008586951401373406
+       0.1306300212974858
+    -0.001170512553873492
+   -0.0008802950027165125
+     -0.02243216302675866
+       0.1295529996304763
+ 1.61e+10    
+       0.1306390305401232
+     -0.02254195474932262
+       0.1314009615951968
+   -0.0008956869251052608
+    -0.008641222167683905
+       0.1314140837492022
+    -0.001189480409469147
+   -0.0008946374835056463
+     -0.02256343611718773
+       0.1303233695372649
+ 1.62e+10    
+       0.1314111512635937
+     -0.02267359341859521
+       0.1321850057619512
+   -0.0009099647199636608
+     -0.00869624592543799
+       0.1321977000684638
+    -0.001208338651103084
+   -0.0009088848418702389
+     -0.02269503205396314
+       0.1310933800384848
+ 1.63e+10    
+       0.1321828811845679
+     -0.02280554714174507
+       0.1329685747341679
+   -0.0009241514191551614
+    -0.008752012620045669
+       0.1329808602689709
+    -0.001227085701729623
+   -0.0009230400113789229
+     -0.02282695187124777
+       0.1318630293076156
+ 1.64e+10    
+       0.1329542179940524
+     -0.02293781624519396
+       0.1337516579121629
+   -0.0009382502546852697
+    -0.008808511152973188
+        0.133763554385995
+    -0.001245720138831079
+   -0.0009371062224644228
+     -0.02295919605718017
+       0.1326323153449856
+ 1.65e+10    
+       0.1337251592615522
+      -0.0230704005416962
+       0.1345342447537145
+   -0.0009522647365106733
+    -0.008865729455058353
+       0.1345457724972204
+    -0.001264240690477461
+   -0.0009510869837519951
+      -0.0230917645743256
+       0.1334012359856984
+ 1.66e+10    
+       0.1344957024420952
+      -0.0232032993508197
+       0.1353163247942088
+   -0.0009661986340786823
+    -0.008923654558968337
+       0.1353275047429845
+    -0.001282646231441638
+   -0.0009649860635635226
+     -0.02322465688042535
+       0.1341697889075285
+ 1.67e+10    
+       0.1352658448831514
+     -0.02333651151964757
+       0.1360978876661685
+   -0.0009800559580889149
+    -0.008982272670580532
+       0.1361087413458796
+    -0.001300935779364394
+   -0.0009788074716452592
+     -0.02335787194937157
+       0.1349379716387578
+ 1.68e+10    
+       0.1360355838314391
+     -0.02347003544363401
+       0.1368789231181351
+   -0.0009938409425247897
+    -0.009041569239086736
+       0.1368894726296812
+    -0.001319108490962697
+   -0.0009925554411702227
+     -0.02349140829233733
+       0.1357057815659441
+ 1.69e+10    
+       0.1368049164396009
+     -0.02360386908754864
+       0.1376594210328765
+     -0.00100755802699764
+    -0.009101529025641968
+       0.1376696890375777
+    -0.001337163658276054
+    -0.001006234411055425
+     -0.02362526397899712
+       0.1364732159416009
+ 1.7e+10     
+       0.1375738397727462
+     -0.02373801000645081
+       0.1384393714448971
+    -0.001021211839442131
+    -0.009162136170398828
+       0.1384493811496748
+    -0.001355100704946221
+    -0.001019849008633749
+     -0.02375943665877629
+       0.1372402718917763
+ 1.71e+10    
+       0.1383423508148459
+     -0.02387245536663606
+       0.1392187645572279
+    -0.001034807179196651
+    -0.009223374257786609
+       0.1392285396997548
+    -0.001372919182526088
+    -0.001033404032713106
+     -0.02389392358207117
+       0.1380069464235174
+ 1.72e+10    
+        0.139110446474976
+     -0.02400720196650224
+       0.1399975907574806
+    -0.001048349000499203
+    -0.009285226379912094
+       0.1400071555912695
+     -0.00139061876681389
+    -0.001046904437055379
+     -0.02402872162138618
+       0.1387732364322082
+ 1.73e+10    
+       0.1398781235933997
+     -0.02414224625728549
+       0.1407758406331506
+    -0.001061842396425864
+    -0.009347675197976968
+       0.1407852199125581
+    -0.001408199254209726
+    -0.001060355314299597
+     -0.02416382729233744
+       0.1395391387087701
+ 1.74e+10    
+       0.1406453789474825
+      -0.0242775843636209
+       0.1415535049861597
+    -0.001075292583293325
+    -0.009410703001622566
+       0.1415627239512716
+    -0.001425660558091913
+    -0.001073761880352987
+     -0.02429923677447551
+       0.1403046499467135
+ 1.75e+10    
+       0.1414122092574375
+     -0.02441321210388385
+       0.1423305748466235
+     -0.00108870488554596
+    -0.009474291766127779
+       0.1423396592080033
+    -0.001443002705210778
+     -0.00108712945926925
+     -0.02443494593188546
+       0.1410697667490356
+ 1.76e+10    
+       0.1421786111918923
+     -0.02454912501027422
+       0.1431070414858472
+    -0.001102084721142997
+    -0.009538423207401166
+       0.1431160174091101
+    -0.001460225832098509
+    -0.001100463468629002
+     -0.02457095033352142
+         0.14183448563495
+ 1.77e+10    
+       0.1429445813732787
+     -0.02468531834860674
+       0.1438828964285377
+    -0.001115437587459313
+     -0.00960307883472121
+        0.143891790518731
+    -0.001477330181493255
+    -0.001113769405437537
+     -0.02470724527324238
+       0.1425988030464501
+ 1.78e+10    
+        0.143710116383036
+     -0.02482178713777382
+       0.1446581314642348
+     -0.00112876904770835
+    -0.009668240001192308
+        0.144666970749997
+    -0.001494316098777429
+    -0.001127052832546896
+     -0.02484382578951272
+       0.1433627153546904
+ 1.79e+10    
+       0.1444752127666319
+     -0.02495852616885191
+       0.1454327386579624
+    -0.001142084717896712
+    -0.009733887951894556
+        0.145441550575435
+    -0.001511184028428964
+    -0.001140319365612079
+     -0.02498068668473855
+       0.1441262188661882
+ 1.8e+10     
+       0.1452398670383958
+     -0.02509553002382353
+       0.1462067103601035
+    -0.001155390254314099
+    -0.009800003869717924
+       0.1462155227365705
+    -0.001527934510485549
+    -0.001153574660584787
+     -0.02511782254421226
+       0.1448893098288379
+ 1.81e+10    
+        0.146004075686163
+     -0.02523279309389054
+       0.1469800392154992
+    -0.001168691341560909
+    -0.009866568918879702
+       0.1469888802527357
+     -0.00154456817702207
+    -0.001166824401748428
+     -0.02525522775463915
+       0.1456519844377331
+ 1.82e+10    
+       0.1467678351757314
+     -0.02537030959735715
+       0.1477527181717876
+    -0.001181993681113793
+    -0.009933564286135885
+       0.1477616164290885
+    -0.001561085748642007
+    -0.001180074290291525
+     -0.02539289652222636
+       0.1464142388407983
+ 1.83e+10    
+       0.1475311419551293
+     -0.02550807359706276
+       0.1485247404869797
+    -0.001195302980429194
+     -0.01000097121970187
+       0.1485337248638566
+    -0.001577488030982346
+    -0.001193330033423022
+     -0.02553082289031269
+       0.1471760691442239
+ 1.84e+10    
+        0.148293992458696
+     -0.02564607901734894
+       0.1492960997362928
+    -0.001208624942579331
+     -0.01006877106590992
+       0.1493051994548114
+    -0.001593775911234179
+    -0.001206597334020403
+     -0.02566900075652289
+       0.1479374714177022
+ 1.85e+10    
+        0.149056383110973
+     -0.02578431966054385
+       0.1500667898182439
+    -0.001221965256416489
+      -0.0101369453036333
+       0.1500760344049908
+    -0.001609950354679086
+    -0.001219881880809831
+     -0.02580742388943238
+       0.1486984416994689
+ 1.86e+10    
+       0.1498183103304135
+      -0.0259227892229543
+       0.1508368049600207
+    -0.001235329587259515
+     -0.01020547557651701
+       0.1508462242276811
+    -0.001626012401243183
+     -0.00123318933906867
+     -0.02594608594472925
+       0.1494589760011444
+ 1.87e+10    
+       0.1505797705329044
+     -0.02606148131035261
+       0.1516061397221418
+    -0.001248723568093658
+     -0.01027434372305748
+       0.1516157637506734
+    -0.001641963162069784
+    -0.001246525341844149
+     -0.02608498048086345
+       0.1502190703123769
+ 1.88e+10    
+       0.1513407601351085
+     -0.02620038945295154
+       0.1523747890024203
+    -0.001262152791275608
+     -0.01034353180458009
+       0.1523846481198118
+    -0.001657803816112412
+    -0.001259895481678363
+     -0.02622410097417494
+       0.1509787206052906
+ 1.89e+10    
+       0.1521012755576281
+     -0.02633950711985932
+       0.1531427480392454
+    -0.001275622800733269
+     -0.01041302213116675
+       0.1531528728018487
+     -0.00167353560674955
+    -0.001273305302830048
+      -0.0263634408334941
+       0.1517379228387349
+ 1.9e+10     
+       0.1528613132279907
+     -0.02647882773301136
+       0.1539100124142007
+    -0.001289139084649145
+     -0.01048279728559035
+       0.1539204335866284
+    -0.001689159838423356
+    -0.001286760293979772
+     -0.02650299341421022
+       0.1524966729623409
+ 1.91e+10    
+       0.1536208695834634
+     -0.02661834468057387
+       0.1546765780540297
+     -0.00130270706861517
+     -0.01055284014531379
+       0.1546873265886105
+    -0.001704677873303404
+    -0.001300265881410224
+     -0.02664275203180411
+       0.1532549669203858
+ 1.92e+10    
+       0.1543799410736955
+      -0.0267580513298183
+       0.1554424412319743
+    -0.001316332109248012
+     -0.01062313390261684
+        0.155453548247762
+    -0.001720091127977732
+    -0.001313827422645496
+     -0.02678270997484474
+       0.1540128006554668
+ 1.93e+10    
+       0.1551385241631979
+     -0.02689794103946691
+       0.1562075985684946
+    -0.001330019488249756
+     -0.01069366208291231
+       0.1562190953298279
+    -0.001735401070172803
+    -0.001327450200538923
+     -0.02692286051744808
+       0.1547701701119873
+ 1.94e+10    
+       0.1558966153336555
+     -0.02703800717150841
+       0.1569720470313931
+    -0.001343774406901485
+       -0.010764408561319
+       0.1569839649260061
+     -0.00175060921550455
+     -0.00134113941779332
+     -0.02706319693120122
+       0.1555270712394598
+ 1.95e+10    
+        0.156654211086086
+     -0.02717824310248823
+        0.157735783935362
+    -0.001357601980976672
+      -0.0108353575775555
+       0.1577481544520462
+    -0.001765717124261851
+    -0.001354900191901882
+     -0.02720371249655316
+       0.1562834999956272
+ 1.96e+10    
+       0.1574113079428408
+     -0.02731864223427522
+        0.158498806940968
+    -0.001371507236058077
+     -0.01090649374922335
+       0.1585116616467896
+    -0.001780726398224733
+    -0.001368737550494006
+     -0.02734440051367642
+       0.1570394523494077
+ 1.97e+10    
+       0.1581679024494579
+     -0.02745919800430915
+       0.1592611140530961
+     -0.00138549510324615
+     -0.01097780208354608
+       0.1592744845701753
+    -0.001795638677518937
+    -0.001382656427071703
+     -0.02748525431280384
+       0.1577949242836646
+ 1.98e+10    
+       0.1589239911763671
+     -0.02759990389533499
+       0.1600227036188699
+     -0.00139957041524201
+     -0.01104926798763216
+       0.1600366216007297
+    -0.001810455637508637
+    -0.001396661657122798
+     -0.02762626726404735
+       0.1585499117978079
+ 1.99e+10    
+       0.1596795707204553
+     -0.02774075344462933
+       0.1607835743250668
+    -0.001413737902792966
+     -0.01112087727732872
+       0.1607980714325607
+    -0.001825178985729044
+    -0.001410757974594923
+     -0.02776743278670354
+         0.15930441091023
+ 2e+10       
+       0.1604346377064944
+     -0.02788174025272694
+       0.1615437251950482
+     -0.00142800219148377
+     -0.01119261618473328
+       0.1615588330718818
+    -0.001839810458860661
+    -0.001424950008716696
+     -0.02790874435805577
+        0.160058417660579
+ 2.01e+10    
+       0.1611891887884367
+     -0.02802285799165375
+       0.1623031555852199
+    -0.001442367798860222
+     -0.01126447136442953
+       0.1623189058330778
+    -0.001854351819746811
+    -0.001439242281150427
+     -0.02805019552167856
+       0.1608119281118774
+ 2.02e+10    
+       0.1619432206505827
+     -0.02816410041267589
+       0.1630618651810452
+    -0.001456839131870335
+     -0.01133642989851221
+       0.1630782893343429
+    -0.001868804854455979
+    -0.001453639203463266
+     -0.02819177989525551
+       0.1615649383524868
+ 2.03e+10    
+       0.1626967300086252
+     -0.02830546135357268
+       0.1638198539926263
+    -0.001471420484609278
+     -0.01140847930046558
+       0.1638369834929037
+    -0.001883171369390445
+    -0.001468145074900203
+     -0.02833349117791791
+       0.1623174444979238
+ 2.04e+10    
+       0.1634497136105771
+     -0.02844693474544431
+        0.164577122349873
+    -0.001486116036353342
+     -0.01148060751795822
+       0.1645949885198525
+    -0.001897453188442696
+    -0.001482764080447414
+     -0.02847532315711602
+       0.1630694426925371
+ 2.05e+10    
+       0.1642021682375815
+     -0.02858851461906231
+       0.1653336708972767
+    -0.001500929849869164
+     -0.01155280293461593
+       0.1653523049146073
+    -0.001911652150200996
+    -0.001497500289169025
+     -0.02861726971503209
+       0.1638209291110407
+ 2.06e+10    
+       0.1649540907046169
+     -0.02873019511077482
+       0.1660895005883075
+    -0.001515865869984424
+     -0.01162505437083283
+       0.1661089334590223
+    -0.001925770105205544
+    -0.001512357652806015
+     -0.02875932483454668
+        0.164571899959918
+ 2.07e+10    
+       0.1657054778610939
+     -0.02887197046797651
+       0.1668446126794525
+    -0.001530927922408538
+      -0.0116973510836787
+       0.1668648752111644
+    -0.001939808913255651
+    -0.001527340004622832
+     -0.02890148260476904
+       0.1653223514786938
+ 2.08e+10    
+       0.1664563265913546
+      -0.0290138350541544
+       0.1675990087239129
+    -0.001546119712786694
+     -0.01176968276596033
+       0.1676201314987793
+    -0.001953770440770396
+    -0.001542451058487652
+     -0.02904373722614381
+        0.166072279941084
+ 2.09e+10    
+       0.1672066338150749
+     -0.02915578335352044
+       0.1683526905649745
+    -0.001561444825977967
+     -0.01184203954449082
+        0.168374703912461
+     -0.00196765655820236
+    -0.001557694408175938
+     -0.02918608301514457
+        0.166821681656026
+ 2.1e+10     
+       0.1679563964875765
+     -0.02929780997524333
+       0.1691056603290729
+    -0.001576906725543821
+     -0.01191441197762102
+       0.1691285942985509
+    -0.001981469137506355
+    -0.001573073526881677
+     -0.02932851440856787
+       0.1675705529685925
+ 2.11e+10    
+       0.1687056116000502
+     -0.02943990965728933
+       0.1698579204185677
+    -0.001592508753433761
+     -0.01198679105208445
+       0.1698818047517764
+    -0.001995210049663542
+    -0.001588591766927346
+     -0.02947102596743814
+       0.1683188902607978
+ 2.12e+10    
+        0.169454276179701
+     -0.02958207726988678
+       0.1706094735042407
+    -0.001608254129859316
+     -0.01205916817920453
+       0.1706343376076546
+    -0.002008881162261986
+    -0.001604252359657814
+      -0.0296136123805372
+       0.1690666899522976
+ 2.13e+10    
+       0.1702023872898093
+     -0.02972430781862289
+       0.1713603225175388
+    -0.001624145953342316
+     -0.01213153519051314
+       0.1713861954346749
+    -0.002022484337133824
+    -0.001620058415509875
+     -0.02975626846757006
+       0.1698139485009876
+ 2.14e+10    
+       0.1709499420297233
+     -0.02986659644718718
+       0.1721104706425721
+    -0.001640187200928225
+     -0.01220388433282496
+       0.1721373810262791
+    -0.002036021428050293
+    -0.001636012924244038
+     -0.02989898918197925
+       0.1705606624035076
+ 2.15e+10    
+       0.1716969375347785
+     -0.03000893843977306
+       0.1728599213078889
+     -0.00165638072855362
+     -0.01227620826281291
+       0.1728878973926554
+    -0.002049494278474714
+    -0.001652118755328555
+     -0.03004176961342072
+       0.1713068281956523
+ 2.16e+10    
+       0.1724433709761519
+     -0.03015132922314876
+       0.1736086781780382
+    -0.001672729271556949
+     -0.01234850004112572
+       0.1736377477523656
+    -0.002062904719373837
+    -0.001668378658467216
+     -0.03018460498991331
+       0.1720524424526958
+ 2.17e+10    
+       0.1731892395606546
+     -0.03029376436841041
+       0.1743567451449377
+    -0.001689235445324855
+     -0.01242075312608844
+       0.1743869355238193
+    -0.002076254567088084
+    -0.001684795264258093
+     -0.03032749067967449
+       0.1727975017896341
+ 2.18e+10    
+       0.1739345405304659
+     -0.03043623959242903
+       0.1751041263190612
+    -0.001705901746061802
+     -0.01249296136702418
+       0.1751354643166124
+    -0.002089545621260938
+    -0.001701371084976586
+     -0.03047042219265429
+       0.1735420028613467
+ 2.19e+10    
+       0.1746792711628133
+     -0.03057875075900343
+       0.1758508260204626
+    -0.001722730551676909
+     -0.01256511899723373
+       0.1758833379227461
+    -0.002102779662827468
+    -0.001718108515472036
+      -0.0306133951817803
+       0.1742859423626865
+ 2.2e+10     
+       0.1754234287696002
+     -0.03072129387973047
+       0.1765968487696469
+    -0.001739724122777331
+     -0.01263722062666781
+       0.1766305603077413
+    -0.002115958452062298
+    -0.001735009834170187
+     -0.03075640544392509
+       0.1750293170284969
+ 2.21e+10    
+       0.1761670106969887
+      -0.0308638651146052
+        0.177342199278308
+    -0.001756884603761356
+     -0.01270926123432558
+       0.1773771356016645
+    -0.002129083726687066
+    -0.001752077204172356
+     -0.03089944892060936
+       0.1757721236335649
+ 2.22e+10    
+       0.1769100143249365
+     -0.03100646077236165
+       0.1780868824399435
+     -0.00177421402400197
+     -0.01278123616041007
+       0.1781230680900792
+    -0.002142157200037238
+    -0.001769312674444434
+     -0.03104252169845109
+       0.1765143589925103
+ 2.23e+10    
+       0.1776524370666935
+     -0.03114907731056607
+       0.1788309033203604
+     -0.00179171429911527
+     -0.01285314109827093
+       0.1788683622049364
+    -0.002155180559288205
+    -0.001786718181087458
+     -0.03118562000937374
+       0.1772560199596166
+ 2.24e+10    
+       0.1783942763682611
+     -0.03129171133547464
+       0.1795742671480905
+    -0.001809387232304687
+     -0.01292497208616279
+       0.1796130225154223
+    -0.002168155463740499
+    -0.001804295548683155
+      -0.0313287402305847
+       0.1779971034286068
+ 2.25e+10    
+       0.1791355297078183
+     -0.03143435960166579
+        0.180316979304723
+    -0.001827234515775326
+     -0.01299672549884562
+       0.1803570537187711
+    -0.002181083543164239
+    -0.001822046491706139
+       -0.031471878884335
+       0.1787376063323692
+ 2.26e+10    
+       0.1798761945951142
+     -0.03157701901145869
+       0.1810590453151727
+    -0.001845257732211951
+     -0.01306839803905244
+       0.1811004606310637
+    -0.002193966396201816
+    -0.001839972615999221
+     -0.03161503263747197
+       0.1794775256426331
+ 2.27e+10    
+       0.1806162685708337
+      -0.0317196866141291
+       0.1818004708378929
+    -0.001863458356313828
+     -0.01313998672884807
+       0.1818432481780169
+    -0.002206805588829265
+    -0.001858075420302191
+     -0.03175819830079574
+       0.1802168583696022
+ 2.28e+10    
+       0.1813557492059374
+     -0.03186235960493269
+       0.1825412616550507
+    -0.001881837756381022
+     -0.01321148890090164
+       0.1825854213857844
+      -0.0022196026528755
+     -0.00187635629783074
+     -0.03190137282822986
+       0.1809556015615446
+ 2.29e+10    
+       0.1820946341009782
+     -0.03200503532394662
+        0.183281423662673
+    -0.001900397195947065
+     -0.01328290218969333
+       0.1833269853717787
+     -0.00223235908459901
+    -0.001894816537899304
+     -0.03204455331581767
+       0.1816937523043475
+ 2.3e+10     
+       0.1828329208853967
+     -0.03214771125473954
+       0.1840209628607806
+    -0.001919137835451581
+     -0.01335422452267561
+       0.1840679453355209
+    -0.002245076343321747
+    -0.001913457327581821
+     -0.03218773700055316
+       0.1824313077210341
+ 2.31e+10    
+       0.1835706072168004
+     -0.03229038502288032
+       0.1847598853435185
+    -0.001938060733949769
+     -0.01342545411140709
+       0.1848083065495423
+    -0.002257755850119341
+    -0.001932279753406858
+     -0.03233092125905831
+         0.18316826497125
+ 2.32e+10    
+       0.1843076907802265
+     -0.03243305439429537
+       0.1854981972893005
+    -0.001957166850851287
+      -0.0134965894426771
+       0.1855480743503383
+    -0.002270398986567598
+    -0.001951284803081224
+     -0.03247410360611516
+       0.1839046212507209
+ 2.33e+10    
+        0.185044169287391
+     -0.03257571727348397
+       0.1862359049509724
+    -0.001976457047687809
+     -0.01356762926963577
+       0.1862872541293907
+    -0.002283007093544084
+    -0.001970473367238245
+     -0.03261728169306287
+       0.1846403737906822
+ 2.34e+10    
+       0.1857800404759274
+     -0.03271837170160111
+       0.1869730146460147
+    -0.001995932089901549
+     -0.01363857260294641
+       0.1870258513242688
+    -0.002295581470084611
+    -0.001989846241206785
+     -0.03276045330606896
+       0.1853755198572856
+ 2.35e+10    
+       0.1865153021086169
+     -0.03286101585441736
+       0.1877095327467904
+    -0.002015592648653444
+     -0.01370941870197297
+       0.1877638714098224
+    -0.002308123372293627
+     -0.00200940412679722
+      -0.0329036163642845
+       0.1861100567509854
+ 2.36e+10    
+         0.18724995197261
+     -0.03300364804016491
+       0.1884454656708531
+    -0.002035439302645548
+     -0.01378016706601694
+       0.1885013198894702
+    -0.002320634012308324
+     -0.00202914763409889
+     -0.03304676891789055
+       0.1868439818059038
+ 2.37e+10    
+       0.1879839878786458
+     -0.03314626669727736
+       0.1891808198713245
+    -0.002055472539955609
+     -0.01385081742561428
+       0.1892382022866031
+    -0.002333114557314982
+    -0.002049077283289116
+     -0.03318990914604658
+       0.1875772923891821
+ 2.38e+10    
+       0.1887174076602644
+      -0.0332888703920339
+       0.1899156018273552
+    -0.002075692759879537
+     -0.01392136973390521
+       0.1899745241361026
+    -0.002345566128617375
+    -0.002069193506447797
+     -0.03333303535474653
+       0.1883099859003143
+ 2.39e+10    
+       0.1894502091730222
+     -0.03343145781611408
+       0.1906498180346776
+     -0.00209610027477999
+     -0.01399182415808624
+       0.1907102909759909
+    -0.002357989800756234
+     -0.00208949664937505
+     -0.03347614597459365
+       0.1890420597704728
+ 2.4e+10     
+        0.190182390293704
+     -0.03357402778407269
+       0.1913834749962639
+     -0.00211669531193599
+     -0.01406218107095484
+       0.1914455083392186
+    -0.002370386600679206
+     -0.00210998697341035
+     -0.03361923955849917
+       0.1897735114618203
+ 2.41e+10    
+       0.1909139489195388
+     -0.03371657923074212
+       0.1921165792130989
+    -0.002137478015393879
+     -0.01413244104255488
+       0.1921801817455982
+     -0.00238275750696003
+    -0.002130664657249402
+      -0.0337623147793136
+       0.1905043384668143
+ 2.42e+10    
+       0.1916448829674174
+     -0.03385911120856981
+       0.1928491371750779
+    -0.002158448447815208
+     -0.01420260483193157
+       0.1929143166938941
+    -0.002395103449066407
+    -0.002151529798756919
+     -0.03390537042739898
+       0.1912345383075079
+ 2.43e+10    
+       0.1923751903731166
+     -0.03400162288489823
+       0.1935811553520404
+    -0.002179606592318984
+     -0.01427267337900274
+       0.1936479186540732
+    -0.002407425306675902
+    -0.002172582416773209
+     -0.03404840540814606
+        0.191964108534841
+ 2.44e+10    
+       0.1931048690905283
+     -0.03414411353919451
+        0.194312640184951
+     -0.00220095235431872
+     -0.01434264779655412
+       0.1943809930597303
+    -0.002419723909038404
+    -0.002193822452911727
+     -0.03419141873944702
+       0.1926930467279338
+ 2.45e+10    
+       0.1938339170908961
+     -0.03428658256023736
+        0.195043598077234
+    -0.002222485563348281
+      -0.0144125293623639
+       0.1951135453006869
+    -0.002432000034385025
+    -0.002215249773346918
+     -0.03433440954912688
+       0.1934213504933745
+ 2.46e+10    
+       0.1945623323620596
+     -0.03442902944326606
+       0.1957740353862748
+    -0.002244205974878937
+     -0.01448231951146248
+       0.1958455807157796
+    -0.002444254409381802
+    -0.002236864170589974
+     -0.03447737707234239
+       0.1941490174645101
+ 2.47e+10    
+       0.1952901129077109
+     -0.03457145378710091
+       0.1965039584150958
+    -0.002266113272122842
+     -0.01455201982853282
+       0.1965771045858368
+     -0.00245648770862803
+      -0.0022586653652502
+     -0.03462032064895269
+       0.1948760453007386
+ 2.48e+10    
+       0.1960172567466591
+     -0.03471385529123876
+       0.1972333734042145
+    -0.002288207067823042
+      -0.0146216320404551
+       0.1973081221268561
+    -0.002468700554197548
+    -0.002280653007782579
+     -0.03476323972086819
+       0.1956024316868006
+ 2.49e+10    
+        0.196743761912108
+     -0.03485623375293094
+        0.197962286523697
+    -0.002310486906028014
+     -0.01469115800900069
+       0.1980386384833833
+    -0.002480893515222894
+    -0.002302826680217579
+     -0.03490613382938366
+       0.1963281743320804
+ 2.5e+10     
+       0.1974696264509454
+     -0.03499858906424885
+       0.1986907038654075
+    -0.002332952263848945
+     -0.01476059972367781
+        0.198768658722103
+    -0.002493067107520837
+    -0.002325185897874327
+     -0.03504900261249966
+       0.1970532709699078
+ 2.51e+10    
+       0.1981948484230475
+     -0.03514092120914391
+       0.1994186314354714
+    -0.002355602553199943
+     -0.01482995929473318
+       0.1994981878256435
+    -0.002505221793258421
+    -0.002347730111055067
+     -0.03519184580223868
+       0.1977777193568685
+ 2.52e+10    
+       0.1989194259005959
+      -0.0352832302605051
+       0.2001460751469513
+    -0.002378437122519083
+     -0.01489923894631136
+       0.2002272306865994
+    -0.002517357980659024
+    -0.002370458706718972
+      -0.0353346632219593
+       0.1985015172721219
+ 2.53e+10    
+       0.1996433569674106
+      -0.0354255163772214
+       0.2008730408127495
+    -0.002401455258469101
+     -0.01496844100977449
+       0.2009557921017807
+    -0.002529476023746874
+    -0.002393371010137438
+     -0.03547745478367471
+       0.1992246625167269
+ 2.54e+10    
+       0.2003666397182981
+     -0.03556777980125275
+       0.2015995341387389
+    -0.002424656187616972
+     -0.01503756791718495
+       0.2016838767666891
+    -0.002541576222130015
+    -0.002416466286525351
+     -0.03562022048537808
+       0.1999471529129765
+ 2.55e+10    
+       0.2010892722584169
+     -0.03571002085471423
+       0.2023255607171337
+     -0.00244803907809331
+     -0.01510662219495077
+       0.2024114892702253
+     -0.00255365882081964
+    -0.002439743742652937
+     -0.03576296040838035
+       0.2006689863037432
+ 2.56e+10    
+       0.2018112527026589
+     -0.03585223993697858
+       0.2030511260201038
+    -0.002471603041227578
+     -0.01517560645763712
+       0.2031386340896319
+    -0.002565724010085963
+    -0.002463202528433996
+     -0.03590567471466352
+       0.2013901605518361
+ 2.57e+10    
+       0.2025325791750477
+     -0.03599443752180069
+       0.2037762353936362
+     -0.00249534713316158
+     -0.01524452340194336
+       0.2038653155856749
+    -0.002577771925349209
+     -0.00248684173849021
+      -0.0360483636442533
+       0.2021106735393668
+ 2.58e+10    
+       0.2032532498081568
+     -0.03613661415446794
+       0.2045008940516552
+    -0.002519270356438767
+     -0.01531337580084679
+        0.204591537998065
+    -0.002589802647104823
+    -0.002510660413693392
+     -0.03619102751261485
+       0.2028305231671314
+ 2.59e+10    
+       0.2039732627425446
+     -0.03627877044898125
+       0.2052251070704014
+    -0.002543371661569481
+     -0.01538216649791345
+       0.2053173054411213
+    -0.002601816200882163
+    -0.002534657542683318
+     -0.03633366670807414
+       0.2035497073540011
+ 2.6e+10     
+       0.2046926161262072
+     -0.03642090708526877
+       0.2059488793830749
+    -0.002567649948572186
+     -0.01545089840177598
+       0.2060426218996804
+    -0.002613812557235734
+    -0.002558832063360911
+     -0.03647628168926889
+       0.2042682240363302
+ 2.61e+10    
+       0.2054113081140534
+     -0.03656302480643712
+       0.2066722157747489
+    -0.002592104068489327
+      -0.0155195744807785
+       0.2067674912252512
+    -0.002625791631768181
+    -0.002583182864357134
+     -0.03661887298263147
+       0.2049860711673753
+ 2.62e+10    
+        0.206129336867395
+     -0.03670512441606247
+        0.207395120877555
+    -0.002616732824878418
+     -0.01558819775778776
+       0.2074919171324153
+    -0.002637753285183996
+    -0.002607708786477548
+     -0.03676144117990548
+       0.2057032467167288
+ 2.63e+10    
+       0.2068467005534596
+      -0.0368472067755243
+       0.2081175991661459
+    -0.002641534975277256
+     -0.01565677130517068
+       0.2082159031954777
+    -0.002649697323373228
+    -0.002632408624121984
+     -0.03690398693570093
+       0.2064197486697689
+ 2.64e+10    
+       0.2075633973449211
+     -0.03698927280138548
+       0.2088396549534372
+    -0.002666509232643812
+     -0.01572529823993668
+       0.2089394528453616
+    -0.002661623497524433
+    -0.002657281126679057
+     -0.03704651096508696
+       0.2071355750271228
+ 2.65e+10    
+       0.2082794254194513
+     -0.03713132346282005
+       0.2095612923866285
+    -0.002691654266770799
+     -0.01579378171904404
+       0.2096625693667544
+    -0.002673531504265708
+    -0.002682324999895958
+     -0.03718901404122697
+        0.207850723804145
+ 2.66e+10    
+       0.2089947829592917
+     -0.03727335977909227
+       0.2102825154435113
+    -0.002716968705673148
+     -0.01586222493486963
+       0.2103852558954978
+    -0.002685420985833567
+     -0.00270753890722307
+     -0.03733149699305656
+       0.2085651930304135
+ 2.67e+10    
+       0.2097094681508421
+     -0.03741538281708767
+       0.2110033279290587
+    -0.002742451136950885
+     -0.01593063111083989
+       0.2111075154162277
+     -0.00269729153026802
+    -0.002732921471134443
+      -0.0374739607030064
+       0.2092789807492376
+ 2.68e+10    
+       0.2104234791842748
+     -0.03755739368889983
+        0.211723733472304
+    -0.002768100109125263
+      -0.0159990034972219
+       0.2118293507602555
+    -0.002709142671634115
+    -0.002758471274421845
+      -0.0376164061047715
+       0.2099920850171859
+ 2.69e+10    
+       0.2111368142531627
+     -0.03769939354947242
+       0.2124437355235018
+    -0.002793914132948635
+     -0.01606734536707284
+       0.2125507646036955
+    -0.002720973890268019
+    -0.002784186861466463
+     -0.03775883418112772
+       0.2107045039036264
+ 2.7e+10     
+       0.2118494715541321
+     -0.03784138359430056
+       0.2131633373515797
+    -0.002819891682689605
+     -0.01613566001234626
+       0.2132717594658338
+    -0.002732784613047954
+    -0.002810066739483206
+     -0.03790124596179845
+       0.2114162354902851
+ 2.71e+10    
+        0.212561449286532
+     -0.03798336505719103
+       0.2138825420418736
+    -0.002846031197390599
+     -0.01620395074015264
+       0.2139923377077339
+    -0.002744574213688393
+    -0.002836109379743063
+     -0.03804364252136998
+       0.2121272778708203
+ 2.72e+10    
+       0.2132727456521258
+     -0.03812533920808292
+       0.2146013524941479
+    -0.002872331082101593
+     -0.01627222086917268
+       0.2147125015310848
+    -0.002756342013057156
+    -0.002862313218769608
+     -0.03818602497725885
+        0.212837629150411
+ 2.73e+10    
+        0.213983358854801
+     -0.03826730735093109
+       0.2153197714209018
+    -0.002898789709086573
+     -0.01634047372622096
+       0.2154322529772751
+    -0.002768087279514825
+     -0.00288867665951203
+     -0.03832839448772956
+       0.2135472874453637
+ 2.74e+10    
+       0.2146932871002983
+     -0.03840927082165115
+       0.2160378013459551
+     -0.00292540541900514
+     -0.01640871264295783
+        0.216151593926705
+    -0.002779809229275334
+    -0.002915198072494577
+     -0.03847075224996575
+       0.2142562508827343
+ 2.75e+10    
+       0.2154025285959602
+      -0.0385512309861282
+       0.2167554446033148
+    -0.002952176522069094
+     -0.01647694095274684
+       0.2168705260983223
+    -0.002791507026787458
+    -0.002941875796941527
+     -0.03861309949819365
+       0.2149645175999642
+ 2.76e+10    
+       0.2161110815505003
+     -0.03869318923829029
+       0.2174727033363192
+     -0.00297910129917374
+     -0.01654516198765515
+       0.2175890510493807
+    -0.002803179785136123
+    -0.002968708141880008
+      -0.0387554375018581
+       0.2156720857445355
+ 2.77e+10    
+       0.2168189441737872
+     -0.03883514699824449
+       0.2181895794970554
+    -0.003006178003003542
+     -0.01661337907559534
+       0.2183071701754193
+    -0.002814826566463392
+    -0.002995693387218834
+     -0.03889776756385245
+       0.2163789534736387
+ 2.78e+10    
+        0.217526114676651
+     -0.03897710571047901
+       0.2189060748460461
+    -0.003033404859114408
+     -0.01668159553760424
+        0.219024884710456
+    -0.002826446382407836
+    -0.003022829784804898
+     -0.03904009101880123
+       0.2170851189538571
+ 2.79e+10    
+        0.218232591270706
+     -0.03911906684212969
+       0.2196221909522048
+    -0.003060780066990866
+     -0.01674981468525772
+       0.2197421957273907
+    -0.002838038194562099
+    -0.003050115559457134
+     -0.03918240923139641
+       0.2177905803608658
+ 2.8e+10     
+       0.2189383721681914
+     -0.03926103188131047
+       0.2203379291930517
+    -0.003088301801078369
+     -0.01681803981821792
+       0.2204591041386149
+    -0.002849600914948032
+    -0.003077548909978226
+       -0.039324723594787
+       0.2184953358791478
+ 2.81e+10    
+       0.2196434555818295
+     -0.03940300233550868
+       0.2210532907551849
+    -0.003115968211793464
+     -0.01688627422190954
+       0.2211756106968199
+    -0.002861133406508394
+    -0.003105128010144518
+     -0.03946703552902087
+        0.219199383701721
+ 2.82e+10    
+        0.220347839724701
+     -0.03954497973004483
+       0.2217682766350084
+    -0.003143777426508779
+     -0.01695452116532365
+       0.2218917159960011
+    -0.002872634483614906
+    -0.003132851009674299
+     -0.03960934647953955
+       0.2199027220298827
+ 2.83e+10    
+       0.2210515228101371
+     -0.03968696560659549
+       0.2224828876397018
+    -0.003171727550515461
+     -0.01702278389894468
+       0.2226074204726504
+    -0.002884102912592092
+    -0.003160716035174612
+     -0.03975165791572523
+       0.2206053490729685
+ 2.84e+10    
+       0.2217545030516282
+     -0.03982896152177939
+       0.2231971243884312
+    -0.003199816667962885
+     -0.01709106565279829
+       0.2233227244071335
+    -0.002895537412255809
+    -0.003188721191067929
+     -0.03989397132949926
+       0.2213072630481226
+ 2.85e+10    
+       0.2224567786627467
+     -0.03997096904580619
+       0.2239109873137972
+     -0.00322804284277446
+      -0.0171593696346173
+       0.2240376279252417
+    -0.002906936654466764
+    -0.003216864560497376
+     -0.04003628823397091
+       0.2220084621800838
+ 2.86e+10    
+        0.223158347857089
+     -0.04011298976118694
+       0.2246244766635071
+    -0.003256404119543204
+     -0.01722769902812171
+       0.2247521309999184
+    -0.002918299264697511
+    -0.003245144206212353
+     -0.04017861016213752
+       0.2227089447009845
+ 2.87e+10    
+       0.2238592088482273
+     -0.04025502526150487
+       0.2253375925022712
+    -0.003284898524403432
+     -0.01729605699141102
+        0.225466233453149
+    -0.002929623822613261
+    -0.003273558171433703
+     -0.04032093866563319
+       0.2234087088501617
+ 2.88e+10    
+        0.224559359849681
+     -0.04039707715024659
+       0.2260503347139091
+    -0.003313524065881352
+     -0.01736444665546426
+       0.2261799349580094
+    -0.002940908862665539
+    -0.003302104480699914
+     -0.04046327531352654
+       0.2241077528739819
+ 2.89e+10    
+       0.2252587990748981
+     -0.04053914703969128
+       0.2267627030036662
+    -0.003342278735724987
+     -0.01743287112274598
+        0.226893235040866
+    -0.002952152874698021
+    -0.003330781140693566
+     -0.04060562169116589
+        0.224806075025677
+ 2.9e+10     
+       0.2259575247372537
+     -0.04068123654985827
+       0.2274746969007264
+    -0.003371160509712631
+     -0.01750133346591381
+       0.2276061330837227
+    -0.002963354304564631
+    -0.003359586141049182
+     -0.04074797939907152
+       0.2255036735651937
+ 2.91e+10    
+       0.2266555350500577
+     -0.04082334730750965
+       0.2281863157609162
+    -0.003400167348440884
+     -0.01756983672662566
+       0.2283186283267059
+    -0.002974511554758763
+    -0.003388517455142265
+     -0.04089035005187346
+       0.2262005467590515
+ 2.92e+10    
+       0.2273528282265781
+     -0.04096548094520971
+       0.2288975587695929
+    -0.003429297198091672
+     -0.01763838391444233
+       0.2290307198706805
+    -0.002985622985053874
+    -0.003417573040860482
+     -0.04103273527729367
+       0.2268966928802163
+ 2.93e+10    
+       0.2280494024800755
+     -0.04110763910043568
+       0.2296084249447036
+    -0.003458547991180967
+     -0.01770697800582287
+       0.2297424066799919
+    -0.002996686913154219
+    -0.003446750841356235
+     -0.04117513671517245
+       0.2275921102079799
+ 2.94e+10    
+       0.2287452560238486
+     -0.04124982341474273
+        0.230318913140017
+    -0.003487917647286668
+     -0.01777562194320985
+       0.2304536875853254
+    -0.003007701615355914
+    -0.003476048785782395
+     -0.04131755601653607
+       0.2282867970278536
+ 2.95e+10    
+       0.2294403870712907
+     -0.04139203553297809
+       0.2310290220485059
+    -0.003517404073758019
+     -0.01784431863420037
+       0.2311645612866776
+    -0.003018665327217541
+    -0.003505464790010135
+     -0.04145999484270715
+       0.2289807516314688
+ 2.96e+10    
+       0.2301347938359573
+     -0.04153427710254481
+       0.2317387502058835
+     -0.00354700516640549
+      -0.0179130709508013
+       0.2318750263564305
+    -0.003029576244240216
+    -0.003534996757330159
+     -0.04160245486445352
+       0.2296739723164914
+ 2.97e+10    
+       0.2308284745316434
+     -0.04167654977271325
+        0.232448095994277
+    -0.003576718810173439
+     -0.01798188172876353
+       0.2325850812425228
+    -0.003040432522556087
+    -0.003564642579137276
+     -0.04174493776117626
+       0.2303664573865392
+ 2.98e+10    
+       0.2315214273724699
+     -0.04181885519397748
+       0.2331570576460353
+    -0.003606542879793763
+     -0.01805075376699436
+        0.233294724271713
+    -0.003051232279625705
+    -0.003594400135598152
+     -0.04188744522013526
+       0.2310582051511129
+ 2.99e+10    
+       0.2322136505729794
+     -0.04196119501745672
+       0.2338656332476566
+    -0.003636475240421863
+     -0.01811968982704329
+       0.2340039536529233
+    -0.003061973594943246
+    -0.003624267296303567
+     -0.04202997893571143
+       0.2317492139255353
+ 3e+10       
+       0.2329051423482396
+     -0.04210357089433861
+       0.2345738207438327
+    -0.003666513748255971
+     -0.01818869263265881
+       0.2347127674806608
+    -0.003072654510749348
+    -0.003654241920904721
+     -0.04217254060870218
+       0.2324394820308946
+ 3.01e+10    
+       0.2335959009139556
+     -0.04224598447536306
+       0.2352816179415944
+    -0.003696656251138836
+     -0.01825776486941353
+       0.2354211637385068
+    -0.003083273032751464
+    -0.003684321859733797
+     -0.04231513194565182
+       0.2331290077939993
+ 3.02e+10    
+       0.2342859244865884
+     -0.04238843741034588
+       0.2359890225145567
+    -0.003726900589142709
+     -0.01832690918439402
+       0.2361291403026706
+    -0.003093827130851096
+    -0.003714504954409694
+     -0.04245775465821346
+       0.2338177895473391
+ 3.03e+10    
+       0.2349752112834813
+     -0.04253093134773799
+       0.2366960320072481
+    -0.003757244595139164
+      -0.0183961281859527
+       0.2368366949455971
+     -0.00310431473987749
+    -0.003744789038428689
+     -0.04260041046254161
+       0.2345058256290497
+ 3.04e+10    
+       0.2356637595229913
+      -0.0426734679342216
+       0.2374026438395193
+    -0.003787686095351205
+     -0.01846542444351899
+        0.237543825339622
+    -0.003114733760327938
+     -0.00377517193774061
+     -0.04274310107871458
+       0.2351931143828901
+ 3.05e+10    
+       0.2363515674246275
+     -0.04281604881433877
+       0.2381088553110204
+    -0.003818222909891716
+     -0.01853480048746683
+       0.2382505290606726
+    -0.003125082059113757
+    -0.003805651471310153
+     -0.04288582823018444
+       0.2358796541582183
+ 3.06e+10    
+       0.2370386332091944
+     -0.04295867563015253
+       0.2388146636057412
+    -0.003848852853284662
+     -0.01860425880903597
+       0.2389568035920028
+    -0.003135357470312129
+    -0.003836225451664838
+     -0.04302859364325461
+       0.2365654433099792
+ 3.07e+10    
+       0.2377249550989391
+     -0.04310135002093749
+       0.2395200657965996
+    -0.003879573734973386
+     -0.01867380186030333
+       0.2396626463279559
+    -0.003145557795923023
+    -0.003866891685428697
+     -0.04317139904658188
+       0.2372504801986932
+ 3.08e+10    
+       0.2384105313177042
+     -0.04324407362289885
+       0.2402250588500771
+    -0.003910383359813047
+     -0.01874343205420324
+       0.2403680545777526
+    -0.003155680806631432
+    -0.003897647973842074
+     -0.04331424617070326
+       0.2379347631904524
+ 3.09e+10    
+       0.2390953600910831
+     -0.04338684806891812
+       0.2409296396308881
+    -0.003941279528548874
+     -0.01881315176459276
+       0.2410730255692945
+    -0.003165724242574121
+    -0.003928492113269136
+     -0.04345713674758524
+       0.2386182906569191
+ 3.1e+10     
+       0.2397794396465803
+     -0.04352967498832309
+       0.2416338049066765
+    -0.003972260038281427
+     -0.01888296332635986
+       0.2417775564529808
+    -0.003175685814111011
+    -0.003959421895690656
+     -0.04360007251019497
+       0.2393010609753304
+ 3.11e+10    
+       0.2404627682137728
+      -0.0436725560066816
+       0.2423375513527316
+    -0.004003322682917058
+     -0.01895286903557193
+       0.2424816443055265
+    -0.003185563202600531
+    -0.003990435109185788
+     -0.04374305519209148
+        0.239983072528505
+ 3.12e+10    
+       0.2411453440244744
+     -0.04381549274561543
+       0.2430408755567144
+    -0.004034465253605906
+     -0.01902287114966247
+       0.2431852861337838
+    -0.003195354061179109
+    -0.004021529538399772
+     -0.04388608652703591
+       0.2406643237048543
+ 3.13e+10    
+       0.2418271653129042
+     -0.04395848682263583
+       0.2437437740233885
+    -0.004065685539166814
+     -0.01909297188765265
+       0.2438884788785549
+    -0.003205056015544121
+    -0.004052702964999787
+     -0.04402916824861954
+       0.2413448128983958
+ 3.14e+10    
+        0.242508230315852
+     -0.04410153985099438
+       0.2444462431793462
+    -0.004096981326499162
+     -0.01916317343040639
+        0.244591219418393
+    -0.003214666664740287
+    -0.004083953168118942
+     -0.04417230208990847
+       0.2420245385087701
+ 3.15e+10    
+       0.2431885372728497
+     -0.04424465343955301
+       0.2451482793777244
+     -0.00412835040098289
+     -0.01923347792091633
+       0.2452935045733904
+    -0.003224183581949208
+    -0.004115277924787714
+     -0.04431548978310388
+         0.24270349894126
+ 3.16e+10    
+       0.2438680844263407
+     -0.04438782919266718
+       0.2458498789029006
+    -0.004159790546865895
+      -0.0193038874646181
+       0.2459953311089388
+      -0.0032336043152818
+    -0.004146675010353894
+     -0.04445873305921607
+       0.2433816926068104
+ 3.17e+10    
+       0.2445468700218498
+     -0.04453106871008267
+       0.2465510379751657
+    -0.004191299547640218
+     -0.01937440412973113
+       0.2466966957394697
+    -0.003242926388573306
+    -0.004178142198891241
+     -0.04460203364775245
+       0.2440591179220529
+ 3.18e+10    
+       0.2452248923081541
+     -0.04467437358684524
+       0.2472517527553646
+    -0.004222875186406233
+     -0.01944502994762408
+       0.2473975951321578
+    -0.003252147302180706
+    -0.004209677263596671
+     -0.04474539327641669
+       0.2447357733093285
+ 3.19e+10    
+       0.2459021495374523
+     -0.04481774541321915
+       0.2479520193494975
+    -0.004254515246225692
+     -0.01951576691320231
+       0.2480980259105937
+    -0.003261264533782522
+    -0.004241277977175797
+     -0.04488881367081984
+       0.2454116571967142
+ 3.2e+10     
+       0.2465786399655351
+     -0.04496118577461612
+       0.2486518338132795
+    -0.004286217510464227
+      -0.0195866169853158
+       0.2487979846584124
+    -0.003270275539180204
+    -0.004272942112218741
+      -0.0450322965542005
+       0.2460867680180494
+ 3.21e+10    
+       0.2472543618519512
+     -0.04510469625153109
+       0.2493511921566489
+    -0.004317979763122409
+     -0.01965758208718587
+       0.2494974679228819
+    -0.003279177753101656
+    -0.004304667441563758
+     -0.04517584364715509
+       0.2467611042129624
+ 3.22e+10    
+        0.247929313460176
+     -0.04524827841948498
+       0.2500500903482205
+    -0.004349799789157342
+     -0.01972866410684815
+       0.2501964722184402
+    -0.003287968590005889
+    -0.004336451738651697
+     -0.04531945666737495
+       0.2474346642268993
+ 3.23e+10    
+       0.2486034930577748
+     -0.04539193384897196
+       0.2507485243196779
+    -0.004381675374792689
+     -0.01979986489761107
+       0.2508949940301853
+     -0.00329664544488943
+    -0.004368292777868975
+     -0.04546313732939204
+       0.2481074465111504
+ 3.24e+10    
+       0.2492768989165674
+     -0.04553566410541138
+       0.2514464899701012
+    -0.004413604307820783
+     -0.01987118627852687
+       0.2515930298173049
+    -0.003305205694093314
+    -0.004400188334881237
+     -0.04560688734432935
+       0.2487794495228786
+ 3.25e+10    
+       0.2499495293127864
+     -0.04567947074910181
+       0.2521439831702234
+     -0.00444558437789265
+     -0.01994263003487516
+       0.2522905760164527
+     -0.00331364669611148
+    -0.004432136186956467
+     -0.04575070841965811
+       0.2494506717251474
+ 3.26e+10    
+       0.2506213825272371
+     -0.04582335533517726
+       0.2528409997666118
+    -0.004477613376800416
+     -0.02001419791865598
+       0.2529876290450607
+    -0.003321965792399582
+    -0.004464134113278674
+     -0.04589460225895892
+       0.2501211115869477
+ 3.27e+10    
+       0.2512924568454519
+     -0.04596731941356421
+       0.2535375355857726
+    -0.004509689098749796
+      -0.0200858916490918
+       0.2536841853045889
+    -0.003330160308184295
+    -0.004496179895251619
+     -0.04603857056168686
+       0.2507907675832232
+ 3.28e+10    
+       0.2519627505578419
+     -0.04611136452893719
+       0.2542335864381673
+    -0.004541809340623367
+     -0.02015771291313655
+       0.2543802411837069
+     -0.00333822755327319
+    -0.004528271316793325
+     -0.04618261502293983
+       0.2514596381948974
+ 3.29e+10    
+       0.2526322619598469
+     -0.04625549222067506
+       0.2549291481221498
+    -0.004573971902235461
+     -0.02022966336599096
+       0.2550757930614071
+    -0.003346164822864505
+     -0.00456040616462098
+     -0.04632673733322928
+       0.2521277219088968
+ 3.3e+10     
+       0.2533009893520786
+     -0.04639970402281292
+       0.2556242164278076
+    -0.004606174586578468
+     -0.02030174463162221
+       0.2557708373100457
+    -0.003353969398356863
+    -0.004592582228527306
+     -0.04647093917825277
+       0.2527950172181753
+ 3.31e+10    
+       0.2539689310404635
+     -0.04654400146399286
+       0.2563187871407127
+    -0.004638415200060132
+     -0.02037395830328681
+       0.2564653702983113
+    -0.003361638548159019
+    -0.004624797301647249
+     -0.04661522223866769
+        0.253461522621735
+ 3.32e+10    
+       0.2546360853363812
+     -0.04668838606740985
+       0.2570128560455758
+    -0.004670691552733649
+     -0.02044630594405656
+       0.2571593883941162
+    -0.003369169528498916
+    -0.004657049180716218
+     -0.04675958818986536
+       0.2541272366246473
+ 3.33e+10    
+       0.2553024505567955
+     -0.04683285935075397
+       0.2577064189298029
+    -0.004703001458518975
+      -0.0205187890873449
+       0.2578528879674115
+    -0.003376559584232312
+    -0.004689335666319645
+     -0.04690403870174568
+       0.2547921577380711
+ 3.34e+10    
+       0.2559680250243869
+     -0.04697742282614673
+       0.2583994715869504
+    -0.004735342735416795
+     -0.02059140923743388
+       0.2585458653929245
+    -0.003383805949650657
+    -0.004721654563134123
+     -0.04704857543849087
+       0.2554562844792699
+ 3.35e+10    
+       0.2566328070676741
+     -0.04712207800007183
+        0.259092009820077
+    -0.004767713205714889
+     -0.02066416786999987
+       0.2592383170528109
+    -0.003390905849287865
+    -0.004754003680160082
+      -0.0471932000583381
+       0.2561196153716268
+ 3.36e+10    
+       0.2572967950211368
+     -0.04726682637330008
+       0.2597840294449926
+    -0.004800110696186764
+     -0.02073706643263842
+       0.2599302393392346
+    -0.003397856498726362
+    -0.004786380830946093
+     -0.04733791421335167
+       0.2567821489446572
+ 3.37e+10    
+       0.2579599872253308
+       -0.047411669440807
+       0.2604755262933997
+    -0.004832533038283298
+     -0.02081010634538592
+       0.2606216286568554
+    -0.003404655105401522
+    -0.004818783833805577
+     -0.04748271954919215
+       0.2574438837340197
+ 3.38e+10    
+       0.2586223820269992
+      -0.0475566086916832
+       0.2611664962159277
+    -0.004864978068317199
+     -0.02088328900123785
+       0.2613124814252394
+    -0.003411298869404914
+    -0.004851210512025153
+     -0.04762761770488436
+       0.2581048182815251
+ 3.39e+10    
+       0.2592839777791788
+     -0.04770164560903725
+       0.2618569350850585
+    -0.004897443627641163
+     -0.02095661576666361
+       0.2620027940811849
+    -0.003417784984285781
+    -0.004883658694065774
+     -0.04777261031258234
+       0.2587649511351417
+ 3.4e+10     
+       0.2599447728412993
+     -0.04784678166988936
+       0.2625468387979438
+    -0.004929927562817894
+     -0.02103008798211619
+       0.2626925630809618
+    -0.003424110637851093
+    -0.004916126213755458
+     -0.04791769899733178
+       0.2594242808489997
+ 3.41e+10    
+       0.2606047655792842
+     -0.04799201834505889
+       0.2632362032791106
+    -0.004962427725785155
+     -0.02110370696253639
+        0.263381784902467
+    -0.003430273012963395
+    -0.004948610910475394
+     -0.04806288537682912
+       0.2600828059833932
+ 3.42e+10    
+       0.2612639543656377
+     -0.04813735709904037
+       0.2639250244830583
+    -0.004994941974013246
+     -0.02117747399785147
+       0.2640704560472953
+    -0.003436269288336859
+    -0.004981110629338027
+     -0.04820817106117747
+       0.2607405251047776
+ 3.43e+10    
+       0.2619223375795324
+     -0.04828279938987243
+       0.2646132983967419
+    -0.005027468170656694
+     -0.02125139035346689
+       0.2647585730427259
+    -0.003442096639330982
+    -0.005013623221358576
+     -0.04835355765263921
+       0.2613974367857669
+ 3.44e+10    
+       0.2625799136068917
+      -0.0484283466689972
+       0.2653010210419503
+    -0.005060004184699992
+     -0.02132545727075162
+       0.2654461324436197
+    -0.003447752238742038
+    -0.005046146543618953
+     -0.04849904674538441
+       0.2620535396051284
+ 3.45e+10    
+       0.2632366808404641
+      -0.0485740003811097
+       0.2659881884775667
+    -0.005092547891096578
+     -0.02139967596751557
+       0.2661331308342376
+    -0.003453233257592074
+    -0.005078678459424934
+     -0.04864463992523552
+       0.2627088321477699
+ 3.46e+10    
+       0.2638926376798951
+     -0.04871976196399842
+       0.2666747968017249
+    -0.005125097170902878
+     -0.02147404763847958
+       0.2668195648299698
+    -0.003458536865915209
+    -0.005111216838456887
+     -0.04879033876940892
+       0.2633633130047339
+ 3.47e+10    
+       0.2645477825317908
+     -0.04886563284837619
+       0.2673608421538537
+    -0.005157649911406113
+     -0.02154857345573721
+       0.2675054310789812
+    -0.003463660233541141
+    -0.005143759556913121
+     -0.04893614484625028
+       0.2640169807731769
+ 3.48e+10    
+       0.2652021138097813
+      -0.0490116144577013
+       0.2680463207166106
+    -0.005190204006246406
+     -0.02162325456920782
+       0.2681907262637757
+    -0.003468600530875903
+    -0.005176304497647522
+     -0.04908205971496825
+       0.2646698340563569
+ 3.49e+10    
+        0.265855629934574
+     -0.04915770820798923
+       0.2687312287177119
+    -0.005222757355533799
+     -0.02169809210708161
+       0.2688754471026744
+    -0.003473354929679368
+    -0.005208849550300123
+     -0.04922808492536217
+       0.2653218714636122
+ 3.5e+10     
+       0.2665083293340031
+     -0.04930391550761457
+       0.2694155624316508
+     -0.00525530786595969
+     -0.02177308717625475
+       0.2695595903512117
+    -0.003477920603839679
+    -0.005241392611421767
+     -0.04937422201754547
+       0.2659730916103375
+ 3.51e+10    
+       0.2671602104430764
+     -0.04945023775710331
+       0.2700993181813132
+    -0.005287853450903237
+     -0.02184824086275644
+        0.270243152803455
+    -0.003482294730144315
+    -0.005273931584592552
+     -0.04952047252166659
+       0.2666234931179601
+ 3.52e+10    
+       0.2678112717040135
+     -0.04959667634891621
+       0.2707824923394865
+    -0.005320392030532337
+     -0.02192355423216565
+       0.2709261312932338
+      -0.0034864744890477
+    -0.005306464380534165
+     -0.04966683795762296
+       0.2672730746139109
+ 3.53e+10    
+       0.2684615115662813
+     -0.04974323266722191
+        0.271465081330266
+    -0.005352921531899719
+     -0.02199902833001928
+       0.2716085226953008
+    -0.003490457065435299
+    -0.005338988917216412
+     -0.04981331983477318
+        0.267921834731595
+ 3.54e+10    
+       0.2691109284866238
+     -0.04988990808766187
+       0.2721470816303624
+     -0.00538543988903448
+     -0.02207466418221044
+       0.2722903239264044
+     -0.00349423964938374
+       -0.005371503119958
+     -0.04995991965164292
+       0.2685697721103554
+ 3.55e+10    
+       0.2697595209290859
+     -0.05003670397710512
+       0.2728284897703025
+    -0.005417945043028421
+     -0.02215046279537674
+       0.2729715319462911
+    -0.003497819436917392
+    -0.005404004921521436
+     -0.05010663889562832
+       0.2692168853954393
+ 3.56e+10    
+       0.2704072873650337
+     -0.05018362169339463
+       0.2735093023355371
+    -0.005450434942117864
+     -0.02222642515727955
+       0.2736521437586278
+    -0.003501193630760732
+    -0.005436492262202634
+      -0.0502534790426943
+       0.2698631732379579
+ 3.57e+10    
+       0.2710542262731708
+     -0.05033066258508567
+       0.2741895159674518
+    -0.005482907541760926
+     -0.02230255223717345
+       0.2743321564118517
+     -0.00350435944108669
+    -0.005468963089915121
+     -0.05040044155706961
+       0.2705086342948463
+ 3.58e+10    
+       0.2717003361395457
+     -0.05047782799117391
+       0.2748691273642806
+    -0.005515360804710279
+     -0.02237884498616556
+       0.2750115669999446
+    -0.003507314086260743
+    -0.005501415360268507
+     -0.05054752789093696
+        0.271153267228817
+ 3.59e+10    
+       0.2723456154575598
+     -0.05062511924081743
+       0.2755481332819291
+    -0.005547792701081545
+     -0.02245530433756599
+       0.2756903726631368
+    -0.003510054793580535
+    -0.005533847036642474
+     -0.05069473948412041
+       0.2717970707083146
+ 3.6e+10     
+        0.272990062727966
+     -0.05077253765304856
+        0.276226530534705
+    -0.005580201208417532
+     -0.02253193120722782
+       0.2763685705885409
+    -0.003512578800011167
+    -0.005566256090255111
+     -0.05084207776376928
+       0.2724400434074671
+ 3.61e+10    
+        0.273633676458867
+     -0.05092008453648009
+       0.2769043159959632
+    -0.005612584311748077
+     -0.02260872649387828
+        0.277046158010716
+    -0.003514883352915787
+    -0.005598640500226341
+     -0.05098954414403752
+       0.2730821840060324
+ 3.62e+10    
+       0.2742764551657056
+     -0.05106776118900241
+       0.2775814865986608
+    -0.005644940003645619
+     -0.02268569107944045
+       0.2777231322121631
+    -0.003516965710781456
+    -0.005630998253636816
+     -0.05113714002576085
+       0.2737234911893462
+ 3.63e+10    
+       0.2749183973712519
+     -0.05121556889747431
+       0.2782580393358309
+    -0.005677266284277574
+     -0.02276282582934494
+       0.2783994905237576
+    -0.003518823143940083
+    -0.005663327345581785
+      -0.0512848667961301
+        0.274363963648264
+ 3.64e+10    
+       0.2755595016055875
+     -0.05136350893740675
+       0.2789339712609731
+      -0.0057095611614537
+     -0.02284013159283331
+       0.2790752303251157
+    -0.003520452935284525
+    -0.005695625779220486
+       -0.051432725828362
+       0.2750036000791016
+ 3.65e+10    
+       0.2761997664060836
+     -0.05151158257264041
+       0.2796092794883655
+    -0.005741822650670644
+     -0.02291760920325166
+       0.2797503490448984
+    -0.003521852380979451
+    -0.005727891565820807
+     -0.05158071848136731
+        0.275642399183577
+ 3.66e+10    
+       0.2768391903173762
+      -0.0516597910550168
+       0.2802839611932982
+    -0.005774048775151868
+     -0.02299525947833602
+       0.2804248441610558
+      -0.0035230187911671
+    -0.005760122724799834
+      -0.0517288460994159
+        0.276280359668743
+ 3.67e+10    
+       0.2774777718913358
+       -0.051808135624043
+        0.280958013612233
+    -0.005806237565884421
+     -0.02307308322048807
+        0.281098713201012
+    -0.003523949490667645
+    -0.005792317283759759
+     -0.05187711001180015
+        0.276917480246925
+ 3.68e+10    
+       0.2781155096870346
+     -0.05195661750655214
+       0.2816314340428899
+    -0.005838387061652017
+     -0.02315108121704333
+       0.2817719537417909
+    -0.003524641819674173
+    -0.005824473278519683
+     -0.05202551153249547
+        0.277553759635651
+ 3.69e+10    
+       0.2787524022707108
+     -0.05210523791635784
+       0.2823042198442639
+    -0.005870495309064578
+     -0.02322925424052994
+       0.2824445634100897
+    -0.003525093134442081
+    -0.005856588753143523
+     -0.05217405195981958
+       0.2781891965575833
+ 3.7e+10     
+       0.2793884482157266
+     -0.05225399805390433
+       0.2829763684365749
+     -0.00590256036258437
+     -0.02330760304892014
+       0.2831165398822943
+    -0.003525300807972715
+    -0.005888661759963627
+     -0.05232273257608964
+       0.2788237897404464
+ 3.71e+10    
+       0.2800236461025229
+     -0.05240289910591138
+       0.2836478773011514
+    -0.005934580284548504
+     -0.02338612838587318
+       0.2837878808844483
+    -0.003525262230691443
+    -0.005920690359600463
+      -0.0524715546472784
+        0.279457537916954
+ 3.72e+10    
+        0.280657994518575
+     -0.05255194224501657
+       0.2843187439802509
+     -0.00596655314518865
+     -0.02346483098097068
+       0.2844585841921661
+    -0.003524974811119677
+    -0.005952672620978846
+     -0.05262051942266863
+       0.2800904398247327
+ 3.73e+10    
+       0.2812914920583374
+     -0.05270112862941227
+       0.2849889660768216
+    -0.005998477022647137
+     -0.02354371154994392
+       0.2851286476304976
+    -0.003524435976540947
+    -0.005984606621340078
+     -0.05276962813450577
+       0.2807224942062447
+ 3.74e+10    
+        0.281924137323192
+     -0.05285045940248058
+       0.2856585412542047
+    -0.006030350002990058
+     -0.02362277079489493
+       0.2857980690737539
+    -0.003523643173660891
+     -0.00601649044625051
+      -0.0529188819976527
+       0.2813536998087112
+ 3.75e+10    
+       0.2825559289213896
+      -0.0529999356924245
+       0.2863274672357803
+    -0.006062170180217388
+     -0.02370200940450888
+       0.2864668464452768
+    -0.003522593869260993
+    -0.006048322189606888
+     -0.05306828220924001
+       0.2819840553840287
+ 3.76e+10    
+       0.2831868654679897
+     -0.05314955861189723
+       0.2869957418045637
+    -0.006093935656269693
+     -0.02378142805426106
+       0.2871349777171724
+    -0.003521285550846119
+    -0.006080099953637936
+       -0.053217829948319
+       0.2826135596886895
+ 3.77e+10    
+       0.2838169455847959
+     -0.05329932925762827
+       0.2876633628027458
+    -0.006125644541032649
+     -0.02386102740661598
+       0.2878024609100013
+    -0.003519715727285494
+    -0.006111821848902606
+     -0.05336752637551327
+       0.2832422114836972
+ 3.78e+10    
+       0.2844461679002906
+     -0.05344924871004854
+       0.2883303281311884
+    -0.006157294952337966
+     -0.02394080811122084
+       0.2884692940924282
+    -0.003517881929447268
+    -0.006143485994285464
+     -0.05351737263267067
+       0.2838700095344819
+ 3.79e+10    
+       0.2850745310495664
+     -0.05359931803291397
+       0.2889966357488718
+    -0.006188885015961811
+     -0.02402077080509216
+        0.289135475380833
+    -0.003515781710826432
+    -0.006175090516988446
+     -0.05366736984251549
+       0.2844969526108136
+ 3.8e+10     
+       0.2857020336742517
+     -0.05374953827292712
+       0.2896622836723005
+    -0.006220412865620504
+      -0.0241009161127972
+       0.2898010029388863
+    -0.003513412648166047
+    -0.006206633552519646
+     -0.05381751910830175
+       0.2851230394867152
+ 3.81e+10    
+       0.2863286744224398
+       -0.053899910459359
+       0.2903272699748622
+     -0.00625187664296367
+     -0.02418124464662877
+       0.2904658749770914
+    -0.003510772342071605
+    -0.006238113244679596
+     -0.05396782151346719
+       0.2857482689403743
+ 3.82e+10    
+        0.286954451948609
+     -0.05405043560366942
+       0.2909915927861523
+    -0.006283274497564474
+     -0.02426175700677492
+       0.2911300897522892
+    -0.003507858417618486
+    -0.006269527745543868
+     -0.05411827812128769
+       0.2863726397540514
+ 3.83e+10    
+        0.287579364913547
+     -0.05420111469912875
+       0.2916552502912597
+    -0.006314604586907678
+      -0.0243424537814837
+        0.291793645567135
+    -0.003504668524952437
+    -0.006300875215443532
+     -0.05426888997453401
+       0.2869961507139914
+ 3.84e+10    
+       0.2882034119842672
+     -0.05435194872043809
+       0.2923182407300151
+    -0.006345865076374723
+     -0.02442333554722212
+       0.2924565407695451
+    -0.003501200339883007
+    -0.006332153822942466
+     -0.05441965809512962
+       0.2876188006103305
+ 3.85e+10    
+       0.2888265918339271
+     -0.05450293862335149
+       0.2929805623962081
+    -0.006377054139226972
+     -0.02450440286883103
+       0.2931187737521121
+    -0.003497451564469606
+    -0.006363361744812241
+     -0.05457058348380991
+        0.288240588237003
+ 3.86e+10    
+       0.2894489031417408
+     -0.05465408534429821
+       0.2936422136367737
+    -0.006408169956586117
+     -0.02458565629967479
+       0.2937803429514966
+    -0.003493419927600422
+    -0.006394497166004501
+     -0.05472166711978386
+       0.2888615123916483
+ 3.87e+10    
+       0.2900703445928958
+     -0.05480538980000664
+       0.2943031928509476
+    -0.006439210717412822
+     -0.02466709638178684
+       0.2944412468477925
+    -0.003489103185563913
+    -0.006425558279620519
+     -0.05487290996039853
+       0.2894815718755172
+ 3.88e+10    
+       0.2906909148784602
+     -0.05495685288712981
+       0.2949634984893958
+    -0.006470174618482304
+     -0.02474872364601134
+       0.2951014839638658
+    -0.003484499122612846
+    -0.006456543286878736
+     -0.05502431294080387
+       0.2901007654933752
+ 3.89e+10    
+       0.2913106126952947
+     -0.05510847548187194
+       0.2956231290533186
+    -0.006501059864358699
+     -0.02483053861214052
+       0.2957610528646785
+    -0.003479605551520683
+    -0.006487450397079663
+     -0.05517587697362306
+       0.2907190920534075
+ 3.9e+10     
+       0.2919294367459603
+     -0.05526025843961861
+       0.2962820830935314
+    -0.006531864667366638
+     -0.02491254178904833
+       0.2964199521565807
+     -0.00347442031413042
+    -0.006518277827568949
+     -0.05532760294862312
+       0.2913365503671234
+ 3.91e+10    
+       0.2925473857386235
+     -0.05541220259456793
+       0.2969403592095234
+     -0.00656258724756094
+     -0.02499473367482087
+       0.2970781804865933
+    -0.003468941281895664
+    -0.006549023803697684
+     -0.05547949173239056
+       0.2919531392492597
+ 3.92e+10    
+        0.293164458386963
+     -0.05556430875936499
+       0.2975979560484967
+    -0.006593225832694482
+     -0.02507711475688318
+        0.297735736541666
+    -0.003463166356413814
+     -0.00657968655878113
+     -0.05563154416800832
+       0.2925688575176812
+ 3.93e+10    
+       0.2937806534100719
+     -0.05571657772473979
+        0.298254872304388
+    -0.006623778658183779
+     -0.02515968551212317
+       0.2983926190479212
+    -0.003457093469951461
+    -0.006610264334055113
+     -0.05578376107473784
+       0.2931837039932851
+ 3.94e+10    
+       0.2943959695323619
+     -0.05586901025914752
+       0.2989111067168726
+    -0.006654243967073133
+     -0.02524244640701252
+       0.2990488267698818
+    -0.003450720585961559
+    -0.006640755378630696
+     -0.05593614324770418
+       0.2937976774999034
+ 3.95e+10    
+       0.2950104054834631
+     -0.05602160710841316
+       0.2995666580703547
+    -0.006684620009996487
+     -0.02532539789772477
+       0.2997043585096834
+    -0.003444045699592842
+    -0.006671157949446734
+     -0.05608869145758422
+       0.2944107768642032
+ 3.96e+10    
+        0.295623959998127
+     -0.05617436899537955
+       0.3002215251929449
+    -0.006714905045137685
+     -0.02540854043025133
+       0.3003592131062786
+    -0.003437066838190837
+    -0.006701470311220793
+     -0.05624140645030055
+         0.29502300091559
+ 3.97e+10    
+       0.2962366318161234
+     -0.05632729661955935
+       0.3008757069554233
+    -0.006745097338189295
+     -0.02549187444051434
+       0.3010133894346218
+    -0.003429782061790643
+    -0.006731690736398156
+     -0.05639428894671752
+       0.2956343484861085
+ 3.98e+10    
+       0.2968484196821411
+     -0.05648039065679136
+       0.3015292022701973
+    -0.006775195162309219
+     -0.02557540035447815
+       0.3016668864048475
+    -0.003422189463601587
+     -0.00676181750509941
+      -0.0565473396423428
+       0.2962448184103439
+ 3.99e+10    
+       0.2974593223456843
+     -0.05663365175890174
+       0.3021820100902448
+    -0.006805196798076117
+     -0.02565911858825828
+       0.3023197029614403
+    -0.003414287170483211
+    -0.006791848905066164
+     -0.05670055920703349
+        0.296854409525324
+ 4e+10       
+       0.2980693385609714
+     -0.05678708055336922
+       0.3028341294080551
+    -0.006835100533443137
+     -0.02574302954822888
+       0.3029718380823944
+     -0.00340607334341298
+     -0.00682178323160545
+     -0.05685394828470679
+       0.2974631206704215
+ 4.01e+10    
+       0.2986784670868313
+      -0.0569406776429958
+       0.3034855592545604
+     -0.00686490466369008
+     -0.02582713363112829
+       0.3036232907783661
+    -0.003397546177945411
+    -0.006851618787532286
+     -0.05700750749305477
+       0.2980709506872534
+ 4.02e+10    
+       0.2992867066865987
+     -0.05709444360558272
+       0.3041362986980649
+    -0.006894607491374181
+     -0.02591143122416303
+       0.3042740600918198
+    -0.003388703904662432
+    -0.006881353883111509
+     -0.05716123742326522
+       0.2986778984195865
+ 4.03e+10    
+       0.2998940561280116
+     -0.05724837899361089
+       0.3047863468431673
+    -0.006924207326279496
+     -0.02599592270511053
+       0.3049241450961683
+    -0.003379544789615229
+    -0.006910986835997324
+     -0.05731513863974624
+       0.2992839627132355
+ 4.04e+10    
+       0.3005005141831054
+     -0.05740248433392786
+        0.305435702829685
+    -0.006953702485364964
+     -0.02608060844242076
+       0.3055735448949117
+    -0.003370067134757228
+     -0.00694051597117238
+     -0.05746921167985837
+       0.2998891424159692
+ 4.05e+10    
+       0.3011060796281082
+     -0.05755676012744004
+       0.3060843658315735
+    -0.006983091292710961
+     -0.02616548879531646
+       0.3062222586207673
+    -0.003360269278368143
+    -0.006969939620885299
+     -0.05762345705364892
+       0.3004934363774107
+ 4.06e+10    
+       0.3017107512433367
+     -0.05771120684881059
+       0.3067323350558469
+    -0.007012372079465054
+     -0.02625056411389256
+       0.3068702854348032
+      -0.0033501495954693
+    -0.006999256124586933
+     -0.05777787524359517
+       0.3010968434489425
+ 4.07e+10    
+       0.3023145278130892
+     -0.05786582494616359
+       0.3073796097415014
+    -0.007041543183785958
+     -0.02633583473921467
+       0.3075176245255654
+    -0.003339706498229825
+    -0.007028463828865598
+     -0.05793246670435058
+       0.3016993624836089
+ 4.08e+10    
+        0.302917408125543
+     -0.05802061484079503
+       0.3080261891584367
+    -0.007070602950786922
+     -0.02642130100341725
+       0.3081642751082059
+    -0.003328938436363821
+    -0.007057561087381391
+     -0.05808723186249781
+       0.3023009923360201
+ 4.09e+10    
+       0.3035193909726463
+     -0.05817557692688828
+       0.3086720726063829
+    -0.007099549732477714
+     -0.02650696322980037
+       0.3088102364236116
+    -0.003317843897518406
+    -0.007086546260799442
+     -0.05824217111630841
+       0.3029017318622586
+ 4.1e+10     
+       0.3041204751500145
+      -0.0583307115712386
+       0.3093172594138316
+    -0.007128381887705611
+     -0.02659282173292665
+        0.309455507737532
+     -0.00330642140765258
+    -0.007115417716722104
+     -0.05839728483550653
+       0.3035015799197822
+ 4.11e+10    
+        0.304720659456825
+      -0.0584860191129821
+       0.3099617489369689
+    -0.007157097782095298
+      -0.0266788768187176
+       0.3101000883397103
+    -0.003294669531406898
+    -0.007144173829620321
+     -0.05855257336104086
+       0.3041005353673308
+ 4.12e+10    
+       0.3053199426957118
+     -0.05864149986333279
+       0.3106055405586184
+     -0.00718569578798819
+     -0.02676512878454974
+       0.3107439775430161
+    -0.003282586872463672
+    -0.007172812980764378
+     -0.05870803700486195
+       0.3046985970648357
+ 4.13e+10    
+        0.305918323672662
+     -0.05879715410532596
+       0.3112486336871856
+    -0.007214174284380263
+     -0.02685157791935028
+       0.3113871746825787
+    -0.003270172073897979
+    -0.007201333558153576
+     -0.05886367604970402
+       0.3052957638733218
+ 4.14e+10    
+       0.3065158011969094
+     -0.05895298209356856
+       0.3118910277556114
+    -0.007242531656859668
+      -0.0269382245036929
+       0.3120296791149287
+    -0.003257423818519015
+    -0.007229733956445362
+     -0.05901949074887711
+       0.3058920346548205
+ 4.15e+10    
+       0.3071123740808319
+     -0.05910898405399638
+        0.312532722220336
+    -0.007270766297543053
+     -0.02702506880989338
+       0.3126714902171374
+    -0.003244340829202203
+    -0.007258012576883837
+     -0.05917548132606133
+       0.3064874082722753
+ 4.16e+10    
+       0.3077080411398477
+      -0.0592651601836398
+       0.3131737165602652
+    -0.007298876605011429
+     -0.02711211110210545
+       0.3133126073859685
+    -0.003230921869211503
+    -0.007286167827227423
+      -0.0593316479751114
+        0.307081883589454
+ 4.17e+10    
+        0.308302801192312
+     -0.05942151065039491
+        0.313814010275751
+    -0.007326860984245076
+     -0.02719935163641653
+       0.3139530300370276
+    -0.003217165742512251
+    -0.007314198121676288
+     -0.05948799085986486
+       0.3076754594708581
+ 4.18e+10    
+       0.3088966530594138
+     -0.05957803559280318
+         0.31445360288758
+    -0.007354717846558152
+     -0.02728679066094371
+       0.3145927576039227
+    -0.003203071294074291
+    -0.007342101880798922
+     -0.05964451011395894
+       0.3082681347816349
+ 4.19e+10    
+       0.3094895955650757
+     -0.05973473511983892
+       0.3150924939359717
+    -0.007382445609532245
+     -0.02737442841593037
+       0.3152317895374291
+     -0.00318863741016533
+    -0.007369877531458553
+     -0.05980120584065374
+       0.3088599083874901
+ 4.2e+10     
+       0.3100816275358487
+     -0.05989160931070256
+       0.3157306829795878
+    -0.007410042696949703
+     -0.02746226513384226
+       0.3158701253046605
+    -0.003173863018634569
+    -0.007397523506739003
+     -0.05995807811266133
+       0.3094507791546016
+ 4.21e+10    
+       0.3106727478008158
+     -0.06004865821462405
+       0.3163681695945523
+     -0.00743750753872629
+     -0.02755030103946504
+       0.3165077643882489
+    -0.003158747089186494
+    -0.007425038245869998
+      -0.0601151269719828
+       0.3100407459495331
+ 4.22e+10    
+       0.3112629551914893
+     -0.06020588185067152
+       0.3170049533734844
+    -0.007464838570843341
+     -0.02763853635000121
+       0.3171447062855319
+    -0.003143288633644712
+    -0.007452420194152692
+     -0.06027235242975252
+       0.3106298076391523
+ 4.23e+10    
+       0.3118522485417113
+     -0.06036328020756918
+       0.3176410339245418
+     -0.00749203423527952
+     -0.02772697127516816
+       0.3177809505077464
+    -0.003127486706205967
+     -0.00747966780288419
+     -0.06042975446608755
+       0.3112179630905446
+ 4.24e+10    
+       0.3124406266875563
+     -0.06052085324352289
+       0.3182764108704793
+    -0.007519092979942345
+     -0.02781560601729668
+       0.3184164965792339
+    -0.003111340403684013
+    -0.007506779529282475
+     -0.06058733302994678
+       0.3118052111709336
+ 4.25e+10    
+       0.3130280884672328
+     -0.06067860088605233
+       0.3189110838477156
+    -0.007546013258598894
+     -0.02790444077142958
+       0.3190513440366515
+    -0.003094848865743662
+    -0.007533753836410834
+     -0.06074508803899448
+       0.3123915507475998
+ 4.26e+10    
+       0.3136146327209862
+     -0.06083652303183281
+       0.3195450525054186
+    -0.007572793530806957
+     -0.02799347572542131
+       0.3196854924281944
+    -0.003078011275124477
+    -0.007560589193102128
+     -0.06090301937947361
+       0.3129769806878004
+ 4.27e+10    
+       0.3142002582910052
+     -0.06099461954654421
+       0.3201783165046011
+     -0.00759943226184502
+     -0.02808271106003821
+       0.3203189413128273
+    -0.003060826857854652
+    -0.007587284073883205
+     -0.06106112690608344
+       0.3135614998586899
+ 4.28e+10    
+        0.314784964021322
+     -0.06115289026472713
+       0.3208108755172307
+    -0.007625927922642843
+     -0.02817214694905902
+       0.3209516902595243
+    -0.003043294883454468
+    -0.007613836958898919
+     -0.06121941044186756
+       0.3141451071272468
+ 4.29e+10    
+       0.3153687487577232
+     -0.06131133498964807
+       0.3214427292253546
+    -0.007652278989711361
+     -0.02826178355937651
+       0.3215837388465225
+    -0.003025414665129667
+    -0.007640246333836394
+     -0.06137786977810644
+       0.3147278013601939
+ 4.3e+10     
+       0.3159516113476546
+      -0.0614699534931725
+       0.3220738773202375
+    -0.007678483945072698
+     -0.02835162105109924
+       0.3222150866605814
+    -0.003007185559954515
+     -0.00766651068984934
+     -0.06153650467421841
+       0.3153095814239253
+ 4.31e+10    
+       0.3165335506401286
+     -0.06162874551564575
+       0.3227043195015171
+    -0.007704541276189882
+     -0.02844165957765494
+       0.3228457332962555
+    -0.002988606969044659
+    -0.007692628523482174
+     -0.06169531485766853
+       0.3158904461844351
+ 4.32e+10    
+       0.3171145654856353
+      -0.0617877107657814
+       0.3233340554763675
+    -0.007730449475896626
+     -0.02853189928589353
+       0.3234756783551803
+    -0.002969678337719547
+    -0.007718598336594426
+      -0.0618543000238837
+       0.3164703945072416
+ 4.33e+10    
+        0.317694654736052
+     -0.06194684892055908
+       0.3239630849586875
+    -0.007756207042327261
+     -0.02862234031619139
+       0.3241049214453619
+    -0.002950399155654532
+     -0.00774441863628548
+     -0.06201345983617544
+       0.3170494252573211
+ 4.34e+10    
+       0.3182738172445537
+     -0.06210615962512882
+       0.3245914076682954
+    -0.007781812478846164
+     -0.02871298280255682
+       0.3247334621804867
+    -0.002930768957022629
+    -0.007770087934819045
+     -0.06217279392567036
+       0.3176275372990369
+ 4.35e+10    
+       0.3188520518655277
+     -0.06226564249272518
+       0.3252190233301429
+    -0.007807264293977933
+     -0.02880382687273523
+       0.3253613001792356
+    -0.002910787320625692
+    -0.007795604749548339
+     -0.06233230189124762
+       0.3182047294960723
+ 4.36e+10    
+       0.3194293574544859
+     -0.06242529710458743
+       0.3258459316735439
+     -0.00783256100133721
+     -0.02889487264831606
+       0.3259884350646154
+    -0.002890453870015335
+    -0.007820967602841115
+     -0.06249198329948469
+       0.3187810007113651
+ 4.37e+10    
+       0.3200057328679801
+     -0.06258512300988969
+       0.3264721324314178
+    -0.007857701119558648
+      -0.0289861202448397
+        0.326614866463297
+    -0.002869768273603068
+    -0.007846175022005391
+     -0.06265183768460858
+        0.319356349807042
+ 4.38e+10    
+       0.3205811769635211
+     -0.06274511972567834
+       0.3270976253395497
+    -0.007882683172227315
+      -0.0290775697719057
+       0.3272405940049671
+    -0.002848730244760266
+    -0.007871225539215123
+     -0.06281186454845654
+       0.3199307756443573
+ 4.39e+10    
+       0.3211556885994913
+     -0.06290528673681696
+       0.3277224101358653
+     -0.00790750568780909
+     -0.02916922133328138
+       0.3278656173216948
+    -0.002827339541907209
+    -0.007896117691436581
+      -0.0629720633604431
+       0.3205042770836311
+ 4.4e+10     
+        0.321729266635069
+     -0.06306562349594125
+       0.3283464865597214
+    -0.007932167199581503
+     -0.02926107502701152
+       0.3284899360473069
+    -0.002805595968591823
+    -0.007920850020354911
+     -0.06313243355753455
+       0.3210768529841876
+ 4.41e+10    
+       0.3223019099301462
+     -0.06322612942341883
+       0.3289698543512115
+    -0.007956666245564577
+     -0.02935313094552821
+       0.3291135498167755
+    -0.002783499373557694
+    -0.007945421072301222
+      -0.0632929745442313
+       0.3216485022042995
+ 4.42e+10    
+       0.3228736173452508
+     -0.06338680390732136
+       0.3295925132504902
+    -0.007981001368452229
+     -0.02944538917576225
+       0.3297364582656198
+    -0.002761049650801401
+     -0.00796982939818025
+     -0.06345368569255724
+       0.3222192236011311
+ 4.43e+10    
+       0.3234443877414693
+     -0.06354764630340001
+       0.3302144629971068
+    -0.008005171115544054
+      -0.0295378497992544
+       0.3303586610293194
+    -0.002738246739619364
+     -0.00799407355339829
+     -0.06361456634205609
+       0.3227890160306807
+ 4.44e+10    
+       0.3240142199803731
+     -0.06370865593507279
+       0.3308357033293624
+    -0.008029174038677336
+      -0.0296305128922679
+       0.3309801577427381
+     -0.00271509062464385
+    -0.008018152097792004
+     -0.06377561579979682
+       0.3233578783477315
+ 4.45e+10    
+       0.3245831129239439
+     -0.06386983209341829
+       0.3314562339836766
+     -0.00805300869415952
+     -0.02972337852590168
+       0.3316009480395646
+    -0.002691581335868341
+    -0.008042063595557297
+     -0.06393683334038405
+       0.3239258094057949
+ 4.46e+10    
+          0.3251510654345
+     -0.06403117403717651
+       0.3320760546939722
+    -0.008076673642701256
+     -0.02981644676620364
+       0.3322210315517606
+     -0.00266771894866231
+    -0.008065806615179461
+     -0.06409821820597827
+       0.3244928080570658
+ 4.47e+10    
+        0.325718076374628
+      -0.0641926809927601
+       0.3326951651910772
+    -0.008100167449349939
+     -0.02990971767428548
+       0.3328404079090233
+     -0.00264350358377504
+    -0.008089379729363477
+     -0.06425976960632103
+       0.3250588731523703
+ 4.48e+10    
+       0.3262841446071101
+     -0.06435435215427017
+       0.3333135652021365
+     -0.00812348868342358
+     -0.03000319130643736
+        0.333459076738263
+    -0.002618935407328939
+    -0.008112781514964989
+     -0.06442148671876978
+       0.3256240035411204
+ 4.49e+10    
+       0.3268492689948613
+     -0.06451618668352427
+       0.3339312544500476
+    -0.008146635918445458
+     -0.03009686771424369
+       0.3340770376630888
+    -0.002594014630801991
+    -0.008136010552922429
+     -0.06458336868833831
+       0.3261881980712704
+ 4.5e+10     
+        0.327413448400857
+     -0.06467818371008761
+       0.3345482326529025
+    -0.008169607732079219
+     -0.03019074694469918
+       0.3346942903033094
+    -0.002568741510999458
+    -0.008159065428189199
+     -0.06474541462774527
+       0.3267514555892718
+ 4.51e+10    
+       0.3279766816880738
+     -0.06484034233131598
+       0.3351644995234521
+      -0.0081924027060648
+     -0.03028482904032566
+       0.3353108342744464
+    -0.002543116350014807
+    -0.008181944729667212
+     -0.06490762361747018
+       0.3273137749400329
+ 4.52e+10    
+       0.3285389677194223
+     -0.06500266161240387
+       0.3357800547685827
+    -0.008215019426154647
+     -0.03037911403928942
+       0.3359266691872579
+    -0.002517139495179941
+    -0.008204647050140871
+     -0.06506999470581618
+       0.3278751549668795
+ 4.53e+10    
+       0.3291003053576894
+     -0.06516514058644228
+       0.3363948980888066
+    -0.008237456482051009
+     -0.03047360197551892
+       0.3365417946472782
+     -0.00249081133900453
+     -0.00822717098621195
+     -0.06523252690898021
+       0.3284355945115164
+ 4.54e+10    
+       0.3296606934654751
+     -0.06532777825448259
+       0.3370090291777701
+    -0.008259712467343725
+     -0.03056829287882324
+       0.3371562102543648
+    -0.002464132319104701
+    -0.008249515138235427
+     -0.06539521921113081
+       0.3289950924139929
+ 4.55e+10    
+       0.3302201309051372
+     -0.06549057358560964
+       0.3376224477217755
+    -0.008281785979448774
+     -0.03066318677501083
+       0.3377699156022644
+    -0.002437102918120825
+    -0.008271678110255911
+     -0.06555807056449268
+       0.3295536475126666
+ 4.56e+10    
+       0.3307786165387321
+     -0.06565352551702111
+       0.3382351533993159
+    -0.008303675619547713
+     -0.03075828368600851
+       0.3383829102781828
+    -0.002409723663624551
+    -0.008293658509945394
+     -0.06572107988943851
+       0.3301112586441722
+ 4.57e+10    
+        0.331336149227963
+      -0.0658166329541158
+       0.3388471458806287
+    -0.008325379992527821
+     -0.03085358362998139
+       0.3389951938623757
+    -0.002381995128015122
+    -0.008315454948541339
+     -0.06588424607458809
+         0.33066792464339
+ 4.58e+10    
+       0.3318927278341242
+     -0.06597989477058855
+       0.3394584248272587
+    -0.008346897706922896
+     -0.03094908662145283
+       0.3396067659277451
+     -0.00235391792840489
+    -0.008337066040786314
+     -0.06604756797691501
+       0.3312236443434204
+ 4.59e+10    
+       0.3324483512180518
+     -0.06614330980853322
+       0.3400689898916406
+    -0.008368227374855396
+     -0.03104479267142466
+        0.340217626039451
+    -0.002325492726494022
+    -0.008358490404868281
+     -0.06621104442185916
+       0.3317784165755534
+ 4.6e+10     
+       0.3330030182400728
+     -0.06630687687855323
+       0.3406788407166913
+    -0.008389367611978936
+     -0.03114070178749785
+       0.3408277737545336
+    -0.002296720228434428
+    -0.008379726662361742
+     -0.06637467420344793
+       0.3323322401692456
+ 4.61e+10    
+       0.3335567277599581
+     -0.06647059475987903
+        0.341287976935419
+    -0.008410317037422109
+     -0.03123681397399378
+       0.3414372086215496
+    -0.002267601184683088
+    -0.008400773438170236
+     -0.06653845608442313
+       0.3328851139520962
+ 4.62e+10    
+       0.3341094786368751
+     -0.06663446220049338
+       0.3418963981705457
+     -0.00843107427373279
+     -0.03133312923207517
+        0.342045930180217
+    -0.002238136389844447
+    -0.008421629360469715
+     -0.06670238879637595
+       0.3334370367498281
+ 4.63e+10    
+       0.3346612697293455
+     -0.06679847791726436
+       0.3425041040341427
+    -0.008451637946823989
+     -0.03142964755986775
+       0.3426539379610747
+    -0.002208326682502225
+    -0.008442293060652938
+     -0.06686647103988805
+       0.3339880073862654
+ 4.64e+10    
+       0.3352120998952015
+     -0.06696264059608524
+         0.34311109412728
+     -0.00847200668592004
+     -0.03152636895258187
+       0.3432612314851528
+    -0.002178172945040442
+    -0.008462763173274976
+     -0.06703070148468038
+       0.3345380246833196
+ 4.65e+10    
+       0.3357619679915444
+     -0.06712694889202124
+       0.3437173680396906
+    -0.008492179123504435
+     -0.03162329340263446
+       0.3438678102636537
+    -0.002147676103453765
+    -0.008483038335999856
+     -0.06719507876976874
+       0.3350870874609725
+ 4.66e+10    
+       0.3363108728747086
+     -0.06729140142946508
+       0.3443229253494455
+    -0.008512153895268099
+     -0.03172042089977077
+       0.3444736737976457
+    -0.002116837127147273
+     -0.00850311718954843
+     -0.06735960150362542
+       0.3356351945372623
+ 4.67e+10    
+       0.3368588134002198
+     -0.06745599680229751
+        0.344927765622644
+    -0.008531929640059093
+     -0.03181775143118688
+       0.3450788215777664
+    -0.002085657028725397
+    -0.008522998377647003
+     -0.06752426826434874
+       0.3361823447282734
+ 4.68e+10    
+       0.3374057884227659
+     -0.06762073357405733
+       0.3455318884131172
+    -0.008551504999833408
+     -0.03191528498165157
+       0.3456832530839403
+    -0.002054136863770417
+    -0.008542680546977776
+     -0.06768907759983958
+       0.3367285368481276
+ 4.69e+10    
+       0.3379517967961584
+     -0.06778561027811704
+       0.3461352932621423
+    -0.008570878619606493
+     -0.03201302153362871
+       0.3462869677851045
+    -0.002022277730610228
+     -0.00856216234712971
+     -0.06785402802798307
+       0.3372737697089743
+ 4.7e+10     
+       0.3384968373733043
+     -0.06795062541786548
+       0.3467379796981703
+    -0.008590049147406414
+     -0.03211096106739939
+       0.3468899651389472
+    -0.001990080770075596
+    -0.008581442430551301
+     -0.06801911803683908
+       0.3378180421209874
+ 4.71e+10    
+       0.3390409090061743
+     -0.06811577746689844
+       0.3473399472365675
+    -0.008609015234227621
+     -0.03220910356118428
+       0.3474922445916566
+    -0.001957547165246913
+    -0.008600519452504028
+     -0.06818434608483823
+       0.3383613528923612
+ 4.72e+10    
+       0.3395840105457776
+     -0.06828106486921606
+        0.347941195379369
+    -0.008627775533986319
+     -0.03230744899126588
+       0.3480938055776815
+    -0.001924678141190314
+    -0.008619392071017373
+     -0.06834971060098473
+       0.3389037008293083
+ 4.73e+10    
+       0.3401261408421341
+     -0.06844648603942573
+       0.3485417236150412
+    -0.008646328703476772
+     -0.03240599733211032
+       0.3486946475195002
+    -0.001891474964683456
+    -0.008638058946845047
+     -0.06851520998506616
+       0.3394450847360609
+ 4.74e+10    
+       0.3406672987442524
+     -0.06861203936295449
+       0.3491415314182623
+    -0.008664673402328885
+     -0.03250474855648983
+       0.3492947698274035
+    -0.001857938943930761
+    -0.008656518743422209
+     -0.06868084260786964
+        0.339985503414873
+ 4.75e+10    
+       0.3412074831001061
+     -0.06877772319626549
+       0.3497406182497084
+    -0.008682808292966906
+     -0.03260370263560418
+       0.3498941718992856
+    -0.001824071428268363
+    -0.008674770126824449
+     -0.06884660681140475
+       0.3405249556660263
+ 4.76e+10    
+       0.3417466927566153
+     -0.06894353586708307
+       0.3503389835558566
+     -0.00870073204056945
+     -0.03270285953920278
+       0.3504928531204455
+    -0.001789873807858533
+    -0.008692811765727747
+     -0.06901250090913272
+       0.3410634402878351
+ 4.77e+10    
+       0.3422849265596289
+     -0.06910947567462448
+       0.3509366267687936
+    -0.008718443313030807
+     -0.03280221923570573
+       0.3510908128634008
+    -0.001755347513374024
+    -0.008710642331369626
+     -0.06917852318620241
+       0.3416009560766556
+ 4.78e+10    
+        0.342822183353907
+     -0.06927554088983667
+       0.3515335473060421
+    -0.008735940780923417
+     -0.03290178169232551
+       0.3516880504877093
+    -0.001720494015671852
+    -0.008728260497512146
+     -0.06934467189969253
+       0.3421375018268978
+ 4.79e+10    
+       0.3433584619831094
+     -0.06944172975564213
+       0.3521297445703939
+    -0.008753223117461646
+     -0.03300154687518777
+       0.3522845653398016
+    -0.001685314825457167
+    -0.008745664940405627
+     -0.06951094527886109
+       0.3426730763310384
+ 4.8e+10     
+       0.3438937612897808
+     -0.06960804048718905
+       0.3527252179497561
+    -0.008770288998466871
+     -0.03310151474945217
+       0.3528803567528238
+    -0.001649811492936688
+    -0.008762854338754313
+     -0.06967734152539928
+       0.3432076783796342
+ 4.81e+10    
+       0.3444280801153431
+     -0.06977447127210962
+       0.3533199668170056
+    -0.008787137102333909
+     -0.03320168527943264
+       0.3534754240464883
+    -0.001613985607462173
+    -0.008779827373682828
+     -0.06984385881369352
+       0.3437413067613393
+ 4.82e+10    
+        0.344961417300088
+     -0.06994102027078469
+       0.3539139905298587
+    -0.008803766109998652
+     -0.03330205842871767
+        0.354069766526938
+     -0.00157783879716377
+     -0.00879658272870453
+      -0.0700104952910941
+       0.3442739602629278
+ 4.83e+10    
+       0.3454937716831672
+     -0.07010768561661275
+       0.3545072884307456
+    -0.008820174704907252
+     -0.03340263416028974
+       0.3546633834866159
+    -0.001541372728573317
+    -0.008813119089690943
+     -0.07017724907818788
+       0.3448056376693098
+ 4.84e+10    
+       0.3460251421025937
+     -0.07027446541628911
+       0.3550998598466996
+    -0.008836361572986376
+     -0.03350341243664486
+        0.355256274204146
+    -0.001504589106237813
+    -0.008829435144842683
+     -0.07034411826907941
+       0.3453363377635593
+ 4.85e+10    
+       0.3465555273952357
+     -0.07044135775008795
+        0.355691704089256
+     -0.00885232540261505
+     -0.03360439321991134
+       0.3558484379442243
+    -0.001467489672322795
+    -0.008845529584661855
+      -0.0705111009316768
+       0.3458660593269364
+ 4.86e+10    
+         0.34708492639682
+     -0.07060836067215229
+       0.3562828204543562
+    -0.008868064884597807
+     -0.03370557647196817
+       0.3564398739575165
+    -0.001430076206206161
+    -0.008861401101925657
+     -0.07067819510798529
+       0.3463948011389184
+ 4.87e+10    
+        0.347613337941933
+     -0.07077547221079039
+       0.3568732082222698
+     -0.00888357871213909
+      -0.0338069621545629
+       0.3570305814805679
+    -0.001392350524061884
+    -0.008877048391661837
+     -0.07084539881440484
+       0.3469225619772267
+ 4.88e+10    
+        0.348140760864024
+     -0.07094269036877715
+       0.3574628666575177
+    -0.008898865580819247
+     -0.03390855022942932
+       0.3576205597357196
+    -0.001354314478434416
+    -0.008892470151124963
+     -0.07101271004203577
+       0.3474493406178596
+ 4.89e+10    
+       0.3486671939954129
+     -0.07111001312366297
+       0.3580517950088108
+    -0.008913924188571822
+     -0.03401034065840391
+       0.3582098079310336
+    -0.001315969957803087
+    -0.008907665079774828
+      -0.0711801267569887
+       0.3479751358351266
+ 4.9e+10     
+       0.3491926361673007
+     -0.07127743842808838
+       0.3586399925089973
+    -0.008928753235662213
+     -0.03411233340354261
+       0.3587983252602295
+    -0.001277318886137287
+    -0.008922631879255905
+     -0.07134764690070254
+       0.3484999464016862
+ 4.91e+10    
+       0.3497170862097758
+       -0.071444964210104
+       0.3592274583750147
+    -0.008943351424667855
+     -0.03421452842723656
+        0.359386110902626
+    -0.001238363222441848
+    -0.008937369253378119
+     -0.07151526839026588
+       0.3490237710885808
+ 4.92e+10    
+       0.3502405429518305
+     -0.07161258837349702
+       0.3598141918078567
+    -0.008957717460459791
+     -0.03431692569232685
+       0.3599731640230932
+    -0.001199104960293356
+    -0.008951875908099585
+     -0.07168298911874647
+       0.3495466086652808
+ 4.93e+10    
+       0.3507630052213745
+     -0.07178030879812397
+       0.3604001919925442
+    -0.008971850050185526
+     -0.03441952516221915
+       0.3605594837720121
+    -0.001159546127366819
+    -0.008966150551510387
+     -0.07185080695552561
+        0.350068457899726
+ 4.94e+10    
+       0.3512844718452526
+     -0.07194812334024919
+       0.3609854580981091
+    -0.008985747903253632
+     -0.03452232680099823
+       0.3611450692852431
+    -0.001119688784953338
+    -0.008980191893817952
+     -0.07201871974663791
+       0.3505893175583699
+ 4.95e+10    
+       0.3518049416492627
+     -0.07211602983288865
+       0.3615699892775827
+    -0.008999409731319479
+     -0.03462533057354005
+       0.3617299196841013
+    -0.001079535027468477
+    -0.008993998647334108
+     -0.07218672531511759
+        0.351109186406228
+ 4.96e+10    
+       0.3523244134581782
+     -0.07228402608615983
+        0.362153784667996
+    -0.009012834248272558
+     -0.03472853644562532
+       0.3623140340753413
+    -0.001039086981951621
+    -0.009007569526463177
+     -0.07235482146135087
+       0.3516280632069272
+ 4.97e+10    
+       0.3528428860957723
+     -0.07245210988763823
+       0.3627368433903844
+    -0.009026020170225369
+     -0.03483194438405052
+       0.3628974115511497
+    -0.000998346807556331
+    -0.009020903247692051
+      -0.0725230059634325
+       0.3521459467227571
+ 4.98e+10    
+       0.3533603583848421
+      -0.0726202790027187
+       0.3633191645498069
+    -0.009038966215503487
+     -0.03493555435673949
+       0.3634800511891433
+   -0.0009573166950317632
+    -0.009033998529581474
+     -0.07269127657752938
+       0.3526628357147222
+ 4.99e+10    
+       0.3538768291472371
+     -0.07278853117498159
+       0.3639007472353643
+    -0.009051671104637362
+     -0.03503936633285323
+       0.3640619520523766
+   -0.0009159988661954009
+    -0.009046854092758785
+     -0.07285963103824897
+        0.353178728942602
+ 5e+10       
+       0.3543922972038894
+     -0.07295686412656735
+       0.3644815905202333
+    -0.009064133560355282
+     -0.03514338028290001
+       0.3646431131893575
+   -0.0008743955733969623
+    -0.009059468659912289
+     -0.07302806705901398
+        0.353693625165005
+ 5.01e+10    
+       0.3549067613748469
+      -0.0731252755585534
+       0.3650616934617043
+    -0.009076352307578216
+     -0.03524759617884347
+        0.365223533634069
+    -0.000832509098973771
+      -0.0090718409557871
+     -0.07319658233244217
+       0.3542075231394325
+ 5.02e+10    
+       0.3554202204793054
+     -0.07329376315133868
+       0.3656410551012254
+    -0.009088326073415734
+     -0.03535201399421103
+       0.3658032124059977
+   -0.0007903417546975425
+    -0.009083969707182315
+     -0.07336517453073049
+       0.3547204216223377
+ 5.03e+10    
+       0.3559326733356487
+     -0.07346232456503327
+       0.3662196744644612
+     -0.00910005358716352
+     -0.03545663370420072
+       0.3663821485101702
+   -0.0007478958812128769
+    -0.009095853642949972
+     -0.07353384130604762
+       0.3552323193691958
+ 5.04e+10    
+       0.3564441187614836
+     -0.07363095743985254
+       0.3667975505613469
+    -0.009111533580302447
+     -0.03556145528578753
+       0.3669603409371993
+   -0.0007051738474673794
+    -0.009107491493995106
+     -0.07370258029092851
+       0.3557432151345665
+ 5.05e+10    
+       0.3569545555736847
+     -0.07379965939651792
+       0.3673746823861617
+     -0.00912276478649897
+     -0.03566647871782854
+       0.3675377886633296
+   -0.0006621780501335007
+    -0.009118881993277785
+     -0.07387138909867616
+       0.3562531076721649
+ 5.06e+10    
+       0.3574639825884357
+     -0.07396842803666252
+       0.3679510689176002
+     -0.00913374594160705
+     -0.03577170398116805
+       0.3681144906504997
+   -0.0006189109130225318
+    -0.009130023875815988
+     -0.07404026532376931
+       0.3567619957349364
+ 5.07e+10    
+       0.3579723986212763
+     -0.07413726094324145
+       0.3685267091188574
+    -0.009144475783671573
+     -0.03587713105874052
+       0.3686904458464028
+   -0.0005753748864903401
+    -0.009140915878690658
+     -0.07420920654227289
+       0.3572698780751256
+ 5.08e+10    
+       0.3584798024871478
+     -0.07430615568094816
+       0.3691016019377134
+    -0.009154953052933099
+     -0.03598275993567353
+       0.3692656531845585
+    -0.000531572446835478
+    -0.009151556741051611
+      -0.0743782103122563
+       0.3577767534443568
+ 5.09e+10    
+        0.358986193000446
+     -0.07447510979663591
+       0.3696757463066327
+    -0.009165176491834176
+     -0.03608859059938958
+       0.3698401115843895
+   -0.0004875060956893581
+    -0.009161945204125468
+     -0.07454727417421522
+       0.3582826205937098
+ 5.1e+10     
+       0.3594915689750731
+     -0.07464412081974407
+       0.3702491411428631
+    -0.009175144845027067
+     -0.03619462303970705
+       0.3704138199513048
+   -0.0004431783593989919
+    -0.009172080011224465
+      -0.0747163956514996
+       0.3587874782738033
+ 5.11e+10    
+       0.3599959292244896
+     -0.07481318626272951
+       0.3708217853485444
+    -0.009184856859382973
+     -0.03630085724893976
+       0.3709867771767907
+   -0.0003985917884019739
+    -0.009181959907757383
+      -0.0748855722507458
+       0.3592913252348769
+ 5.12e+10    
+       0.3604992725617765
+     -0.07498230362150324
+       0.3713936778108243
+    -0.009194311284002507
+     -0.03640729322199645
+       0.3715589821385045
+   -0.0003537489565944138
+    -0.009191583641241218
+     -0.07505480146231419
+        0.359794160226875
+ 5.13e+10    
+        0.361001597799689
+     -0.07515147037587214
+       0.3719648174019767
+    -0.009203506870227859
+     -0.03651393095647818
+       0.3721304337003793
+    -0.000308652460691221
+    -0.009200949961314923
+     -0.07522408076073239
+       0.3602959819995385
+ 5.14e+10    
+       0.3615029037507213
+     -0.07532068398998537
+       0.3725352029795304
+    -0.009212442371656105
+     -0.03662077045277581
+       0.3727011307127278
+   -0.0002633049195796136
+    -0.009210057619754203
+     -0.07539340760514182
+       0.3607967893024905
+ 5.15e+10    
+       0.3620031892271711
+     -0.07548994191278602
+       0.3731048333864005
+    -0.009221116544154247
+     -0.03672781171416564
+       0.3732710720123605
+   -0.0002177089736653717
+    -0.009218905370487878
+     -0.07556277943975109
+       0.3612965808853323
+ 5.16e+10    
+       0.3625024530412029
+     -0.07565924157846707
+       0.3736737074510263
+    -0.009229528145875415
+      -0.0368350547469047
+       0.3738402564227038
+    -0.000171867284212341
+      -0.0092274919696156
+     -0.07573219369429289
+       0.3617953554977359
+ 5.17e+10    
+       0.3630006940049189
+     -0.07582858040693295
+        0.374241823987516
+    -0.009237675937276441
+     -0.03694249956032454
+       0.3744086827539226
+   -0.0001257825326751757
+    -0.009235816175427075
+     -0.07590164778448616
+       0.3622931118895432
+ 5.18e+10    
+       0.3634979109304278
+     -0.07599795580426495
+        0.374809181795797
+    -0.009245558681137103
+     -0.03705014616692433
+       0.3749763498030559
+   -7.945742002542677e-05
+    -0.009243876748422655
+       -0.076071139112503
+       0.3627898488108614
+ 5.19e+10    
+       0.3639941026299209
+     -0.07616736516319247
+       0.3753757796617698
+    -0.009253175142580474
+     -0.03715799458246285
+         0.37554325635415
+   -3.289466607127463e-05
+    -0.009251672451335111
+      -0.0762406650674409
+       0.3632855650121708
+ 5.2e+10     
+       0.3644892679157446
+     -0.07633680586356821
+       0.3759416163574695
+    -0.009260524089094651
+     -0.03726604482604942
+       0.3761094011784007
+    1.390299122921773e-05
+    -0.009259202049153141
+     -0.07641022302579797
+       0.3637802592444226
+ 5.21e+10    
+         0.36498340560048
+     -0.07650627527284747
+       0.3765066906412295
+     -0.00926760429055617
+     -0.03737429692023344
+        0.376674783034302
+    6.093279646088756e-05
+    -0.009266464309146001
+     -0.07657981035195499
+       0.3642739302591496
+ 5.22e+10    
+       0.3654765144970219
+     -0.07667577074657377
+       0.3770710012578566
+    -0.009274414519254188
+     -0.03748275089109389
+       0.3772394006677964
+    0.0001081919774504011
+    -0.009273458000889578
+     -0.07674942439866046
+       0.3647665768085733
+ 5.23e+10    
+       0.3659685934186613
+     -0.07684528962886675
+       0.3776345469388028
+    -0.009280953549916536
+     -0.03759140676832664
+       0.3778032528124343
+    0.0001556777459709962
+    -0.009280181896293576
+     -0.07691906250752098
+       0.3652581976457146
+ 5.24e+10    
+       0.3664596411791724
+     -0.07701482925291672
+       0.3781973264023485
+    -0.009287220159736931
+     -0.03770026458533119
+        0.378366338189535
+    0.0002033872984530726
+    -0.009286634769630531
+     -0.07708872200949547
+       0.3657487915245082
+ 5.25e+10    
+       0.3669496565928971
+     -0.07718438694148247
+       0.3787593383537882
+     -0.00929321312840317
+     -0.03780932437929664
+       0.3789286555083551
+     0.000251317816700281
+    -0.009292815397565544
+      -0.0772584002253951
+       0.3662383571999188
+ 5.26e+10    
+       0.3674386384748348
+     -0.07735396000739261
+       0.3793205814856206
+    -0.009298931238127186
+     -0.03791858619128623
+       0.3794902034662621
+    0.0002994664686110709
+    -0.009298722559187653
+     -0.07742809446638596
+       0.3667268934280565
+ 5.27e+10    
+       0.3679265856407367
+     -0.07752354575405412
+       0.3798810544777456
+    -0.009304373273675807
+     -0.03802805006632057
+       0.3800509807489083
+    0.0003478304089056361
+     -0.00930435503604252
+     -0.07759780203449718
+       0.3672143989663003
+ 5.28e+10    
+       0.3684134969071977
+     -0.07769314147596218
+       0.3804407559976611
+    -0.009309538022403282
+     -0.03813771605346056
+       0.3806109860304163
+    0.0003964067798578731
+    -0.009309711612166108
+     -0.07776752022313384
+         0.36770087257342
+ 5.29e+10    
+       0.3688993710917536
+     -0.07786274445921552
+       0.3809996847006727
+    -0.009314424274284505
+     -0.03824758420588883
+       0.3811702179735639
+    0.0004451927120323062
+    -0.009314791074119822
+     -0.07793724631759219
+       0.3681863130097002
+ 5.3e+10     
+       0.3693842070129809
+     -0.07803235198203674
+       0.3815578392300976
+    -0.009319030821950125
+     -0.03835765458098948
+       0.3817286752299762
+    0.0004941853250260263
+     -0.00931959221102684
+     -0.07810697759558208
+       0.3686707190370704
+ 5.31e+10    
+       0.3698680034905967
+     -0.07820196131529455
+       0.3821152182174794
+    -0.009323356460722149
+     -0.03846792724042798
+       0.3822863564403186
+    0.0005433817282149795
+    -0.009324113814609536
+     -0.07827671132774983
+       0.3691540894192316
+ 5.32e+10    
+       0.3703507593455653
+     -0.07837156972303365
+       0.3826718202828092
+    -0.009327399988651302
+     -0.03857840225022934
+       0.3828432602345008
+    0.0005927790215050647
+    -0.009328354679228273
+     -0.07844644477820936
+       0.3696364229217916
+ 5.33e+10    
+       0.3708324734002002
+     -0.07854117446300438
+       0.3832276440347425
+    -0.009331160206555231
+     -0.03868907968085494
+       0.3833993852318789
+    0.0006423742960873695
+    -0.009332313601921216
+     -0.07861617520507388
+       0.3701177183123976
+ 5.34e+10    
+       0.3713131444782772
+     -0.07871077278720033
+        0.383782688070827
+    -0.009334635918058004
+      -0.0387999596072786
+       0.3839547300414632
+    0.0006921646351975644
+    -0.009335989382445248
+     -0.07878589986099367
+       0.3705979743608747
+ 5.35e+10    
+       0.3717927714051416
+      -0.0788803619423968
+       0.3843369509777337
+    -0.009337825929630696
+     -0.03891104210906181
+       0.3845092932621332
+    0.0007421471148794439
+    -0.009339380823318347
+     -0.07895561599369742
+       0.3710771898393643
+ 5.36e+10    
+       0.3722713530078239
+     -0.07904993917069621
+       0.3848904313314902
+    -0.009340729050632955
+     -0.03902232727042769
+       0.3850630734828534
+     0.000792318804752105
+    -0.009342486729862584
+     -0.07912532084653717
+       0.3715553635224658
+ 5.37e+10    
+       0.3727488881151543
+     -0.07921950171007393
+       0.3854431276977173
+    -0.009343344093356016
+     -0.03913381518033357
+       0.3856160692828939
+    0.0008426767687809338
+     -0.00934530591024856
+     -0.07929501165903743
+       0.3720324941873812
+ 5.38e+10    
+       0.3732253755578818
+     -0.07938904679493099
+       0.3859950386318706
+    -0.009345669873066377
+     -0.03924550593254289
+        0.386168279232056
+    0.0008932180660520292
+    -0.009347837175540793
+     -0.07946468566744823
+       0.3725085806140616
+ 5.39e+10    
+       0.3737008141687932
+     -0.07955857165664881
+       0.3865461626794873
+    -0.009347705208050646
+       -0.039357399625696
+       0.3867197018909007
+    0.0009439397515498568
+     -0.00935007933974407
+     -0.07963434010530202
+       0.3729836215853564
+ 5.4e+10     
+       0.3741752027828377
+     -0.07972807352414861
+       0.3870964983764344
+     -0.00934944891966155
+     -0.03946949636337978
+       0.3872703358109802
+    0.0009948388769381259
+    -0.009352031219851085
+     -0.07980397220397348
+       0.3734576158871631
+ 5.41e+10    
+       0.3746485402372512
+      -0.0798975496244536
+       0.3876460442491606
+    -0.009350899832364775
+     -0.03958179625419628
+       0.3878201795350771
+     0.001045912491343594
+    -0.009353691635890567
+     -0.07997357919324491
+       0.3739305623085825
+ 5.42e+10    
+       0.3751208253716846
+     -0.08006699718325544
+       0.3881947988149514
+    -0.009352056773786923
+     -0.03969429941183035
+       0.3883692315974415
+     0.001097157642142697
+    -0.009355059410976935
+     -0.08014315830187335
+       0.3744024596420734
+ 5.43e+10    
+       0.3755920570283326
+     -0.08023641342548446
+       0.3887427605821918
+    -0.009352918574764061
+     -0.03980700595511603
+       0.3889174905240348
+     0.001148571375750583
+    -0.009356133371360504
+     -0.08031270675816177
+       0.3748733066836116
+ 5.44e+10    
+       0.3760622340520688
+     -0.08040579557588273
+       0.3892899280506247
+    -0.009353484069391868
+     -0.03991991600810212
+        0.389464954832781
+     0.001200150738412879
+     -0.00935691234647882
+     -0.08048222179053595
+       0.3753431022328512
+ 5.45e+10    
+       0.3765313552905774
+     -0.08057514085958097
+        0.389836299711621
+    -0.009353752095075853
+     -0.04003302970011691
+       0.3900116230338108
+      0.00125189277699939
+      -0.0093573951690087
+     -0.08065170062812088
+       0.3758118450932856
+ 5.46e+10    
+       0.3769994195944927
+     -0.08074444650267916
+       0.3903818740484459
+    -0.009353721492583138
+      -0.0401463471658309
+       0.3905574936297208
+     0.001303794539799991
+    -0.009357580674919402
+     -0.08082114050132438
+        0.376279534072415
+ 5.47e+10    
+       0.3774664258175381
+      -0.0809137097328301
+       0.3909266495365322
+    -0.009353391106094625
+     -0.04025986854532015
+       0.3911025651158295
+     0.001355853077322358
+    -0.009357467703526197
+     -0.08099053864242259
+       0.3767461679819135
+ 5.48e+10    
+       0.3779323728166685
+     -0.08108292777982658
+       0.3914706246437558
+    -0.009352759783258282
+     -0.04037359398412681
+       0.3916468359804365
+     0.001408065443091373
+    -0.009357055097545303
+     -0.08115989228614789
+       0.3772117456377983
+ 5.49e+10    
+       0.3783972594522135
+       -0.081252097876192
+       0.3920137978307153
+    -0.009351826375242869
+     -0.04048752363332035
+       0.3921903047050898
+      0.00146042869445007
+    -0.009356341703149152
+     -0.08132919867028274
+        0.377676265860604
+ 5.5e+10     
+       0.3788610845880261
+     -0.08142121725777331
+       0.3925561675510112
+    -0.009350589736792963
+     -0.04060165764955612
+       0.3927329697648492
+     0.001512939893361675
+    -0.009355326370022543
+     -0.08149845503625394
+       0.3781397274755551
+ 5.51e+10    
+       0.3793238470916308
+     -0.08159028316433893
+       0.3930977322515329
+    -0.009349048726284072
+     -0.04071599619513449
+        0.393274829628559
+     0.001565596107213131
+    -0.009354007951419755
+     -0.08166765862973177
+       0.3786021293127447
+ 5.52e+10    
+       0.3797855458343751
+     -0.08175929284017777
+       0.3936384903727448
+    -0.009347202205778869
+      -0.0408305394380581
+       0.3938158827591209
+     0.001618394409619101
+    -0.009352385304221757
+      -0.0818368067012326
+       0.3790634702073134
+ 5.53e+10    
+       0.3802461796915838
+     -0.08192824353470265
+       0.3941784403489753
+    -0.009345049041084064
+     -0.04094528755208793
+       0.3943561276137699
+     0.001671331881227017
+    -0.009350457288994861
+     -0.08200589650672349
+       0.3795237489996322
+ 5.54e+10    
+        0.380705747542716
+     -0.08209713250305652
+       0.3947175806087109
+     -0.00934258810180769
+     -0.04106024071679945
+       0.3948955626443535
+     0.001724405610522572
+    -0.009348222770049304
+      -0.0821749253082302
+        0.379982964535485
+ 5.55e+10    
+       0.3811642482715227
+     -0.08226595700672167
+       0.3952559095748919
+    -0.009339818261417297
+     -0.04117539911763672
+       0.3954341862976155
+     0.001777612694635545
+     -0.00934568061549893
+     -0.08234389037444928
+       0.3804411156662559
+ 5.56e+10    
+       0.3816216807662073
+     -0.08243471431413132
+       0.3957934256652104
+    -0.009336738397298426
+     -0.04129076294596627
+        0.395971997015478
+       0.0018309502401457
+    -0.009342829697321076
+     -0.08251278898136151
+       0.3808982012491174
+ 5.57e+10    
+       0.3820780439195922
+     -0.08260340170128526
+       0.3963301272924093
+    -0.009333347390813871
+     -0.04140633239912968
+       0.3965089932353314
+      0.00188441536388879
+     -0.00933966889141731
+     -0.08268161841284945
+       0.3813542201472236
+ 5.58e+10    
+       0.3825333366292809
+     -0.08277201645236712
+       0.3968660128645873
+    -0.009329644127363286
+     -0.04152210768049547
+       0.3970451733903248
+     0.001938005193762193
+    -0.009336197077674385
+     -0.08285037596131745
+       0.3818091712298998
+ 5.59e+10    
+       0.3829875577978288
+     -0.08294055586036546
+        0.397401080785505
+    -0.009325627496443396
+     -0.04163808899950992
+       0.3975805359096569
+     0.001991716869530209
+    -0.009332413140025898
+     -0.08301905892831435
+       0.3822630533728414
+ 5.6e+10     
+       0.3834407063329117
+     -0.08310901722769616
+       0.3979353294548903
+    -0.009321296391708655
+      -0.0417542765717471
+       0.3981150792188775
+     0.002045547543628587
+    -0.009328315966514199
+     -0.08318766462516031
+       0.3827158654583115
+ 5.61e+10    
+       0.3838927811475004
+     -0.08327739786682993
+       0.3984687572687508
+    -0.009316649711032082
+     -0.04187067061895792
+       0.3986488017401765
+     0.002099494381968387
+    -0.009323904449352874
+     -0.08335619037357306
+        0.383167606375339
+ 5.62e+10    
+        0.384343781160034
+     -0.08344569510091972
+       0.3990013626196874
+     -0.00931168635656681
+     -0.04198727136911852
+       0.3991817018926943
+     0.002153554564738653
+    -0.009319177484989524
+     -0.08352463350630134
+       0.3836182750199235
+ 5.63e+10    
+       0.3847937052946001
+     -0.08361390626443291
+       0.3995331438972075
+    -0.009306405234807824
+     -0.04210407905647749
+       0.3997137780928188
+     0.002207725287207999
+    -0.009314133974168791
+     -0.08369299136775707
+       0.3840678702952393
+ 5.64e+10    
+       0.3852425524811113
+     -0.08378202870378408
+       0.4000640994880411
+    -0.009300805256654021
+     -0.04222109392160266
+       0.4002450287544938
+     0.002262003760524611
+    -0.009308772821995799
+     -0.08386126131465232
+       0.3845163911118412
+ 5.65e+10    
+       0.3856903216554897
+     -0.08395005977797272
+       0.4005942277764636
+    -0.009294885337470469
+     -0.04233831621142634
+       0.4007754522895266
+      0.00231638721251485
+    -0.009303092937999932
+     -0.08402944071663818
+       0.3849638363878769
+ 5.66e+10    
+       0.3861370117598499
+     -0.08411799685922024
+       0.4011235271446142
+    -0.009288644397151068
+     -0.04245574617929092
+       0.4013050471078977
+     0.002370872888479775
+    -0.009297093236198602
+      -0.0841975269569458
+        0.385410205049295
+ 5.67e+10    
+       0.3865826217426871
+     -0.08428583733361331
+       0.4016519959728218
+    -0.009282081360181316
+      -0.0425733840849926
+       0.4018338116180754
+     0.002425458051989818
+    -0.009290772635161386
+     -0.08436551743303071
+       0.3858554960300615
+ 5.68e+10    
+       0.3870271505590645
+     -0.08445357860174478
+       0.4021796326399272
+    -0.009275195155701303
+     -0.04269123019482441
+       0.4023617442273268
+     0.002480139985677165
+     -0.00928413005807447
+     -0.08453340955721793
+       0.3862997082723736
+ 5.69e+10    
+       0.3874705971708059
+     -0.08462121807936168
+       0.4027064355236145
+    -0.009267984717568714
+     -0.04280928478161952
+       0.4028888433420397
+     0.002534915992025775
+    -0.009277164432804722
+     -0.08470120075735144
+         0.38674284072688
+ 5.7e+10     
+       0.3879129605466882
+     -0.08478875319801162
+       0.4032324030007368
+    -0.009260448984422104
+     -0.04292754812479225
+       0.4034151073680379
+     0.002589783394158665
+    -0.009269874691964417
+      -0.0848688884774443
+       0.3871848923528995
+ 5.71e+10    
+       0.3883542396626373
+     -0.08495618140569358
+       0.4037575334476504
+    -0.009252586899744243
+      -0.0430460205103799
+       0.4039405347109046
+     0.002644739536622588
+     -0.00926225977297573
+     -0.08503647017833213
+       0.3876258621186457
+ 5.72e+10    
+       0.3887944335019265
+      -0.0851235001675104
+        0.404281825240546
+    -0.009244397411925107
+     -0.04316470223108221
+       0.4044651237763043
+     0.002699781786169352
+    -0.009254318618135153
+     -0.08520394333832708
+       0.3880657490014481
+ 5.73e+10    
+       0.3892335410553765
+     -0.08529070696632257
+       0.4048052767557851
+    -0.009235879474325477
+     -0.04328359358630193
+       0.4049888729703091
+     0.002754907532534319
+    -0.009246050174678182
+     -0.08537130545387639
+        0.388504551987984
+ 5.74e+10    
+       0.3896715613215577
+     -0.08545779930340475
+       0.4053278863702346
+    -0.009227032045339976
+     -0.04340269488218302
+       0.4055117806997254
+     0.002810114189211158
+     -0.00923745339484364
+      -0.0855385540402207
+       0.3889422700745033
+ 5.75e+10    
+       0.3901084933069948
+     -0.08562477469910412
+       0.4058496524616065
+    -0.009217854088460271
+     -0.04352200643164913
+       0.4060338453724223
+     0.002865399194223199
+    -0.009228527235938085
+     -0.08570568663205537
+       0.3893789022670614
+ 5.76e+10    
+       0.3905443360263739
+     -0.08579163069350075
+       0.4063705734087981
+     -0.00920834457233805
+     -0.04364152855444138
+       0.4065550653976643
+      0.00292076001089087
+    -0.009219270660400087
+     -0.08587270078419451
+       0.3898144475817539
+ 5.77e+10    
+       0.3909790885027509
+     -0.08595836484706951
+       0.4068906475922333
+    -0.009198502470847853
+     -0.04376126157715518
+       0.4070754391864417
+     0.002976194128595098
+    -0.009209682635864101
+     -0.08603959407223435
+       0.3902489050449484
+ 5.78e+10    
+       0.3914127497677631
+      -0.0861249747413436
+       0.4074098733942041
+    -0.009188326763149842
+     -0.04388120583327645
+       0.4075949651518081
+     0.003031699063536629
+    -0.009199762135224505
+     -0.08620636409322208
+       0.3906822736935261
+ 5.79e+10    
+       0.3918453188618415
+     -0.08629145797958075
+       0.4079282491992192
+    -0.009177816433752052
+     -0.04400136166321757
+       0.4081136417092131
+      0.00308727235949088
+    -0.009189508136699106
+     -0.08637300846632318
+       0.3911145525751184
+ 5.8e+10     
+       0.3922767948344283
+     -0.08645781218743023
+       0.4084457733943456
+    -0.009166970472572587
+     -0.04412172941435229
+       0.4086314672768431
+     0.003142911588558049
+    -0.009178919623892289
+     -0.08653952483349246
+       0.3915457407483503
+ 5.81e+10    
+        0.392707176744193
+     -0.08662403501360164
+       0.4089624443695588
+     -0.00915578787500154
+     -0.04424230944105013
+       0.4091484402759587
+     0.003198614351908714
+    -0.009167995585858216
+     -0.08670591086014591
+       0.3919758372830832
+ 5.82e+10    
+       0.3931364636592505
+     -0.08679012413053563
+       0.4094782605180929
+    -0.009144267641962231
+     -0.04436310210471109
+       0.4096645591312375
+     0.003254378280524161
+    -0.009156735017163263
+     -0.08687216423583412
+       0.3924048412606605
+ 5.83e+10    
+        0.393564654657387
+     -0.08695607723507626
+       0.4099932202367878
+    -0.009132408779972481
+     -0.04448410777379832
+       0.4101798222711159
+     0.003310201035931766
+    -0.009145136917948195
+     -0.08703828267491821
+       0.3928327517741564
+ 5.84e+10    
+       0.3939917488262786
+     -0.08712189204914367
+        0.410507321926444
+    -0.009120210301205141
+     -0.04460532682387128
+       0.4106942281281335
+      0.00336608031093482
+    -0.009133200293990007
+     -0.08720426391724638
+       0.3932595679286254
+ 5.85e+10    
+       0.3944177452637211
+      -0.0872875663204097
+       0.4110205639921744
+    -0.009107671223548171
+     -0.04472675963761848
+       0.4112077751392788
+     0.003422013830336786
+    -0.009120924156763015
+     -0.08737010572883158
+       0.3936852888413521
+ 5.86e+10    
+        0.394842643077856
+     -0.08745309782297385
+       0.4115329448437572
+    -0.009094790570664568
+     -0.04484840660488882
+        0.411720461746336
+     0.003477999351660072
+    -0.009108307523499736
+     -0.08753580590253149
+       0.3941099136421075
+ 5.87e+10    
+       0.3952664413874011
+     -0.08761848435804129
+       0.4120444628959944
+    -0.009081567372051159
+     -0.04497026812272382
+        0.412232286396235
+     0.003534034665858409
+    -0.009095349417250894
+      -0.0877013622587301
+       0.3945334414734027
+ 5.88e+10    
+       0.3956891393218808
+     -0.08778372375460115
+       0.4125551165690674
+    -0.009068000663097184
+     -0.04509234459538807
+       0.4127432475413984
+     0.003590117598023477
+    -0.009082048866945172
+     -0.08786677264601879
+       0.3949558714907486
+ 5.89e+10    
+       0.3961107360218626
+     -0.08794881387010701
+       0.4130649042888925
+    -0.009054089485142292
+     -0.04521463643439994
+       0.4132533436400952
+     0.003646246008084967
+    -0.009068404907447841
+     -0.08803203494188055
+       0.3953772028629126
+ 5.9e+10     
+       0.3965312306391906
+     -0.08811375259115804
+       0.4135738244874845
+    -0.009039832885533595
+      -0.0453371440585621
+       0.4137625731567923
+     0.003702417791504232
+    -0.009054416579619215
+     -0.08819714705337428
+       0.3957974347721814
+ 5.91e+10    
+        0.396950622337223
+     -0.08827853783418084
+       0.4140818756033123
+    -0.009025229917682237
+      -0.0454598678939908
+       0.4142709345625079
+      0.00375863087996126
+    -0.009040082930372111
+     -0.08836210691782052
+       0.3962165664146234
+ 5.92e+10    
+       0.3973689102910747
+     -0.08844316754611359
+        0.414589056081662
+    -0.009010279641119117
+      -0.0455828083741457
+       0.4147784263351679
+     0.003814883242034658
+    -0.009025403012728403
+     -0.08852691250348882
+       0.3966345970003564
+ 5.93e+10    
+       0.3977860936878548
+     -0.08860763970508896
+       0.4150953643749996
+    -0.008994981121549875
+     -0.04570596593985871
+       0.4152850469599589
+     0.003871172883874595
+    -0.009010375885875258
+     -0.08869156181028437
+       0.3970515257538099
+ 5.94e+10    
+       0.3982021717269127
+     -0.08877195232112113
+       0.4156007989433333
+    -0.008979333430908915
+     -0.04582934103936313
+       0.4157907949296904
+     0.003927497849868697
+    -0.008995000615219873
+     -0.08885605287043824
+       0.3974673519139971
+ 5.95e+10    
+       0.3986171436200823
+     -0.08893610343678988
+       0.4161053582545778
+    -0.008963335647412782
+     -0.04595293412832151
+       0.4162956687451466
+     0.003983856223300099
+    -0.008979276272443985
+     -0.08902038374919552
+       0.3978820747347843
+ 5.96e+10    
+       0.3990310085919294
+     -0.08910009112792901
+       0.4166090407849182
+    -0.008946986855612449
+     -0.04607674566985416
+       0.4167996669154514
+     0.004040246126998338
+    -0.008963201935556969
+     -0.08918455254550683
+       0.3982956934851627
+ 5.97e+10    
+       0.3994437658800002
+     -0.08926391350431302
+       0.4171118450191765
+    -0.008930286146444774
+     -0.04620077613456679
+        0.417302787958426
+     0.004096665723982188
+    -0.008946776688948303
+     -0.08934855739271895
+       0.3987082074495234
+ 5.98e+10    
+       0.3998554147350714
+     -0.08942756871034536
+        0.417613769451179
+    -0.008913232617282784
+     -0.04632502600057852
+       0.4178050304009506
+     0.004153113218094501
+    -0.008929999623438567
+      -0.0895123964592672
+       0.3991196159279297
+ 5.99e+10    
+       0.4002659544214049
+     -0.08959105492574838
+       0.4181148125841224
+    -0.008895825371985274
+     -0.04644949575354867
+       0.4183063927793267
+     0.004209586854629259
+    -0.008912869836330276
+     -0.08967606794936749
+       0.3995299182363994
+ 6e+10       
+       0.4006753842169982
+     -0.08975437036625129
+       0.4186149729309432
+    -0.008878063520944855
+     -0.04657418588670448
+       0.4188068736396406
+     0.004266084920949847
+    -0.008895386431456574
+     -0.08983957010370999
+       0.3999391137071788
+ 6.01e+10    
+       0.4010837034138433
+     -0.08991751328428108
+       0.4191142490146842
+    -0.008859946181135527
+     -0.04669909690086764
+       0.4193064715381279
+     0.004322605747099197
+    -0.008877548519229495
+     -0.09000290120015261
+        0.400347201689026
+ 6.02e+10    
+       0.4014909113181828
+      -0.0900804819696526
+       0.4196126393688667
+    -0.008841472476158466
+     -0.04682422930448114
+       0.4198051850415359
+     0.004379147706401146
+     -0.00885935521668698
+      -0.0901660595544152
+       0.4007541815474925
+ 6.03e+10    
+       0.4018970072507698
+     -0.09024327475026023
+       0.4201101425378608
+    -0.008822641536287062
+     -0.04694958361363642
+       0.4203030127274936
+     0.004435709216053089
+    -0.008840805647538506
+     -0.09032904352077466
+       0.4011600526652065
+ 6.04e+10    
+       0.4023019905471268
+      -0.0904058899927675
+       0.4206067570772531
+    -0.008803452498510533
+       -0.047075160352099
+       0.4207999531848732
+     0.004492288737709492
+     -0.00882189894220959
+     -0.09049185149275896
+       0.4015648144421581
+ 6.05e+10    
+       0.4027058605578105
+     -0.09056832610329989
+       0.4211024815542205
+    -0.008783904506576413
+     -0.04720096005133526
+        0.421296005014161
+     0.004548884778056383
+     -0.00880263423788513
+     -0.09065448190384302
+       0.4019684662959854
+ 6.06e+10    
+       0.4031086166486744
+     -0.09073058152813585
+       0.4215973145479033
+    -0.008763996711031742
+     -0.04732698325053934
+       0.4217911668278252
+     0.004605495889376645
+    -0.008783010678550982
+     -0.09081693322814516
+       0.4023710076622643
+ 6.07e+10    
+       0.4035102582011337
+     -0.09089265475439948
+       0.4220912546497756
+    -0.008743728269262632
+     -0.04745323049665819
+       0.4222854372506807
+     0.004662120670105627
+    -0.008763027415035074
+     -0.09097920398112085
+       0.4027724379947974
+ 6.08e+10    
+       0.4039107846124336
+     -0.09105454431075091
+       0.4225843004640171
+    -0.008723098345532924
+     -0.04757970234441844
+       0.4227788149202628
+     0.004718757765377267
+    -0.008742683605046011
+     -0.09114129272026017
+       0.4031727567659031
+ 6.09e+10    
+       0.4043101952959169
+     -0.09121624876807995
+       0.4230764506078913
+    -0.008702106111021089
+     -0.04770639935635248
+       0.4232712984871935
+     0.004775405867560565
+    -0.008721978413211241
+     -0.09130319804578307
+       0.4035719634667117
+ 6.1e+10     
+       0.4047084896812942
+     -0.09137776674019733
+       0.4235677037121149
+    -0.008680750743855846
+      -0.0478333221028243
+       0.4237628866155548
+     0.004832063716785947
+    -0.008700911011113156
+     -0.09146491860133613
+       0.4039700576074568
+ 6.11e+10    
+       0.4051056672149146
+     -0.09153909688452665
+       0.4240580584212334
+    -0.008659031429150223
+     -0.04796047116205573
+       0.4242535779832569
+     0.004888730101461729
+     -0.00867948057732397
+     -0.09162645307468696
+       0.4043670387177704
+ 6.12e+10    
+       0.4055017273600395
+     -0.09170023790279623
+       0.4245475133939972
+    -0.008636947359034159
+      -0.0480878471201526
+       0.4247433712824104
+     0.004945403858780216
+    -0.008657686297438891
+     -0.09178780019842156
+       0.4047629063469813
+ 6.13e+10    
+       0.4058966695971161
+     -0.09186118854173134
+       0.4250360673037358
+    -0.008614497732685385
+     -0.04821545057113113
+       0.4252322652196995
+     0.005002083875213657
+    -0.008635527364107937
+     -0.09194895875063935
+        0.405157660064411
+ 6.14e+10    
+       0.4062904934240524
+     -0.09202194759374445
+       0.4255237188387307
+    -0.008591681756359097
+     -0.04834328211694342
+       0.4257202585167515
+     0.005058769086999523
+    -0.008613002977065942
+     -0.09210992755564831
+       0.4055512994596733
+ 6.15e+10    
+       0.4066831983564942
+     -0.09218251389762719
+       0.4260104667025945
+     -0.00856849864341554
+     -0.04847134236750447
+       0.4262073499105116
+     0.005115458480615276
+    -0.008590112343160962
+     -0.09227070548466014
+       0.4059438241429737
+ 6.16e+10    
+       0.4070747839281031
+     -0.09234288633924062
+       0.4264963096146445
+    -0.008544947614346217
+     -0.04859963194071849
+        0.426693538153615
+     0.005172151093242353
+    -0.008566854676381162
+     -0.09243129145648615
+       0.4063352337454137
+ 6.17e+10    
+       0.4074652496908374
+     -0.09250306385220655
+        0.426981246310281
+     -0.00852102789679832
+     -0.04872815146250514
+       0.4271788220147602
+     0.005228846013219168
+    -0.008543229197879781
+     -0.09259168443823049
+       0.4067255279192902
+ 6.18e+10    
+       0.4078545952152282
+      -0.0926630454185955
+       0.4274652755413597
+    -0.008496738725597461
+     -0.04885690156682654
+       0.4276632002790828
+      0.00528554238048326
+     -0.00851923513599848
+     -0.09275188344598426
+       0.4071147063384004
+ 6.19e+10    
+       0.4082428200906654
+     -0.09282283006961803
+       0.4279483960765712
+     -0.00847207934276855
+     -0.04898588289571383
+       0.4281466717485272
+     0.005342239387002075
+    -0.008494871726288851
+     -0.09291188754551892
+       0.4075027686983463
+ 6.2e+10     
+       0.4086299239256786
+     -0.09298241688631195
+       0.4284306067018161
+    -0.008447048997555051
+     -0.04911509609929433
+       0.4286292352422252
+     0.005398936277192713
+    -0.008470138211532035
+     -0.09307169585298029
+       0.4078897147168413
+ 6.21e+10    
+        0.409015906348219
+     -0.09314180500023106
+       0.4289119062205828
+    -0.008421646946436092
+     -0.04924454183581906
+       0.4291108895968657
+     0.005455632348330029
+    -0.008445033841756839
+     -0.09323130753557893
+       0.4082755441340158
+ 6.22e+10    
+       0.4094007670059496
+     -0.09330099359413264
+       0.4293922934543214
+    -0.008395872453142111
+     -0.04937422077168967
+        0.429591633667071
+     0.005512326950943439
+    -0.008419557874255405
+      -0.0933907218122831
+       0.4086602567127261
+ 6.23e+10    
+       0.4097845055665238
+     -0.09345998190266337
+       0.4298717672428231
+    -0.008369724788668315
+     -0.04950413358148631
+       0.4300714663257709
+     0.005569019489201863
+    -0.008393709573597525
+     -0.09354993795450878
+       0.4090438522388622
+ 6.24e+10    
+       0.4101671217178793
+     -0.09361876921304582
+       0.4303503264445956
+    -0.008343203231286275
+     -0.04963428094799573
+        0.430550386464578
+     0.005625709421287127
+    -0.008367488211642616
+     -0.09370895528680984
+       0.4094263305216582
+ 6.25e+10    
+       0.4105486151685211
+     -0.09377735486576273
+       0.4308279699372383
+    -0.008316307066553555
+     -0.04976466356223944
+       0.4310283929941617
+     0.005682396259755487
+    -0.008340893067549943
+     -0.09386777318756737
+       0.4098076913940024
+ 6.26e+10    
+       0.4109289856478129
+     -0.09393573825524136
+       0.4313046966178227
+    -0.008289035587321466
+     -0.04989528212350231
+        0.431505484844622
+     0.005739079571886987
+    -0.008313923427786736
+     -0.09402639108967716
+       0.4101879347127487
+ 6.27e+10    
+       0.4113082329062641
+     -0.09409391883053557
+       0.4317805054032625
+    -0.008261388093740607
+     -0.05002613733936071
+       0.4319816609658644
+     0.005795758980022977
+    -0.008286578586134227
+     -0.09418480848123714
+       0.4105670603590285
+ 6.28e+10    
+       0.4116863567158235
+     -0.09425189609600872
+       0.4322553952306963
+    -0.008233363893264489
+     -0.05015722992571316
+       0.4324569203279776
+      0.00585243416189137
+    -0.008258857843691677
+     -0.09434302490623435
+       0.4109450682385639
+ 6.29e+10    
+        0.412063356870169
+     -0.09440966961201355
+       0.4327293650578584
+     -0.00820496230065107
+     -0.05028856060680802
+       0.4329312619216037
+     0.005909104850919658
+    -0.008230760508878537
+     -0.09450103996522852
+       0.4113219582819822
+ 6.3e+10     
+       0.4124392331849989
+     -0.09456723899557272
+       0.4332024138634608
+    -0.008176182637961906
+     -0.05042013011527539
+       0.4334046847583145
+     0.005965770836535485
+    -0.008202285897433843
+     -0.09465885331603642
+       0.4116977304451275
+ 6.31e+10    
+        0.412813985498326
+     -0.09472460392105514
+       0.4336745406475602
+    -0.008147024234559845
+     -0.05055193919215515
+       0.4338771878709858
+     0.006022431964454952
+    -0.008173433332414166
+     -0.09481646467441501
+       0.4120723847093787
+ 6.32e+10    
+       0.4131876136707706
+     -0.09488176412085512
+       0.4341457444319407
+    -0.008117486427103617
+     -0.05068398858692982
+       0.4343487703141726
+     0.006079088136958139
+    -0.008144202144188973
+      -0.0949738738147419
+       0.4124459210819635
+ 6.33e+10    
+       0.4135601175858533
+      -0.0950387193860662
+       0.4346160242604866
+    -0.008087568559541033
+     -0.05081627905755406
+       0.4348194311644789
+     0.006135739313152238
+    -0.008114591670433878
+     -0.09513108057069519
+       0.4128183395962737
+ 6.34e+10    
+       0.4139314971502931
+     -0.09519546956715697
+       0.4350853791995554
+    -0.008057269983099432
+     -0.05094881137048728
+       0.4352891695209377
+     0.006192385509221902
+    -0.008084601256121607
+     -0.09528808483593329
+       0.4131896403121847
+ 6.35e+10    
+       0.4143017522942991
+     -0.09535201457464221
+       0.4355538083383546
+    -0.008026590056274308
+     -0.05108158630072476
+       0.4357579845053787
+     0.006249026798666658
+    -0.008054230253510816
+     -0.09544488656477033
+       0.4135598233163684
+ 6.36e+10    
+       0.4146708829718692
+     -0.09550835437975533
+       0.4360213107893147
+    -0.007995528144815163
+     -0.05121460463183104
+       0.4362258752628044
+     0.006305663312525712
+    -0.008023478022132441
+     -0.09560148577285296
+       0.4139288887226152
+ 6.37e+10    
+       0.4150388891610829
+     -0.09566448901511622
+       0.4364878856884628
+    -0.007964083621709589
+     -0.05134786715597234
+       0.4366928409617624
+     0.006362295239589666
+    -0.007992343928773907
+      -0.0957578825378331
+       0.4142968366721483
+ 6.38e+10    
+       0.4154057708644027
+     -0.09582041857540173
+       0.4369535321957952
+    -0.007932255867164562
+     -0.05148137467395033
+       0.4371588807947184
+     0.006418922826599407
+    -0.007960827347460874
+     -0.09591407700004172
+       0.4146636673339444
+ 6.39e+10    
+       0.4157715281089671
+     -0.09597614321800899
+       0.4374182494956519
+    -0.007900044268585765
+     -0.05161512799523596
+       0.4376239939784259
+     0.006475546378431596
+    -0.007928927659436662
+     -0.09607006936315778
+       0.4150293809050511
+ 6.4e+10     
+        0.416136160946891
+       -0.096131663163722
+       0.4378820367970868
+    -0.007867448220554235
+     -0.05174912793800403
+       0.4380881797542993
+     0.006532166258271538
+    -0.007896644253139372
+     -0.09622585989487815
+       0.4153939776109068
+ 6.41e+10    
+       0.4164996694555621
+     -0.09628697869737282
+       0.4383448933342408
+    -0.007834467124800832
+     -0.05188337532916884
+       0.4385514373887876
+     0.006588782887772388
+    -0.007863976524176386
+      -0.0963814489275845
+        0.415757457705658
+ 6.42e+10    
+       0.4168620537379404
+     -0.09644209016850365
+       0.4388068183667114
+    -0.007801100390178079
+     -0.05201787100441925
+       0.4390137661737407
+     0.006645396747201479
+    -0.007830923875296563
+     -0.09653683685900753
+       0.4161198214724807
+ 6.43e+10    
+       0.4172233139228544
+     -0.09659699799202373
+       0.4392678111799262
+    -0.007767347432629895
+     -0.05215261580825541
+       0.4394751654267814
+     0.006702008375573183
+    -0.007797485716360179
+     -0.09669202415289133
+       0.4164810692238993
+ 6.44e+10    
+       0.4175834501653014
+     -0.09675170264886741
+       0.4397278710855084
+    -0.007733207675158449
+     -0.05228761059402552
+       0.4399356344916762
+     0.006758618370768531
+    -0.007763661464305844
+      -0.0968470113396537
+       0.4168412013021051
+ 6.45e+10    
+       0.4179424626467457
+     -0.09690620468664796
+       0.4401869974216498
+     -0.00769868054778891
+     -0.05242285622396336
+       0.4403951727387025
+     0.006815227389641427
+    -0.007729450543115642
+     -0.09700179901704556
+       0.4172002180792779
+ 6.46e+10    
+       0.4183003515754196
+     -0.09706050472031141
+       0.4406451895534785
+     -0.00766376548753146
+     -0.05255835356922686
+       0.4408537795650186
+     0.006871836148111531
+     -0.00769485238377713
+     -0.09715638785080802
+       0.4175581199579038
+ 6.47e+10    
+       0.4186571171866177
+      -0.0972146034327851
+       0.4411024468734256
+     -0.00762846193834082
+     -0.05269410350993646
+       0.4413114543950291
+     0.006928445421243587
+    -0.007659866424243147
+     -0.09731077857532658
+       0.4179149073710966
+ 6.48e+10    
+       0.4190127597430004
+     -0.09736850157562688
+       0.4415587688015934
+     -0.00759276935107346
+     -0.05283010693521502
+       0.4417681966807565
+     0.006985056043313315
+     -0.00762449210938896
+     -0.09746497199428469
+       0.4182705807829158
+ 6.49e+10    
+       0.4193672795348907
+      -0.0975221999696706
+       0.4420141547861208
+    -0.007556687183441821
+     -0.05296636474322781
+       0.4422240059022018
+     0.007041668907859852
+    -0.007588728890966876
+     -0.09761896898131311
+       0.4186251406886871
+ 6.5e+10     
+       0.4197206768805734
+     -0.09767569950566973
+       0.4424686043035509
+    -0.007520214899966531
+      -0.0531028778412236
+       0.4426788815677147
+     0.007098284967724687
+    -0.007552576227558345
+     -0.09777277048063795
+       0.4189785876153213
+ 6.51e+10    
+       0.4200729521265934
+     -0.09782900114493749
+       0.4429221168591932
+    -0.007483351971925506
+     -0.05323964714557614
+       0.4431328232143569
+     0.007154905235076933
+    -0.007516033584523224
+     -0.09792637750772708
+        0.419330922121635
+ 6.52e+10    
+       0.4204241056480554
+     -0.09798210591998678
+       0.4433746919874894
+    -0.007446097877300764
+     -0.05337667358182685
+       0.4435858304082654
+     0.007211530781425094
+    -0.007479100433946635
+     -0.09807979114993162
+       0.4196821447986655
+ 6.53e+10    
+       0.4207741378489228
+     -0.09813501493516541
+       0.4438263292523761
+    -0.007408452100722596
+     -0.05351395808472754
+        0.444037902745018
+     0.007268162737615378
+     -0.00744177625458328
+     -0.09823301256712778
+       0.4200322562699943
+ 6.54e+10    
+       0.4211230491623139
+     -0.09828772936728918
+       0.4442770282476454
+    -0.007370414133410929
+     -0.05365150159828468
+       0.4444890398499932
+     0.007324802293816099
+    -0.007404060531798692
+     -0.09838604299235411
+       0.4203812571920634
+ 6.55e+10    
+          0.4214708400508
+     -0.09844025046627254
+       0.4447267885973078
+    -0.007331983473114395
+     -0.05378930507580355
+       0.4449392413787343
+     0.007381450699488943
+    -0.007365952757508454
+     -0.09853888373244729
+       0.4207291482544915
+ 6.56e+10    
+       0.4218175110067058
+     -0.09859257955575802
+       0.4451756099559523
+    -0.007293159624046267
+     -0.05392736947993434
+       0.4453885070173069
+      0.00743810926334619
+    -0.007327452430114085
+      -0.0986915361686734
+       0.4210759301803939
+ 6.57e+10    
+       0.4221630625524038
+     -0.09874471803374003
+       0.4456234920091051
+    -0.007253942096818196
+      -0.0540656957827179
+       0.4458368364826625
+     0.007494779353294674
+    -0.007288559054436762
+      -0.0988440017573599
+       0.4214216037266993
+ 6.58e+10    
+       0.4225074952406115
+     -0.09889666737318779
+       0.4460704344735862
+    -0.007214330408370962
+     -0.05420428496563286
+       0.4462842295229932
+     0.007551462396365893
+    -0.007249272141648083
+     -0.09899628203052033
+        0.421766169684464
+ 6.59e+10    
+       0.4228508096546887
+     -0.09904842912266515
+       0.4465164370978698
+    -0.007174324081902765
+     -0.05434313801964369
+       0.4467306859180925
+     0.007608159878632883
+    -0.007209591209198299
+     -0.09914837859648003
+       0.4221096288791908
+ 6.6e+10     
+       0.4231930064089328
+     -0.09920000490694676
+       0.4469614996624375
+    -0.007133922646794529
+     -0.05448225594524931
+       0.4471762054797107
+      0.00766487334511294
+    -0.007169515780741605
+     -0.09930029314049696
+       0.4224519821711447
+ 6.61e+10    
+       0.4235340861488726
+     -0.09935139642763192
+       0.4474056219801338
+    -0.007093125638532978
+     -0.05462163975253242
+       0.4476207880519096
+     0.007721604399657698
+    -0.007129045386058934
+     -0.09945202742537945
+       0.4227932304556626
+ 6.62e+10    
+       0.4238740495515682
+     -0.09950260546375611
+       0.4478488038965218
+    -0.007051932598630402
+     -0.05476129046121047
+       0.4480644335114196
+     0.007778354704828541
+    -0.007088179560977993
+     -0.09960358329210184
+       0.4231333746634734
+ 6.63e+10    
+       0.4242128973258961
+     -0.09965363387239655
+       0.4482910452902329
+    -0.007010343074542168
+     -0.05490120910068652
+       0.4485071417679898
+     0.007835125981759498
+    -0.007046917847290439
+     -0.09975496266041617
+       0.4234724157610075
+ 6.64e+10    
+        0.424550630212851
+     -0.09980448358927851
+       0.4487323460733199
+    -0.006968356619581394
+     -0.05504139671010118
+       0.4489489127647418
+     0.007891920010006076
+    -0.007005259792666505
+     -0.09990616752946151
+        0.423810354750712
+ 6.65e+10    
+       0.4248872489858339
+     -0.09995515662937507
+       0.4491727061916054
+    -0.006925972792830882
+     -0.05518185433838652
+       0.4493897464785232
+     0.007948738627380917
+    -0.006963204950566612
+      -0.1000571999783696
+       0.4241471926713581
+ 6.66e+10    
+       0.4252227544509445
+      -0.1001056550875058
+       0.4496121256250336
+     -0.00688319115905218
+     -0.05532258304431908
+       0.4498296429202522
+     0.008005583729775832
+    -0.006920752880150588
+      -0.1002080621668673
+       0.4244829305983578
+ 6.67e+10    
+       0.4255571474472736
+      -0.1002559811389313
+       0.4500506043880149
+    -0.006840011288592117
+     -0.05546358389657535
+        0.450268602135269
+     0.008062457270970654
+    -0.006877903146183955
+       -0.100358756335875
+       0.4248175696440688
+ 6.68e+10    
+       0.4258904288471898
+      -0.1004061370399433
+       0.4504881425297739
+    -0.006796432757286547
+     -0.05560485797378736
+       0.4507066242036851
+      0.00811936126242852
+    -0.006834655318941235
+      -0.1005092848081033
+       0.4251511109581049
+ 6.69e+10    
+       0.4262225995566331
+      -0.1005561251284542
+        0.450924740134693
+    -0.006752455146361247
+     -0.05574640636459965
+       0.4511437092407244
+     0.008176297773078139
+    -0.006791008974107024
+      -0.1006596499886452
+       0.4254835557276453
+ 6.7e+10     
+       0.4265536605153996
+      -0.1007059478245793
+       0.4513603973226566
+    -0.006708078042330314
+     -0.05588823016772616
+       0.4515798573970723
+      0.00823326892908253
+    -0.006746963692673937
+      -0.1008098543655644
+       0.4258149051777402
+ 6.71e+10    
+         0.42688361269743
+      -0.1008556076312193
+       0.4517951142493934
+    -0.006663301036891498
+     -0.05603033049200992
+       0.4520150688592157
+     0.008290276913594883
+    -0.006702519060837749
+       -0.100959900510481
+       0.4261451605716156
+ 6.72e+10    
+        0.427212457111095
+       -0.101005107134636
+       0.4522288911068166
+    -0.006618123726819003
+     -0.05617270845648224
+       0.4524493438497876
+     0.008347323966500817
+    -0.006657674669890017
+      -0.1011097910791528
+        0.426474323210979
+ 6.73e+10    
+       0.4275401947994811
+      -0.1011544490050269
+       0.4526617281233627
+    -0.006572545713853655
+     -0.05631536519042265
+       0.4528826826279049
+     0.008404412384148147
+    -0.006612430116108002
+      -0.1012595288120538
+       0.4268023944363231
+ 6.74e+10    
+       0.4278668268406742
+      -0.1013036359970941
+       0.4530936255643307
+    -0.006526566604589982
+     -0.05645830183342127
+       0.4533150854895087
+     0.008461544519063068
+    -0.006566785000641394
+      -0.1014091165349482
+       0.4271293756272273
+ 6.75e+10    
+       0.4281923543480405
+      -0.1014526709506101
+       0.4535245837322157
+    -0.006480186010360999
+     -0.05660151953544086
+       0.4537465527677019
+     0.008518722779653768
+    -0.006520738929396808
+      -0.1015585571594615
+       0.4274552682026582
+ 6.76e+10    
+       0.4285167784705107
+      -0.1016015567909813
+       0.4539546029670455
+    -0.006433403547119835
+     -0.05674501945688054
+       0.4541770848330858
+     0.008575949629901014
+    -0.006474291512919155
+      -0.1017078536836464
+       0.4277800736212687
+ 6.77e+10    
+       0.4288401003928576
+      -0.1017502965298051
+       0.4543836836467136
+    -0.006386218835318912
+     -0.05688880276864013
+       0.4546066820940912
+     0.008633227589035983
+    -0.006427442366270633
+      -0.1018570091925459
+       0.4281037933816986
+ 6.78e+10    
+       0.4291623213359755
+      -0.1018988932654242
+       0.4548118261873098
+    -0.006338631499786494
+     -0.05703287065218554
+        0.455035344997315
+     0.008690559231205191
+    -0.006380191108906636
+      -0.1020060268587531
+       0.4284264290228668
+ 6.79e+10    
+       0.4294834425571574
+      -0.1020473501834774
+       0.4552390310434479
+    -0.006290641169600212
+     -0.05717722429961556
+       0.4554630740278501
+     0.008747947185123017
+    -0.006332537364549024
+      -0.1021549099429652
+       0.4287479821242703
+ 6.8e+10     
+       0.4298034653503719
+      -0.1021956705574469
+       0.4556652987086001
+    -0.006242247477957911
+     -0.05732186491372929
+       0.4558898697096139
+     0.008805394133711494
+     -0.00628448076105692
+      -0.1023036617945351
+       0.4290684543062773
+ 6.81e+10    
+       0.4301223910465366
+       -0.102343857749199
+       0.4560906297154161
+    -0.006193450062046182
+     -0.05746679370809459
+        0.456315732605677
+     0.008862902813727728
+    -0.006236020930294541
+      -0.1024522858520177
+       0.4293878472304166
+ 6.82e+10    
+       0.4304402210137893
+      -0.1024919152095225
+       0.4565150246360517
+    -0.006144248562905985
+     -0.05761201190711777
+       0.4567406633185905
+     0.008920476015378676
+     -0.00618715750799626
+      -0.1026007856437134
+       0.4297061625996708
+ 6.83e+10    
+       0.4307569566577628
+      -0.1026398464786643
+        0.456938484082491
+    -0.006094642625295216
+     -0.05775752074611409
+       0.4571646624907088
+     0.008978116581923989
+    -0.006137890133629325
+      -0.1027491647882063
+       0.4300234021587644
+ 6.84e+10    
+       0.4310725994218515
+      -0.1027876551868569
+       0.4573610087068673
+    -0.006044631897549261
+     -0.05790332147137927
+       0.4575877308045117
+     0.009035827409266291
+    -0.006088218450253499
+       -0.102897426994898
+       0.4303395676944486
+ 6.85e+10    
+       0.4313871507874805
+      -0.1029353450548457
+       0.4577825992017829
+    -0.005994216031438576
+     -0.05804941534026294
+       0.4580098689829294
+     0.009093611445529625
+    -0.006038142104378235
+      -0.1030455760645393
+       0.4306546610357917
+ 6.86e+10    
+       0.4317006122743723
+      -0.1030829198944094
+       0.4582032563006255
+    -0.005943394682023295
+     -0.05819580362124128
+       0.4584310777896559
+     0.009151471690625645
+    -0.005987660745817266
+      -0.1031936158897536
+       0.4309686840544557
+ 6.87e+10    
+       0.4320129854408102
+      -0.1032303836088765
+       0.4586229807778848
+    -0.005892167507506025
+     -0.05834248759399268
+       0.4588513580294708
+     0.009209411195808254
+    -0.005936774027540297
+      -0.1033415504555606
+       0.4312816386649845
+ 6.88e+10    
+       0.4323242718839017
+      -0.1033777401936379
+       0.4590417734494657
+    -0.005840534169081173
+       -0.058489468549473
+       0.4592707105485537
+     0.009267433063215978
+    -0.005885481605522307
+      -0.1034893838398918
+         0.43159352682508
+ 6.89e+10    
+       0.4326344732398387
+      -0.1035249937366551
+       0.4594596351730006
+    -0.005788494330782134
+     -0.05863674778999294
+       0.4596891362347945
+     0.009325540445403051
+    -0.005833783138590074
+      -0.1036371202141027
+       0.4319043505358791
+ 6.9e+10     
+       0.4329435911841575
+      -0.1036721484189631
+       0.4598765668481587
+    -0.005736047659325814
+     -0.05878432662929576
+       0.4601066360181105
+     0.009383736544858854
+    -0.005781678288266214
+      -0.1037847638434821
+       0.4322141118422334
+ 6.91e+10    
+       0.4332516274319952
+       -0.103819208515169
+       0.4602925694169527
+    -0.005683193823954501
+     -0.05893220639263628
+       0.4605232108707522
+     0.009442024613515622
+    -0.005729166718610321
+      -0.1039323190877543
+       0.4325228128329797
+ 6.92e+10    
+       0.4335585837383437
+      -0.1039661783939464
+       0.4607076438640476
+    -0.005629932496275305
+     -0.05908038841686103
+       0.4609388618076122
+     0.009500407952245295
+    -0.005676248096058159
+      -0.1040797904015778
+       0.4328304556412123
+ 6.93e+10    
+       0.4338644618983041
+      -0.1041130625185246
+       0.4611217912170626
+    -0.005576263350096682
+     -0.05922887405048964
+       0.4613535898865293
+     0.009558889910344568
+    -0.005622922089257587
+      -0.1042271823350397
+        0.433137042444554
+ 6.94e+10    
+       0.4341692637473379
+      -0.1042598654471737
+       0.4615350125468715
+    -0.005522186061263313
+     -0.05937766465379632
+       0.4617673962085945
+     0.009617473885009713
+    -0.005569188368902489
+      -0.1043744995341448
+       0.4334425754654215
+ 6.95e+10    
+       0.4344729911615139
+      -0.1044065918336836
+       0.4619473089679058
+    -0.005467700307487104
+     -0.05952676159889433
+       0.4621802819184523
+     0.009676163320799271
+    -0.005515046607563721
+      -0.1045217467413001
+       0.4337470569712942
+ 6.96e+10    
+       0.4347756460577573
+      -0.1045532464278405
+       0.4623586816384496
+    -0.005412805768177232
+     -0.05967616626981941
+       0.4625922482045981
+     0.009734961709087239
+    -0.005460496479518082
+      -0.1046689287957943
+       0.4340504892749711
+ 6.97e+10    
+       0.4350772303940915
+      -0.1046998340758954
+       0.4627691317609349
+    -0.005357502124266449
+     -0.05982588006261551
+        0.463003296299677
+      0.00979387258750433
+    -0.005405537660574276
+      -0.1048160506342727
+       0.4343528747348391
+ 6.98e+10    
+       0.4353777461698824
+      -0.1048463597210307
+       0.4631786605822377
+    -0.005301789058035741
+     -0.05997590438542168
+       0.4634134274807797
+     0.009852899539369612
+    -0.005350169827896769
+      -0.1049631172912072
+       0.4346542157551251
+ 6.99e+10    
+       0.4356771954260767
+      -0.1049928284038197
+       0.4635872693939636
+    -0.005245666252936243
+     -0.06012624065855876
+       0.4638226430697341
+     0.009912046193111257
+    -0.005294392659827174
+      -0.1051101338993613
+       0.4349545147861562
+ 7e+10       
+        0.435975580245442
+      -0.1051392452626825
+       0.4639949595327433
+    -0.005189133393408644
+     -0.06027689031461914
+       0.4642309444333952
+     0.009971316221677054
+    -0.005238205835702979
+      -0.1052571056902485
+       0.4352537743246102
* NOTE: Solution at 1e+08 Hz used as DC point.

.model c_m4lines_HFSS_W_1 sp N=4 SPACING=nonuniform VALTYPE=real
+ INTERPOLATION=spline
+ INFINITY =
+    7.938621322074103e-11
+   -2.234686778922564e-11
+    8.350721157248263e-11
+   -1.872746540418529e-12
+   -1.142445181304755e-11
+    8.352938776572516e-11
+   -2.203335273976321e-13
+   -1.872043010176729e-12
+   -2.235002713338225e-11
+     7.92698254841625e-11
+ DATA = 700
+ 0           
+    8.640174920590117e-11
+    -2.14416090728894e-11
+    8.793408763567512e-11
+   -8.389673395611541e-13
+   -1.021175218891604e-11
+    8.796128153242538e-11
+   -3.023047060529615e-13
+   -8.359493564182524e-13
+   -2.144637104119777e-11
+    8.625786243188311e-11
+ 2e+08       
+    8.579356517807833e-11
+   -2.133018481287351e-11
+    8.732273804978702e-11
+   -8.409745571171349e-13
+   -1.015945392081564e-11
+    8.734928774723289e-11
+   -3.017209077407336e-13
+   -8.379727382415652e-13
+   -2.133396863163589e-11
+    8.565048805585838e-11
+ 3e+08       
+    8.543439129147498e-11
+   -2.125919358636875e-11
+    8.696147697909173e-11
+   -8.388714817469942e-13
+   -1.013212095931011e-11
+    8.698809761386621e-11
+   -3.016053761501185e-13
+   -8.358583481642005e-13
+   -2.126333912016844e-11
+    8.529262847560166e-11
+ 4e+08       
+     8.51973785006239e-11
+   -2.121611624896911e-11
+    8.672397360039697e-11
+   -8.370576263106825e-13
+    -1.01144905578764e-11
+    8.675056048629885e-11
+   -3.015461469017349e-13
+   -8.340441696890575e-13
+   -2.122041112324275e-11
+    8.505609369460387e-11
+ 5e+08       
+    8.501308142501136e-11
+   -2.118240268346723e-11
+    8.653926817497166e-11
+   -8.358747223385644e-13
+   -1.009992154090721e-11
+    8.656576400727495e-11
+   -3.012893316516853e-13
+   -8.328633203687275e-13
+   -2.118669760698499e-11
+    8.487204370126886e-11
+ 6e+08       
+    8.485906137203432e-11
+    -2.11533346653181e-11
+    8.638463937856391e-11
+   -8.349758688101932e-13
+   -1.008711758231931e-11
+    8.641104847680747e-11
+   -3.008173216221576e-13
+   -8.319664423778381e-13
+   -2.115758882075701e-11
+     8.47182727872951e-11
+ 7e+08       
+    8.472695307073616e-11
+   -2.112780632516672e-11
+    8.625179551406494e-11
+   -8.341174077938374e-13
+   -1.007578659555687e-11
+    8.627813731849719e-11
+   -3.001762091430381e-13
+   -8.311096585892238e-13
+   -2.113201709725078e-11
+     8.45864327515991e-11
+ 8e+08       
+    8.461229945786495e-11
+   -2.110531332881669e-11
+    8.613639890603737e-11
+   -8.331937424130681e-13
+   -1.006572106061007e-11
+    8.616268716773436e-11
+   -2.994151589074017e-13
+   -8.301876066807383e-13
+   -2.110948556650975e-11
+    8.447203040662894e-11
+ 9e+08       
+    8.451184222347195e-11
+   -2.108535962900842e-11
+    8.603526482545168e-11
+   -8.321766378163135e-13
+    -1.00566835807289e-11
+    8.606150428414358e-11
+    -2.98570621181589e-13
+   -8.291723195167683e-13
+   -2.108949872180673e-11
+    8.437178184932172e-11
+ 1e+09       
+    8.442288424772558e-11
+   -2.106742960264604e-11
+    8.594571214091148e-11
+   -8.310706423844269e-13
+    -1.00484331775308e-11
+    8.597190206687965e-11
+   -2.976659995362326e-13
+   -8.280685677340599e-13
+   -2.107154255125035e-11
+    8.428298725200001e-11
+ 1.1e+09     
+     8.43467868730977e-11
+    -2.10565228623004e-11
+    8.586308826004625e-11
+   -8.281628259677012e-13
+   -1.003958634525061e-11
+    8.588917790565399e-11
+   -2.960355782910471e-13
+    -8.25189830716901e-13
+   -2.106047083897488e-11
+    8.420677187963953e-11
+ 1.2e+09     
+    8.427560112040294e-11
+   -2.104531648908617e-11
+    8.578861755273247e-11
+   -8.258107749972172e-13
+   -1.003110455660544e-11
+    8.581461431009167e-11
+   -2.943374349957208e-13
+   -8.228623551389135e-13
+   -2.104911734365513e-11
+    8.413546455588259e-11
+ 1.3e+09     
+     8.42091616663341e-11
+   -2.103391629169333e-11
+    8.572096557110643e-11
+    -8.23910114686463e-13
+   -1.002299692517252e-11
+    8.574687619515703e-11
+   -2.925778086449991e-13
+   -8.209814938667681e-13
+   -2.103758862656038e-11
+    8.406890735365205e-11
+ 1.4e+09     
+    8.414718833313966e-11
+    -2.10224124183306e-11
+    8.565902860698295e-11
+   -8.223749517380232e-13
+   -1.001524287917462e-11
+    8.568485988398318e-11
+    -2.90760460813667e-13
+   -8.194611942612129e-13
+   -2.102597484440859e-11
+     8.40068265529164e-11
+ 1.5e+09     
+    8.408935010925876e-11
+   -2.101087923387924e-11
+    8.560191245326208e-11
+   -8.211345504708737e-13
+   -1.000781060000423e-11
+    8.562767142527594e-11
+   -2.888883548318776e-13
+   -8.182306493311775e-13
+   -2.101434981594957e-11
+     8.39488962336872e-11
+ 1.6e+09     
+     8.40353038819955e-11
+   -2.099937662633938e-11
+    8.554889937433408e-11
+   -8.201301960001971e-13
+   -1.000066620488537e-11
+    8.557459332286059e-11
+   -2.869646325365739e-13
+   -8.172311477916213e-13
+   -2.100277248311014e-11
+    8.389477687333485e-11
+ 1.7e+09     
+    8.398471638884087e-11
+    -2.09879518897071e-11
+    8.549941457564891e-11
+   -8.193124118802404e-13
+   -9.993778051297988e-12
+    8.552505089392479e-11
+   -2.849931483163632e-13
+   -8.164132880334446e-13
+   -2.099128892074878e-11
+    8.384413736389615e-11
+ 1.8e+09     
+    8.393727555926306e-11
+   -2.097664171934448e-11
+    8.545299660823854e-11
+   -8.186385935626231e-13
+   -9.987118534804766e-12
+    8.547858263831369e-11
+   -2.829787324064353e-13
+   -8.157346146746119e-13
+   -2.097993443536364e-11
+    8.379666653690576e-11
+ 1.9e+09     
+    8.389269543049556e-11
+   -2.096547409245719e-11
+    8.540927291211442e-11
+   -8.180710652131057e-13
+   -9.980664634545427e-12
+    8.543481578756385e-11
+   -2.809272895364934e-13
+   -8.151576826202957e-13
+   -2.096873552814151e-11
+    8.375207831420818e-11
+ 2e+09       
+    8.385071734239634e-11
+   -2.095446993710375e-11
+    8.536794030843047e-11
+   -8.175755431437786e-13
+   -9.974397854915927e-12
+    8.539344682180946e-11
+   -2.788457941687409e-13
+   -8.146485294207177e-13
+   -2.095771162804384e-11
+    8.371011314570396e-11
+ 2.1e+09     
+    8.381110909779752e-11
+   -2.094364456079859e-11
+     8.53287497440674e-11
+   -8.171199805780336e-13
+   -9.968303889455178e-12
+    8.535422624558459e-11
+   -2.767422149456995e-13
+   -8.141755283079569e-13
+    -2.09468765682861e-11
+    8.367053739410404e-11
+ 2.2e+09     
+     8.37736631067195e-11
+   -2.093300884264838e-11
+    8.529149448992127e-11
+   -8.166737671497549e-13
+   -9.962372164147643e-12
+    8.531694681701685e-11
+   -2.746253838968883e-13
+    -8.13708593099877e-13
+   -2.093623981259313e-11
+    8.363314167187041e-11
+ 2.3e+09     
+    8.373819410985685e-11
+   -2.092257020770033e-11
+    8.525600105809871e-11
+   -8.162072571927939e-13
+   -9.956595331085987e-12
+    8.528143449241183e-11
+   -2.725048168294584e-13
+   -8.132187069869776e-13
+   -2.092580745242712e-11
+    8.359773872134086e-11
+ 2.4e+09     
+    8.370453681623286e-11
+   -2.091233340787329e-11
+    8.522212222165464e-11
+   -8.156916003909332e-13
+   -9.950968741367886e-12
+    8.524754146874447e-11
+   -2.703904876636825e-13
+   -8.126777470272222e-13
+   -2.091558300200351e-11
+    8.356416117382966e-11
+ 2.5e+09     
+    8.367254363323448e-11
+    -2.09023011352358e-11
+    8.518973164409307e-11
+   -8.150988451068987e-13
+   -9.945489907704494e-12
+    8.521514083128877e-11
+   -2.682925595980215e-13
+   -8.120585734028408e-13
+   -2.090556801909052e-11
+    8.353225936963638e-11
+ 2.6e+09     
+    8.364208257517254e-11
+   -2.089247449290517e-11
+    8.515871973532149e-11
+   -8.144022782200718e-13
+   -9.940157961492351e-12
+    8.518412242362024e-11
+   -2.662210787077826e-13
+   -8.113353467103044e-13
+   -2.089576257877927e-11
+    8.350189933001299e-11
+ 2.7e+09     
+    8.361303538379102e-11
+   -2.088285334762375e-11
+    8.512899044068244e-11
+   -8.135769560894266e-13
+   -9.934973109995162e-12
+     8.51543896473313e-11
+   -2.641856399157917e-13
+   -8.104840282581321e-13
+   -2.088616562581853e-11
+    8.347296091961255e-11
+ 2.8e+09     
+    8.358529586497227e-11
+   -2.087343658662818e-11
+    8.510045874060466e-11
+   -8.126003706864111e-13
+   -9.929936103268278e-12
+    8.512585696969518e-11
+   -2.621950402773749e-13
+   -8.094830088297163e-13
+   -2.087677522927202e-11
+    8.344533620841709e-11
+ 2.9e+09     
+    8.355876843055214e-11
+   -2.086422229989436e-11
+    8.507304869301057e-11
+   -8.114531850225188e-13
+   -9.925047725259528e-12
+    8.509844797197123e-11
+   -2.602569392203373e-13
+   -8.083138025112066e-13
+    -2.08675887613484e-11
+    8.341892802621142e-11
+ 3e+09       
+    8.353336682686228e-11
+   -2.085520790717069e-11
+    8.504669189201685e-11
+   -8.101199650800886e-13
+   -9.920308327521527e-12
+    8.507209381228789e-11
+   -2.583775487954478e-13
+   -8.069617361564391e-13
+   -2.085860302025754e-11
+    8.339364869469498e-11
+ 3.1e+09     
+    8.350901302891646e-11
+   -2.084639024728118e-11
+     8.50213262475852e-11
+   -8.085898337677164e-13
+    -9.91571742600566e-12
+    8.504673200800132e-11
+    -2.56561378257628e-13
+   -8.054165639061087e-13
+   -2.084981431475978e-11
+    8.336941891895915e-11
+ 3.2e+09     
+    8.348563627904544e-11
+    -2.08377656448696e-11
+    8.499689501403472e-11
+    -8.06856977569252e-13
+   -9.911273380748351e-12
+    8.502230546557291e-11
+   -2.548110558155666e-13
+   -8.036729413463831e-13
+   -2.084121852559902e-11
+    8.334616681934766e-11
+ 3.3e+09     
+    8.346317225011358e-11
+   -2.082932996703402e-11
+    8.497334601265863e-11
+   -8.049209490566221e-13
+   -9.906973174674848e-12
+    8.499876170328194e-11
+   -2.531272459749971e-13
+   -8.017307058436758e-13
+   -2.083281115621012e-11
+    8.332382708551703e-11
+ 3.4e+09     
+    8.344156231550942e-11
+   -2.082107867922011e-11
+    8.495063100659096e-11
+   -8.027867274778783e-13
+   -9.902812301546719e-12
+     8.49760522249848e-11
+   -2.515086738815035e-13
+   -7.995949275497881e-13
+   -2.082458738201409e-11
+    8.330234023612577e-11
+ 3.5e+09     
+    8.342075291048813e-11
+   -2.081300690648183e-11
+    8.492870519568585e-11
+   -8.004645230871731e-13
+   -9.898784765074136e-12
+    8.495413201278549e-11
+   -2.499522592489527e-13
+   -7.972757175833067e-13
+   -2.081654210442079e-11
+    8.328165196959121e-11
+ 3.6e+09     
+    8.340069497186114e-11
+   -2.080510950303099e-11
+    8.490752680636543e-11
+    -7.97969335709457e-13
+   -9.894883182561917e-12
+    8.493295911373987e-11
+   -2.484533529950076e-13
+   -7.947878031510941e-13
+   -2.080867001256672e-11
+    8.326171259346187e-11
+ 3.7e+09     
+    8.338134344528164e-11
+   -2.079738113015868e-11
+    8.488705675681445e-11
+    -7.95320300851444e-13
+    -9.89109897843455e-12
+    8.491249430119443e-11
+   -2.470060608791506e-13
+   -7.921499007762461e-13
+   -2.080096565307735e-11
+    8.324247652197642e-11
+ 3.8e+09     
+    8.336265685135723e-11
+   -2.078981634037557e-11
+    8.486725838202209e-11
+   -7.925398744905056e-13
+   -9.887422646725285e-12
+    8.489270079553441e-11
+   -2.456036314048512e-13
+   -7.893839355876449e-13
+   -2.079342350598018e-11
+    8.322390183317244e-11
+ 3.9e+09     
+     8.33445969034289e-11
+    -2.07824096641374e-11
+    8.484809720635924e-11
+   -7.896529184711778e-13
+    -9.88384405788997e-12
+     8.48735440323116e-11
+   -2.442388808144999e-13
+   -7.865141649131792e-13
+   -2.078603806344786e-11
+    8.320594987841278e-11
+ 4e+09       
+    8.332712817110979e-11
+    -2.07751556948483e-11
+     8.48295407538712e-11
+   -7.866857514752294e-13
+   -9.880352784412325e-12
+    8.485499146820462e-11
+   -2.429046265164639e-13
+   -7.835662674981746e-13
+   -2.077880390736361e-11
+    8.318858493836503e-11
+ 4.1e+09     
+    8.331021778457777e-11
+   -2.076804916789404e-11
+    8.481155838845545e-11
+   -7.836652263792309e-13
+   -9.876938421409246e-12
+    8.483701241720172e-11
+    -2.41594101603732e-13
+   -7.805664560245552e-13
+   -2.077171578170797e-11
+    8.317177392035016e-11
+ 4.2e+09     
+    8.329383517524265e-11
+   -2.076108503009252e-11
+    8.479412117769679e-11
+   -7.806178850424695e-13
+   -9.873590882252177e-12
+    8.481957791093498e-11
+   -2.403013267434422e-13
+   -7.775406616591851e-13
+   -2.076476865632123e-11
+    8.315548609259007e-11
+ 4.3e+09     
+     8.32779518488296e-11
+   -2.075425849694954e-11
+    8.477720177543095e-11
+   -7.775692283272442e-13
+   -9.870300654303922e-12
+    8.480266057832507e-11
+   -2.390214209026477e-13
+   -7.745138270699772e-13
+   -2.075795777950634e-11
+    8.313969285132128e-11
+ 4.4e+09     
+    8.326254118721959e-11
+   -2.074756509626167e-11
+    8.476077431916846e-11
+   -7.745431246587499e-13
+   -9.867059005408072e-12
+    8.478623454068717e-11
+   -2.377508383429134e-13
+   -7.715093307742125e-13
+   -2.075127871800734e-11
+    8.312436751705781e-11
+ 4.5e+09     
+    8.324757827562424e-11
+   -2.074100069772934e-11
+    8.474481433936865e-11
+   -7.715613665979386e-13
+   -9.863858137047949e-12
+     8.47702753192519e-11
+    -2.36487525362525e-13
+   -7.685485526126467e-13
+   -2.074472738394836e-11
+    8.310948515654179e-11
+ 4.6e+09     
+    8.323303975189616e-11
+   -2.073456152919983e-11
+    8.472929867823983e-11
+   -7.686433730991402e-13
+   -9.860691284598886e-12
+    8.475475975270307e-11
+   -2.352309958517864e-13
+   -7.656505788866734e-13
+   -2.073830004922832e-11
+    8.309502242716312e-11
+ 4.7e+09     
+    8.321890367501613e-11
+   -2.072824418087668e-11
+    8.471420541628067e-11
+   -7.658060261080592e-13
+   -9.857552768547585e-12
+    8.473966592286036e-11
+   -2.339823295079998e-13
+   -7.628320369906219e-13
+   -2.073199334855865e-11
+    8.308095744087725e-11
+ 4.8e+09     
+    8.320514941005949e-11
+    -2.07220455992893e-11
+    8.469951380520837e-11
+   -7.630636241308486e-13
+   -9.854438002867819e-12
+    8.472497308704347e-11
+   -2.327441003565363e-13
+   -7.601070434531788e-13
+   -2.072580427278121e-11
+    8.306726964491829e-11
+ 4.9e+09     
+    8.319175752722661e-11
+   -2.071596307302764e-11
+    8.468520420622796e-11
+   -7.604279321566447e-13
+   -9.851343467999696e-12
+    8.471066161598935e-11
+   -2.315202459991144e-13
+   -7.574872460013266e-13
+   -2.071973015432653e-11
+    8.305393971688959e-11
+ 5e+09       
+    8.317870971281685e-11
+   -2.070999421226018e-11
+    8.467125803284704e-11
+   -7.579083063817382e-13
+   -9.848266656259631e-12
+    8.469671293643868e-11
+   -2.303158897979714e-13
+   -7.549819391698383e-13
+   -2.071376864670302e-11
+    8.304094947210472e-11
+ 5.1e+09     
+    8.316598869031374e-11
+   -2.070413692391864e-11
+    8.465765769761337e-11
+   -7.555118729854027e-13
+    -9.84520599722711e-12
+    8.468310947770781e-11
+    -2.29137129090247e-13
+   -7.525982335740065e-13
+   -2.070791769979729e-11
+    8.302828178133877e-11
+ 5.2e+09     
+    8.315357815002914e-11
+    -2.06983893842054e-11
+    8.464438656228085e-11
+    -7.53243742179206e-13
+   -9.842160769931171e-12
+    8.466983462170295e-11
+   -2.279908026144303e-13
+   -7.503412607124395e-13
+   -2.070217553256325e-11
+    8.301592049742602e-11
+ 5.3e+09     
+    8.314146268600067e-11
+   -2.069275000980549e-11
+    8.463142889100558e-11
+   -7.511072413917803e-13
+   -9.839131007687456e-12
+    8.465687265594662e-11
+   -2.268842497333865e-13
+   -7.482143976006246e-13
+   -2.069654060442565e-11
+    8.300385038938559e-11
+ 5.4e+09     
+    8.312962773906538e-11
+   -2.068721742890317e-11
+    8.461876980624155e-11
+   -7.491041543669228e-13
+   -9.836117400365886e-12
+    8.464420872926747e-11
+   -2.258250728754499e-13
+   -7.462194982742112e-13
+   -2.069101158646195e-11
+    8.299205708297902e-11
+ 5.5e+09     
+    8.311805954521732e-11
+   -2.068179045283539e-11
+    8.460639524705884e-11
+   -7.472349558550189e-13
+   -9.833121197811067e-12
+    8.463182880986402e-11
+   -2.248209130136789e-13
+   -7.443571219641143e-13
+   -2.068558733317268e-11
+    8.298052700679099e-11
+ 5.6e+09     
+    8.310674508851859e-11
+   -2.067646804897899e-11
+    8.459429192964472e-11
+   -7.454990342818355e-13
+   -9.830144117162473e-12
+    8.461971964550867e-11
+   -2.238792460971187e-13
+   -7.426267503441456e-13
+   -2.068026685542988e-11
+    8.296924734308576e-11
+ 5.7e+09     
+     8.30956720579588e-11
+   -2.067124931527206e-11
+    8.458244730978532e-11
+   -7.438948971678478e-13
+   -9.827188255969483e-12
+    8.460786872568548e-11
+    -2.23007206276729e-13
+   -7.410269885734807e-13
+   -2.067504929500078e-11
+    8.295820598281467e-11
+ 5.8e+09     
+    8.308482880776482e-11
+   -2.066613345661267e-11
+    8.457084954715002e-11
+   -7.424203560992548e-13
+   -9.824256012285885e-12
+    8.459626424549887e-11
+   -2.222114396704024e-13
+   -7.395557468383245e-13
+   -2.066993390089613e-11
+    8.294739148426145e-11
+ 5.9e+09     
+    8.307420432074112e-11
+   -2.066111976325794e-11
+    8.455948747122555e-11
+   -7.410726897044789e-13
+   -9.821350012356642e-12
+    8.458489507120574e-11
+   -2.214979904121151e-13
+   -7.382104007289779e-13
+   -2.066492000767228e-11
+    8.293679303488783e-11
+ 6e+09       
+    8.306378817428843e-11
+   -2.065620759125908e-11
+     8.45483505487702e-11
+   -7.398487843821565e-13
+   -9.818473046071573e-12
+    8.457375070725162e-11
+   -2.208722189388819e-13
+   -7.369879300733638e-13
+   -2.066000701573253e-11
+     8.29264004160161e-11
+ 6.1e+09     
+    8.305357050880051e-11
+     -2.0651396344906e-11
+     8.45374288526747e-11
+   -7.387452534921371e-13
+   -9.815628010037857e-12
+    8.456282126470759e-11
+   -2.203387509641124e-13
+   -7.358850368162056e-13
+      -2.065519437361e-11
+    8.291620397003158e-11
+ 6.2e+09     
+    8.304354199817823e-11
+   -2.064668546111399e-11
+    8.452671303213361e-11
+   -7.377585363990234e-13
+   -9.812817857899652e-12
+    8.455209743102164e-11
+   -2.199014544167509e-13
+   -7.348982432208522e-13
+   -2.065048156217415e-11
+    8.290619456983656e-11
+ 6.3e+09     
+    8.303369382223941e-11
+   -2.064207439565916e-11
+    8.451619428404551e-11
+   -7.368849791927793e-13
+   -9.810045557390665e-12
+    8.454157044101093e-11
+   -2.195634408081342e-13
+   -7.340239721176974e-13
+   -2.064586808067543e-11
+    8.289636359032069e-11
+ 6.4e+09     
+    8.302401764082743e-11
+    -2.06375626111547e-11
+    8.450586432557219e-11
+   -7.361208991458624e-13
+   -9.807314053528103e-12
+    8.453123204902951e-11
+   -2.193270870114888e-13
+   -7.332586111738171e-13
+   -2.064135343452691e-11
+    8.288670288164431e-11
+ 6.5e+09     
+    8.301450556945162e-11
+   -2.063314956665158e-11
+    8.449571536779594e-11
+   -7.354626350488566e-13
+   -9.804626237326436e-12
+    8.452107450226112e-11
+   -2.191940732660615e-13
+   -7.325985632523979e-13
+   -2.063693712471339e-11
+    8.287720474415749e-11
+ 6.6e+09     
+    8.300515015631112e-11
+   -2.062883470874639e-11
+    8.448574009042425e-11
+   -7.349065855275557e-13
+   -9.801984919416743e-12
+    8.451109051508646e-11
+   -2.191654333002623e-13
+   -7.320402849066275e-13
+   -2.063261863871445e-11
+    8.286786190480007e-11
+ 6.7e+09     
+    8.299594436057332e-11
+    -2.06246174640772e-11
+    8.447593161749347e-11
+   -7.344492373262127e-13
+   -9.799392807987039e-12
+    8.450127324448456e-11
+   -2.192416127455933e-13
+   -7.315803149454601e-13
+   -2.062839744282741e-11
+     8.28586674948479e-11
+ 6.8e+09     
+    8.298688153179913e-11
+   -2.062049723309436e-11
+    8.446628349403587e-11
+   -7.340871853680609e-13
+    -9.79685249050685e-12
+    8.449161626643073e-11
+   -2.194225324275818e-13
+   -7.312152948446769e-13
+   -2.062427297577858e-11
+    8.284961502888875e-11
+ 6.9e+09     
+    8.297795539041561e-11
+   -2.061647338499297e-11
+    8.445678966366869e-11
+   -7.338171462012492e-13
+   -9.794366418751615e-12
+    8.448211355325603e-11
+   -2.197076536141217e-13
+   -7.309419825830329e-13
+   -2.062024464351323e-11
+    8.284069838492696e-11
+ 7e+09       
+    8.296916000915631e-11
+   -2.061254525370117e-11
+    8.444744444707626e-11
+   -7.336359662236944e-13
+   -9.791936896701368e-12
+    8.447275945193773e-11
+   -2.200960428295389e-13
+   -7.307572612750123e-13
+   -2.061631181505868e-11
+    8.283191178552706e-11
+ 7.1e+09     
+    8.296048979539618e-11
+   -2.060871213482193e-11
+    8.443824252135456e-11
+   -7.335406258688516e-13
+   -9.789566070943215e-12
+    8.446354866328922e-11
+   -2.205864343639636e-13
+    -7.30658143766608e-13
+   -2.061247381935916e-11
+    8.282324977992163e-11
+ 7.2e+09     
+    8.295193947431875e-11
+   -2.060497328343066e-11
+    8.442917890018799e-11
+   -7.335282407341791e-13
+   -9.787255923259813e-12
+    8.445447622202334e-11
+   -2.211772890963884e-13
+    -7.30641774164319e-13
+   -2.060872994298607e-11
+    8.281470722701565e-11
+ 7.3e+09     
+    8.294350407286396e-11
+   -2.060132791263755e-11
+    8.442024891483766e-11
+   -7.335960604529556e-13
+   -9.785008265133644e-12
+    8.444553747766187e-11
+     -2.2186684868547e-13
+   -7.307054270902496e-13
+   -2.060507942863101e-11
+    8.280627927922902e-11
+ 7.4e+09     
+    8.293517890440739e-11
+   -2.059777519282721e-11
+    8.441144819591146e-11
+   -7.337414659490713e-13
+   -9.782824733937299e-12
+    8.443672807626416e-11
+   -2.226531845563777e-13
+   -7.308465052980486e-13
+   -2.060152147429504e-11
+    8.279796136712674e-11
+ 7.5e+09     
+    8.292695955413125e-11
+   -2.059431425149498e-11
+    8.440277265589745e-11
+   -7.339619655775338e-13
+   -9.780706790615885e-12
+    8.442804394295308e-11
+   -2.235342414197255e-13
+   -7.310625361493073e-13
+   -2.059805523309196e-11
+     8.27897491847897e-11
+ 7.6e+09     
+    8.291884186504975e-11
+   -2.059094417360386e-11
+    8.439421847243781e-11
+   -7.342551905366623e-13
+   -9.778655718696219e-12
+    8.441948126521253e-11
+   -2.245078753026358e-13
+   -7.313511673352589e-13
+   -2.059467981358938e-11
+    8.278163867588667e-11
+ 7.7e+09     
+    8.291082192465665e-11
+   -2.058766400239161e-11
+    8.438578207232266e-11
+   -7.346188898435958e-13
+   -9.776672624481151e-12
+    8.441103647693589e-11
+   -2.255718862561564e-13
+   -7.317101621349047e-13
+   -2.059139428061569e-11
+     8.27736260204101e-11
+ 7.8e+09     
+    8.290289605216548e-11
+   -2.058447274056305e-11
+    8.437746011618489e-11
+   -7.350509250874243e-13
+   -9.774758438305945e-12
+    8.440270624320086e-11
+   -2.267240460353344e-13
+   -7.321373944247276e-13
+   -2.058819765646697e-11
+    8.276570762204221e-11
+ 7.9e+09     
+    8.289506078631492e-11
+   -2.058136935180781e-11
+     8.43692494838778e-11
+   -7.355492651137914e-13
+   -9.772913916748523e-12
+    8.439448744575239e-11
+   -2.279621211356931e-13
+   -7.326308435947843e-13
+   -2.058508892245284e-11
+    8.275788009612102e-11
+ 8e+09       
+    8.288731287371565e-11
+   -2.057835276258861e-11
+    8.436114726051725e-11
+   -7.361119807478882e-13
+   -9.771139645696224e-12
+    8.438637716917017e-11
+   -2.292838916208295e-13
+   -7.331885894795856e-13
+   -2.058206702072505e-11
+    8.275014025817709e-11
+ 8.1e+09     
+    8.287964925771409e-11
+   -2.057542186415052e-11
+    8.435315072317059e-11
+   -7.367372396271834e-13
+   -9.769436044180177e-12
+    8.437837268770245e-11
+   -2.306871661982489e-13
+   -7.338088073765693e-13
+   -2.057913085633787e-11
+    8.274248511301475e-11
+ 8.2e+09     
+      8.2872067067753e-11
+   -2.057257551470572e-11
+    8.434525732817568e-11
+   -7.374233011885372e-13
+   -9.767803368894623e-12
+    8.437047145274487e-11
+   -2.321697940008303e-13
+   -7.344897631990123e-13
+   -2.057627929949395e-11
+    8.273491184431272e-11
+ 8.3e+09     
+    8.286456360920813e-11
+   -2.056981254175426e-11
+      8.4337464699074e-11
+   -7.381685118353555e-13
+   -9.766241719323622e-12
+    8.436267108094524e-11
+   -2.337296735161123e-13
+   -7.352298087905691e-13
+   -2.057351118793376e-11
+    8.272741780472123e-11
+ 8.4e+09     
+    8.285713635368056e-11
+   -2.056713174450276e-11
+    8.432977061513934e-11
+   -7.389713002976421e-13
+   -9.764751043400514e-12
+    8.435496934291507e-11
+   -2.353647590790222e-13
+   -7.360273774156238e-13
+   -2.057082532943121e-11
+    8.272000050643147e-11
+ 8.5e+09     
+    8.284978292972875e-11
+   -2.056453189635103e-11
+    8.432217300048764e-11
+   -7.398301731876884e-13
+    -9.76333114362898e-12
+    8.434736415252754e-11
+   -2.370730653108129e-13
+   -7.368809794304842e-13
+   -2.056822050436145e-11
+    8.271265761219784e-11
+ 8.6e+09     
+    8.284250111402093e-11
+   -2.056201174741603e-11
+    8.431466991374977e-11
+   -7.407437107492691e-13
+    -9.76198168359676e-12
+    8.433985355678453e-11
+   -2.388526698499257e-13
+   -7.377891981346516e-13
+   -2.056569546831215e-11
+    8.270538692679268e-11
+ 8.7e+09     
+    8.283528882289212e-11
+   -2.055957002706967e-11
+    8.430725953829159e-11
+    -7.41710562794486e-13
+   -9.760702194815602e-12
+    8.433243572623136e-11
+   -2.407017146826634e-13
+   -7.387506857973301e-13
+    -2.05632489547112e-11
+    8.269818638887303e-11
+ 8.8e+09     
+       8.282814410429e-11
+   -2.055720544646803e-11
+    8.429994017296422e-11
+   -7.427294448207213e-13
+   -9.759492083823131e-12
+    8.432510894590299e-11
+    -2.42618406343612e-13
+      -7.397641598537e-13
+   -2.056087967744868e-11
+    8.269105406324219e-11
+ 8.9e+09     
+    8.282106513009367e-11
+    -2.05549167010532e-11
+    8.429271022336833e-11
+   -7.437991342993799e-13
+   -9.758350639485297e-12
+    8.431787160678059e-11
+    -2.44601015220154e-13
+   -7.408283992631289e-13
+   -2.055858633347284e-11
+    8.268398813348786e-11
+ 9e+09       
+    8.281405018879121e-11
+   -2.055270247301189e-11
+    8.428556819361357e-11
+   -7.449184671286236e-13
+   -9.757277040440022e-12
+    8.431072219774074e-11
+   -2.466478741615504e-13
+   -7.419422410230288e-13
+   -2.055636760534391e-11
+    8.267698689498108e-11
+ 9.1e+09     
+    8.280709767850315e-11
+   -2.055056143367773e-11
+    8.427851267855984e-11
+    -7.46086334242394e-13
+   -9.756270362626751e-12
+    8.430365929797886e-11
+   -2.487573765626942e-13
+   -7.431045768315937e-13
+   -2.055422216373052e-11
+    8.267004874821883e-11
+ 9.2e+09     
+    8.280020610033534e-11
+   -2.054849224586487e-11
+    8.427154235651956e-11
+   -7.473016783690206e-13
+   -9.755329586848789e-12
+    8.429668156988819e-11
+   -2.509279740649792e-13
+   -7.443143498937261e-13
+   -2.055214866983746e-11
+    8.266317219249594e-11
+ 9.3e+09     
+    8.279337405205151e-11
+   -2.054649356612476e-11
+    8.426465598240559e-11
+   -7.485634909338055e-13
+   -9.754453606319402e-12
+    8.428978775237465e-11
+   -2.531581739924908e-13
+   -7.455705518646506e-13
+   -2.055014577775463e-11
+    8.265635581989135e-11
+ 9.4e+09     
+    8.278660022205178e-11
+   -2.054456404691857e-11
+    8.425785238130876e-11
+   -7.498708090999989e-13
+   -9.753641234146741e-12
+    8.428297665459219e-11
+   -2.554465366202721e-13
+   -7.468722199274702e-13
+   -2.054821213671911e-11
+     8.26495983095552e-11
+ 9.5e+09     
+     8.27798833836446e-11
+   -2.054270233869906e-11
+    8.425113044248571e-11
+     -7.5122271294431e-13
+   -9.752891210715776e-12
+    8.427624715007901e-11
+   -2.577916723530592e-13
+    -7.48218434000321e-13
+   -2.054634639328483e-11
+    8.264289842228319e-11
+ 9.6e+09     
+    8.277322238960132e-11
+   -2.054090709189819e-11
+    8.424448911374133e-11
+   -7.526183227625795e-13
+   -9.752202210930072e-12
+    8.426959817127577e-11
+   -2.601922388770835e-13
+   -7.496083140702194e-13
+   -2.054454719339418e-11
+     8.26362549953658e-11
+ 9.7e+09     
+    8.276661616698273e-11
+   -2.053917695881764e-11
+    8.423792739618958e-11
+   -7.540567965030841e-13
+   -9.751572851280487e-12
+    8.426302870441232e-11
+   -2.626469383339731e-13
+   -7.510410176506587e-13
+   -2.054281318434958e-11
+    8.262966693770093e-11
+ 9.8e+09     
+    8.276006371222585e-11
+   -2.053751059542005e-11
+    8.423144433937425e-11
+   -7.555373273234689e-13
+   -9.751001696711713e-12
+    8.425653778474177e-11
+   -2.651545145547818e-13
+   -7.525157373602917e-13
+   -2.054114301668164e-11
+    8.262313322515651e-11
+ 9.9e+09     
+    8.275356408648126e-11
+   -2.053590666302064e-11
+    8.422503903673533e-11
+   -7.570591412694256e-13
+   -9.750487267261814e-12
+    8.425012449210827e-11
+   -2.677137503824256e-13
+   -7.540316986204046e-13
+   -2.053953534591417e-11
+    8.261665289617505e-11
+ 1e+10       
+    8.274711641119144e-11
+   -2.053436382987935e-11
+    8.421871062140328e-11
+   -7.586214950716547e-13
+   -9.750028044454334e-12
+    8.424378794683085e-11
+    -2.70323465103354e-13
+   -7.555881574687884e-13
+   -2.053798883422521e-11
+    8.261022504760704e-11
+ 1.01e+10    
+    8.274071986389953e-11
+   -2.053288077269409e-11
+    8.421245826230615e-11
+    -7.60223674059132e-13
+   -9.749622477425926e-12
+     8.42375273058883e-11
+   -2.729825120026781e-13
+    -7.57184398487321e-13
+    -2.05365021520051e-11
+    8.260384883076423e-11
+ 1.02e+10    
+    8.273437367428003e-11
+    -2.05314561779968e-11
+    8.420628116057298e-11
+    -7.61864990184938e-13
+   -9.749268988776634e-12
+    8.423134175938949e-11
+   -2.756897760521039e-13
+   -7.588197328411404e-13
+   -2.053507397931318e-11
+    8.259752344768416e-11
+ 1.03e+10    
+    8.272807712038279e-11
+   -2.053008874345457e-11
+    8.420017854622046e-11
+   -7.635447801630466e-13
+   -9.748965980133273e-12
+    8.422523052731366e-11
+   -2.784441717354598e-13
+   -7.604934964265266e-13
+   -2.053370300723497e-11
+    8.259124814759471e-11
+ 1.04e+10    
+    8.272182952508031e-11
+   -2.052877717907774e-11
+    8.419414967510482e-11
+   -7.652624037117355e-13
+   -9.748711837419788e-12
+    8.421919285650754e-11
+   -2.812446410139515e-13
+    -7.62205048124552e-13
+   -2.053238793914207e-11
+    8.258502222357092e-11
+ 1.05e+10    
+    8.271563025271107e-11
+   -2.052752020833834e-11
+    8.418819382612807e-11
+   -7.670172419014405e-13
+   -9.748504935831349e-12
+    8.421322801792489e-11
+   -2.840901514300916e-13
+   -7.639537681577954e-13
+   -2.053112749185852e-11
+     8.25788450093771e-11
+ 1.06e+10    
+    8.270947870591124e-11
+   -2.052631656920185e-11
+    8.418231029868188e-11
+   -7.688086956030048e-13
+    -9.74834364451171e-12
+    8.420733530409365e-11
+    -2.86979694347877e-13
+   -7.657390565465514e-13
+   -2.052992039673556e-11
+    8.257271587648275e-11
+ 1.07e+10    
+    8.270337432262482e-11
+   -2.052516501507526e-11
+    8.417649841031721e-11
+   -7.706361840334705e-13
+    -9.74822633093599e-12
+    8.420151402680047e-11
+   -2.899122833248328e-13
+   -7.675603316614672e-13
+   -2.052876540063935e-11
+    8.256663423124824e-11
+ 1.08e+10    
+    8.269731657328734e-11
+   -2.052406431567521e-11
+    8.417075749462493e-11
+    -7.72499143394965e-13
+   -9.748151365002763e-12
+    8.419576351497745e-11
+   -2.928869526109791e-13
+   -7.694170288687409e-13
+   -2.052766126685444e-11
+    8.256059951226955e-11
+ 1.09e+10    
+    8.269130495817304e-11
+   -2.052301325781966e-11
+    8.416508689931695e-11
+   -7.743970256037441e-13
+   -9.748117122841719e-12
+     8.41900831127804e-11
+   -2.959027557685591e-13
+   -7.713085992645234e-13
+     -2.0526606775907e-11
+    8.255461118787754e-11
+ 1.1e+10     
+    8.268533900490068e-11
+   -2.052201064614675e-11
+    8.415948598449442e-11
+   -7.763292971045878e-13
+    -9.74812199034446e-12
+    8.418447217784741e-11
+   -2.989587644063733e-13
+   -7.732345084944179e-13
+   -2.052560072631169e-11
+    8.254866875378305e-11
+ 1.11e+10    
+    8.267941826608984e-11
+   -2.052105530376412e-11
+    8.415395412108978e-11
+   -7.782954377675981e-13
+   -9.748164366426903e-12
+    8.417893007972492e-11
+   -3.020540670219185e-13
+   -7.751942356542155e-13
+    -2.05246419352454e-11
+    8.254277173086157e-11
+ 1.12e+10    
+    8.267354231716008e-11
+   -2.052014607283259e-11
+     8.41484906894748e-11
+   -7.802949398623328e-13
+   -9.748242666033796e-12
+    8.417345619845259e-11
+   -3.051877679446792e-13
+   -7.771872722682745e-13
+   -2.052372923915227e-11
+    8.253691966307196e-11
+ 1.13e+10    
+    8.266771075426937e-11
+    -2.05192818150877e-11
+    8.414309507822037e-11
+   -7.823273071063899e-13
+   -9.748355322895515e-12
+    8.416804992329578e-11
+   -3.083589863737845e-13
+     -7.7921312134108e-13
+   -2.052286149428333e-11
+    8.253111211550179e-11
+ 1.14e+10    
+    8.266192319238196e-11
+   -2.051846141230224e-11
+    8.413776668299914e-11
+   -7.843920537833361e-13
+   -9.748500792048575e-12
+    8.416271065161514e-11
+   -3.115668555035705e-13
+   -7.812712964784734e-13
+    -2.05220375771742e-11
+    8.252534867253409e-11
+ 1.15e+10    
+      8.2656179263462e-11
+   -2.051768376669363e-11
+    8.413250490562172e-11
+   -7.864887039268933e-13
+   -9.748677552131629e-12
+    8.415743778786536e-11
+   -3.148105217305359e-13
+   -7.833613210742242e-13
+   -2.052125638506476e-11
+    8.251962893612955e-11
+ 1.16e+10    
+    8.265047861478578e-11
+   -2.051694780127845e-11
+    8.412730915319436e-11
+   -7.886167905670235e-13
+   -9.748884107468228e-12
+    8.415223074271294e-11
+   -3.180891439355998e-13
+   -7.854827275586204e-13
+   -2.052051683626425e-11
+    8.251395252421884e-11
+ 1.17e+10    
+    8.264482090736762e-11
+   -2.051625246017854e-11
+    8.412217883739158e-11
+   -7.907758550344884e-13
+   -9.749118989948662e-12
+    8.414708893226458e-11
+    -3.21401892835785e-13
+   -7.876350567048538e-13
+    -2.05198178704642e-11
+    8.250831906919888e-11
+ 1.18e+10    
+    8.263920581449307e-11
+   -2.051559670888044e-11
+    8.411711337383356e-11
+    -7.92965446319863e-13
+   -9.749380760722257e-12
+    8.414201177739853e-11
+   -3.247479503997254e-13
+   -7.898178569899622e-13
+   -2.051915844900386e-11
+    8.250272821652988e-11
+ 1.19e+10    
+    8.263363302035482e-11
+    -2.05149795344515e-11
+    8.411211218155967e-11
+   -7.951851204837069e-13
+   -9.749668011711453e-12
+     8.41369987031896e-11
+   -3.281265093218704e-13
+   -7.920306840062884e-13
+   -2.051853755508959e-11
+    8.249717962342519e-11
+ 1.2e+10     
+     8.26281022187846e-11
+   -2.051439994571542e-11
+    8.410717468259106e-11
+   -7.974344401146243e-13
+   -9.749979366959031e-12
+    8.413204913842283e-11
+   -3.315367725501832e-13
+    -7.94273099920991e-13
+   -2.051795419397228e-11
+    8.249167295763257e-11
+ 1.21e+10    
+    8.262261311207876e-11
+   -2.051385697338953e-11
+    8.410230030157428e-11
+   -7.997129738316427e-13
+   -9.750313483818746e-12
+    8.412716251518472e-11
+   -3.349779528630278e-13
+   -7.965446729793949e-13
+   -2.051740739308434e-11
+    8.248620789629894e-11
+ 1.22e+10    
+     8.26171654099099e-11
+   -2.051334967018667e-11
+    8.409748846549845e-11
+   -8.020202958282862e-13
+   -9.750669053999992e-12
+    8.412233826852974e-11
+   -3.384492724906366e-13
+   -7.988449770498887e-13
+   -2.051689620214031e-11
+    8.248078412491715e-11
+ 1.23e+10    
+    8.261175882832146e-11
+   -2.051287711088293e-11
+    8.409273860347875e-11
+   -8.043559854550756e-13
+   -9.751044804475576e-12
+    8.411757583621196e-11
+   -3.419499627773573e-13
+   -8.011735912072217e-13
+   -2.051641969320193e-11
+    8.247540133634853e-11
+ 1.24e+10    
+    8.260639308879977e-11
+   -2.051243839235475e-11
+    8.408805014660152e-11
+   -8.067196268380131e-13
+   -9.751439498262274e-12
+    8.411287465847692e-11
+   -3.454792638808052e-13
+    -8.03530099351522e-13
+     -2.0515976960711e-11
+    8.247005922991752e-11
+ 1.25e+10    
+    8.260106791742072e-11
+   -2.051203263358619e-11
+    8.408342252782215e-11
+   -8.091108085305699e-13
+    -9.75185193508223e-12
+    8.410823417790929e-11
+    -3.49036424504476e-13
+   -8.059140898605311e-13
+   -2.051556712149199e-11
+    8.246475751057526e-11
+ 1.26e+10    
+    8.259578304406516e-11
+   -2.051165897564893e-11
+    8.407885518191198e-11
+   -8.115291231964283e-13
+   -9.752280951913489e-12
+    8.410365383932732e-11
+   -3.526207016607644e-13
+   -8.083251552726716e-13
+   -2.051518931472565e-11
+    8.245949588812721e-11
+ 1.27e+10    
+    8.259053820170013e-11
+   -2.051131658165653e-11
+    8.407434754544791e-11
+   -8.139741673213037e-13
+   -9.752725423436705e-12
+     8.40991330897226e-11
+   -3.562313604611825e-13
+   -8.107628919989104e-13
+   -2.051484270189688e-11
+    8.245427407652187e-11
+ 1.28e+10    
+    8.258533312572158e-11
+   -2.051100463669429e-11
+    8.406989905683934e-11
+   -8.164455409514292e-13
+   -9.753184262385222e-12
+    8.409467137823762e-11
+   -3.598676739312578e-13
+   -8.132269000613702e-13
+   -2.051452646671711e-11
+    8.244909179319716e-11
+ 1.29e+10    
+     8.25801675533551e-11
+   -2.051072234772721e-11
+    8.406550915638812e-11
+   -8.189428474570274e-13
+   -9.753656419804626e-12
+    8.409026815617734e-11
+   -3.635289228475696e-13
+   -8.157167828563568e-13
+   -2.051423981502394e-11
+     8.24439487584805e-11
+ 1.3e+10     
+    8.257504122311152e-11
+   -2.051046894348608e-11
+    8.406117728637681e-11
+   -8.214656933188992e-13
+   -9.754140885227554e-12
+    8.408592287705061e-11
+   -3.672143955945032e-13
+   -8.182321469409991e-13
+   -2.051398197465904e-11
+    8.243884469503976e-11
+ 1.31e+10    
+    8.256995387429211e-11
+   -2.051024367433414e-11
+    8.405690289118012e-11
+   -8.240136879366418e-13
+   -9.754636686769306e-12
+    8.408163499663627e-11
+    -3.70923388038741e-13
+   -8.207726018410119e-13
+   -2.051375219532558e-11
+    8.243377932738226e-11
+ 1.32e+10    
+    8.256490524654398e-11
+   -2.051004581211524e-11
+    8.405268541739701e-11
+   -8.265864434571271e-13
+   -9.755142891148821e-12
+    8.407740397307186e-11
+   -3.746552034194682e-13
+   -8.233377598786204e-13
+    -2.05135497484273e-11
+    8.242875238139868e-11
+ 1.33e+10    
+    8.255989507945757e-11
+   -2.050987464998443e-11
+    8.404852431399928e-11
+   -8.291835746215295e-13
+   -9.755658603640028e-12
+    8.407322926695949e-11
+   -3.784091522525611e-13
+    -8.25927236019237e-13
+    -2.05133739268895e-11
+    8.242376358394855e-11
+ 1.34e+10    
+    8.255492311220794e-11
+   -2.050972950222254e-11
+    8.404441903249258e-11
+   -8.318046986300438e-13
+   -9.756182967957332e-12
+    8.406911034148657e-11
+   -3.821845522470922e-13
+   -8.285406477354672e-13
+   -2.051322404496366e-11
+    8.241881266248523e-11
+ 1.35e+10    
+    8.254998908323385e-11
+   -2.050960970403502e-11
+    8.404036902708665e-11
+    -8.34449435023022e-13
+   -9.756715166079011e-12
+    8.406504666255859e-11
+   -3.859807282327111e-13
+   -8.311776148875923e-13
+   -2.051309943801695e-11
+    8.241389934471872e-11
+ 1.36e+10    
+    8.254509272995396e-11
+   -2.050951461133722e-11
+    8.403637375487373e-11
+   -8.371174055773905e-13
+   -9.757254418012511e-12
+    8.406103769893953e-11
+   -3.897970120965217e-13
+   -8.338377596191861e-13
+   -2.051299946230691e-11
+    8.240902335831124e-11
+ 1.37e+10    
+    8.254023378851626e-11
+   -2.050944360052577e-11
+    8.403243267601081e-11
+   -8.398082342173912e-13
+   -9.757799981504639e-12
+    8.405708292240027e-11
+   -3.936327427282176e-13
+    -8.36520706267192e-13
+   -2.051292349474333e-11
+    8.240418443060612e-11
+ 1.38e+10    
+    8.253541199357904e-11
+   -2.050939606823758e-11
+    8.402854525390252e-11
+    -8.42521546939029e-13
+   -9.758351151699603e-12
+    8.405318180786831e-11
+   -3.974872659723867e-13
+   -8.392260812852891e-13
+   -2.051287093263708e-11
+    8.239938228838595e-11
+ 1.39e+10    
+    8.253062707812078e-11
+   -2.050937143109734e-11
+    8.402471095538584e-11
+   -8.452569717468316e-13
+   -9.758907260748057e-12
+    8.404933383358154e-11
+   -4.013599345869502e-13
+   -8.419535131799685e-13
+   -2.051284119343777e-11
+    8.239461665765912e-11
+ 1.4e+10     
+    8.252587877327766e-11
+   -2.050936912545402e-11
+    8.402092925091097e-11
+   -8.480141386028139e-13
+   -9.759467677369957e-12
+    8.404553848124001e-11
+   -4.052501082067986e-13
+   -8.447026324583342e-13
+    -2.05128337144604e-11
+    8.238988726347156e-11
+ 1.41e+10    
+    8.252116680820505e-11
+   -2.050938860710731e-11
+    8.401719961471912e-11
+   -8.507926793861943e-13
+   -9.760031806373516e-12
+    8.404179523615659e-11
+   -4.091571533118672e-13
+   -8.474730715869946e-13
+   -2.051284795260209e-11
+    8.238519382974297e-11
+ 1.42e+10    
+    8.251649090996254e-11
+   -2.050942935102445e-11
+    8.401352152501382e-11
+   -8.535922278639625e-13
+   -9.760599088132969e-12
+     8.40381035874029e-11
+   -4.130804431987972e-13
+    -8.50264464961375e-13
+   -2.051288338404945e-11
+    8.238053607912491e-11
+ 1.43e+10    
+    8.251185080342002e-11
+   -2.050949085104867e-11
+    8.400989446412764e-11
+   -8.564124196707776e-13
+   -9.761168998027698e-12
+    8.403446302795216e-11
+    -4.17019357955584e-13
+   -8.530764488848136e-13
+   -2.051293950397746e-11
+    8.237591373287957e-11
+ 1.44e+10    
+    8.250724621118315e-11
+   -2.050957261959919e-11
+    8.400631791867802e-11
+   -8.592528922983658e-13
+    -9.76174104584483e-12
+    8.403087305481377e-11
+   -4.209732844386483e-13
+   -8.559086615566535e-13
+   -2.051301582624045e-11
+    8.237132651077781e-11
+ 1.45e+10    
+    8.250267685353662e-11
+   -2.050967418736395e-11
+     8.40027913797166e-11
+   -8.621132850933317e-13
+   -9.762314775147713e-12
+    8.402733316916195e-11
+   -4.249416162516385e-13
+   -8.587607430689951e-13
+    -2.05131118830558e-11
+    8.236677413101381e-11
+ 1.46e+10    
+    8.249814244840364e-11
+   -2.050979510298546e-11
+    8.399931434286763e-11
+   -8.649932392629049e-13
+   -9.762889762612633e-12
+    8.402384287645612e-11
+   -4.289237537256891e-13
+   -8.616323354113398e-13
+   -2.051322722468105e-11
+    8.236225631013684e-11
+ 1.47e+10    
+    8.249364271132073e-11
+    -2.05099349327406e-11
+    8.399588630845614e-11
+   -8.678923978882362e-13
+    -9.76346561733587e-12
+    8.402040168655182e-11
+   -4.329191039005232e-13
+   -8.645230824826745e-13
+   -2.051336141908496e-11
+    8.235777276299691e-11
+ 1.48e+10    
+    8.248917735542554e-11
+   -2.051009326021443e-11
+    8.399250678162578e-11
+   -8.708104059444703e-13
+   -9.764041980113529e-12
+    8.401700911380365e-11
+   -4.369270805061698e-13
+    -8.67432630110399e-13
+    -2.05135140516133e-11
+    8.235332320270431e-11
+ 1.49e+10    
+    8.248474609145679e-11
+   -2.051026968596893e-11
+    8.398917527244394e-11
+   -8.737469103271718e-13
+   -9.764618522695898e-12
+    8.401366467715672e-11
+   -4.409471039448992e-13
+   -8.703606260756423e-13
+   -2.051368472464961e-11
+    8.234890734060189e-11
+ 1.5e+10     
+    8.248034862776677e-11
+   -2.051046382720759e-11
+    8.398589129599691e-11
+    -8.76701559884786e-13
+    -9.76519494701916e-12
+    8.401036790022889e-11
+   -4.449786012730883e-13
+   -8.733067201443597e-13
+   -2.051387305727168e-11
+    8.234452488624776e-11
+ 1.51e+10    
+    8.247598467034185e-11
+   -2.051067531743544e-11
+    8.398265437247211e-11
+   -8.796740054562722e-13
+   -9.765770984416049e-12
+    8.400711831138271e-11
+   -4.490210061827764e-13
+   -8.762705641038978e-13
+   -2.051407868490434e-11
+     8.23401755474086e-11
+ 1.52e+10    
+    8.247165392283326e-11
+    -2.05109038061158e-11
+     8.39794640272288e-11
+   -8.826638999135878e-13
+   -9.766346394808015e-12
+    8.400391544378607e-11
+   -4.530737589827424e-13
+   -8.792518118043598e-13
+   -2.051430125896897e-11
+    8.233585903006311e-11
+ 1.53e+10    
+    8.246735608659612e-11
+   -2.051114895832407e-11
+    8.397631979085684e-11
+   -8.856708982087284e-13
+   -9.766920965880781e-12
+    8.400075883546289e-11
+   -4.571363065788698e-13
+   -8.822501192042973e-13
+   -2.051454044653022e-11
+    8.233157503841229e-11
+ 1.54e+10    
+     8.24630908607346e-11
+   -2.051141045439875e-11
+    8.397322119922389e-11
+    -8.88694657424617e-13
+   -9.767494512245605e-12
+    8.399764802933321e-11
+   -4.612081024536443e-13
+   -8.852651444205019e-13
+   -2.051479592994048e-11
+    8.232732327489854e-11
+ 1.55e+10    
+    8.245885794215461e-11
+   -2.051168798959068e-11
+    8.397016779351053e-11
+   -8.917348368294066e-13
+   -9.768066874588195e-12
+     8.39945825732421e-11
+   -4.652886066447128e-13
+    -8.88296547781126e-13
+   -2.051506740648248e-11
+    8.232310344023114e-11
+ 1.56e+10    
+    8.245465702562132e-11
+   -2.051198127371047e-11
+    8.396715912023504e-11
+   -8.947910979339943e-13
+   -9.768637918807566e-12
+     8.39915620199797e-11
+   -4.693772857223343e-13
+   -8.913439918819376e-13
+   -2.051535458801086e-11
+    8.231891523341799e-11
+ 1.57e+10    
+    8.245048780382204e-11
+   -2.051229003077494e-11
+    8.396419473126561e-11
+   -8.978631045518122e-13
+    -9.76920753514669e-12
+    8.398858592728992e-11
+   -4.734736127657481e-13
+   -8.944071416450828e-13
+   -2.051565720059256e-11
+    8.231475835180236e-11
+ 1.58e+10    
+     8.24463499674333e-11
+   -2.051261399865266e-11
+    8.396127418382353e-11
+   -9.009505228611879e-13
+   -9.769775637316956e-12
+    8.398565385786988e-11
+   -4.775770673382329e-13
+   -8.974856643801799e-13
+   -2.051597498414678e-11
+    8.231063249110526e-11
+ 1.59e+10    
+    8.244224320519138e-11
+   -2.051295292870946e-11
+    8.395839704047479e-11
+   -9.040530214691672e-13
+   -9.770342161618766e-12
+     8.39827653793609e-11
+   -4.816871354609793e-13
+   -9.005792298470421e-13
+   -2.051630769208525e-11
+    8.230653734547125e-11
+ 1.6e+10     
+    8.243816720396615e-11
+   -2.051330658545389e-11
+    8.395556286911218e-11
+   -9.071702714768012e-13
+   -9.770907066059585e-12
+    8.397992006432846e-11
+   -4.858033095856573e-13
+   -9.036875103198834e-13
+   -2.051665509095251e-11
+    8.230247260751849e-11
+ 1.61e+10    
+      8.2434121648838e-11
+   -2.051367474618331e-11
+    8.395277124292848e-11
+   -9.103019465454938e-13
+   -9.771470329471904e-12
+    8.397711749023566e-11
+   -4.899250885656676e-13
+   -9.068101806524155e-13
+   -2.051701696006721e-11
+    8.229843796839175e-11
+ 1.62e+10    
+    8.243010622317575e-11
+    -2.05140572006308e-11
+    8.395002174037974e-11
+   -9.134477229638923e-13
+   -9.772031950632603e-12
+     8.39743572394076e-11
+   -4.940519776260859e-13
+   -9.099469183437116e-13
+   -2.051739309116472e-11
+    8.229443311781893e-11
+ 1.63e+10    
+    8.242612060871763e-11
+   -2.051445375061345e-11
+    8.394731394514079e-11
+   -9.166072797149068e-13
+   -9.772591947385475e-12
+    8.397163889898746e-11
+   -4.981834883323534e-13
+    -9.13097403604229e-13
+   -2.051778328804081e-11
+     8.22904577441684e-11
+ 1.64e+10    
+    8.242216448565298e-11
+   -2.051486420968244e-11
+     8.39446474460532e-11
+   -9.197802985429625e-13
+   -9.773150355768892e-12
+    8.396896206088679e-11
+   -5.023191385575977e-13
+   -9.162613194218693e-13
+   -2.051818736619781e-11
+    8.228651153451069e-11
+ 1.65e+10    
+    8.241823753270483e-11
+   -2.051528840277478e-11
+    8.394202183706459e-11
+   -9.229664640205361e-13
+   -9.773707229149728e-12
+    8.396632632172782e-11
+   -5.064584524487777e-13
+   -9.194383516274688e-13
+   -2.051860515249265e-11
+    8.228259417467931e-11
+ 1.66e+10    
+    8.241433942721358e-11
+   -2.051572616586776e-11
+    8.393943671716211e-11
+   -9.261654636141568e-13
+   -9.774262637365587e-12
+    8.396373128278003e-11
+   -5.106009603915205e-13
+   -9.226281889599126e-13
+   -2.051903648478765e-11
+    8.227870534933517e-11
+ 1.67e+10    
+    8.241046984522073e-11
+   -2.051617734563579e-11
+    8.393689169029949e-11
+   -9.293769877493765e-13
+   -9.774816665876432e-12
+    8.396117654989133e-11
+   -5.147461989738208e-13
+   -9.258305231298719e-13
+   -2.051948121160415e-11
+    8.227484474203042e-11
+ 1.68e+10    
+    8.240662846155314e-11
+    -2.05166417991104e-11
+    8.393438636531775e-11
+   -9.326007298744054e-13
+   -9.775369414927207e-12
+    8.395866173341329e-11
+    -5.18893710948544e-13
+   -9.290450488825942e-13
+   -2.051993919177942e-11
+    8.227101203527445e-11
+ 1.69e+10    
+    8.240281494990677e-11
+   -2.051711939334332e-11
+    8.393192035586102e-11
+   -9.358363865222611e-13
+   -9.775920998722512e-12
+    8.395618644812173e-11
+   -5.230430451948192e-13
+   -9.322714640590487e-13
+   -2.052041029412678e-11
+    8.226720691059903e-11
+ 1.7e+10     
+    8.239902898293044e-11
+   -2.051761000507324e-11
+    8.392949328028786e-11
+   -9.390836573711873e-13
+   -9.776471544614861e-12
+    8.395375031313354e-11
+   -5.271937566783493e-13
+   -9.355094696554098e-13
+   -2.052089439709988e-11
+    8.226342904862529e-11
+ 1.71e+10    
+    8.239527023230905e-11
+   -2.051811352039623e-11
+    8.392710476157748e-11
+   -9.423422453030182e-13
+   -9.777021192307351e-12
+    8.395135295181976e-11
+   -5.313454064107297e-13
+   -9.387587698803892e-13
+   -2.052139138846067e-11
+    8.225967812912953e-11
+ 1.72e+10    
+    8.239153836884569e-11
+   -2.051862983444032e-11
+    8.392475442723314e-11
+   -9.456118564593566e-13
+    -9.77757009307182e-12
+    8.394899399171378e-11
+   -5.354975614077683e-13
+   -9.420190722106207e-13
+   -2.052190116495181e-11
+    8.225595383111054e-11
+ 1.73e+10    
+    8.238783306254408e-11
+   -2.051915885104427e-11
+    8.392244190918159e-11
+   -9.488922002954936e-13
+   -9.778118408983618e-12
+    8.394667306441918e-11
+   -5.396497946468749e-13
+   -9.452900874435806e-13
+   -2.052242363197344e-11
+    8.225225583285514e-11
+ 1.74e+10    
+    8.238415398268857e-11
+   -2.051970048244087e-11
+    8.392016684367028e-11
+    -9.52182989631625e-13
+   -9.778666312173591e-12
+     8.39443898055125e-11
+   -5.438016850235846e-13
+   -9.485715297480023e-13
+    -2.05229587032645e-11
+    8.224858381200432e-11
+ 1.75e+10    
+    8.238050079792422e-11
+   -2.052025464894478e-11
+     8.39179288711612e-11
+   -9.554839407014961e-13
+   -9.779213984098234e-12
+    8.394214385444671e-11
+   -5.479528173072793e-13
+   -9.518631167116237e-13
+   -2.052350630058958e-11
+    8.224493744561946e-11
+ 1.76e+10    
+    8.237687317633524e-11
+   -2.052082127864545e-11
+    8.391572763622438e-11
+   -9.587947731982184e-13
+   -9.779761614828534e-12
+    8.393993485445032e-11
+   -5.521027820961118e-13
+   -9.551645693861556e-13
+   -2.052406635342979e-11
+    8.224131641024609e-11
+ 1.77e+10    
+    8.237327078552254e-11
+   -2.052140030710506e-11
+    8.391356278742817e-11
+   -9.621152103171606e-13
+   -9.780309402358205e-12
+    8.393776245242703e-11
+   -5.562511757712027e-13
+   -9.584756123293945e-13
+   -2.052463879867977e-11
+    8.223772038197994e-11
+ 1.78e+10    
+    8.236969329267933e-11
+   -2.052199167706143e-11
+    8.391143397722937e-11
+   -9.654449787957549e-13
+   -9.780857551931833e-12
+     8.39356262988543e-11
+   -5.603976004502108e-13
+   -9.617959736441701e-13
+   -2.052522358034969e-11
+    8.223414903652921e-11
+ 1.79e+10    
+    8.236614036466556e-11
+    -2.05225953381365e-11
+    8.390934086186241e-11
+   -9.687838089502528e-13
+   -9.781406275393201e-12
+    8.393352604768095e-11
+   -5.645416639402338e-13
+   -9.651253850144023e-13
+   -2.052582064927276e-11
+    8.223060204927814e-11
+ 1.8e+10     
+    8.236261166808186e-11
+   -2.052321124655028e-11
+    8.390728310122819e-11
+   -9.721314347093594e-13
+    -9.78195579055442e-12
+    8.393146135622477e-11
+    -5.68682979690162e-13
+   -9.684635817378412e-13
+   -2.052642996281856e-11
+    8.222707909534927e-11
+ 1.81e+10    
+    8.235910686934052e-11
+   -2.052383936484025e-11
+    8.390526035878203e-11
+   -9.754875936445552e-13
+   -9.782506320585722e-12
+    8.392943188507026e-11
+   -5.728211667424678e-13
+   -9.718103027557846e-13
+   -2.052705148461187e-11
+    8.222357984966368e-11
+ 1.82e+10    
+    8.235562563473583e-11
+   -2.052447966158667e-11
+    8.390327230142335e-11
+   -9.788520269971318e-13
+   -9.783058093426708e-12
+    8.392743729796703e-11
+   -5.769558496845935e-13
+   -9.751652906792877e-13
+   -2.052768518425768e-11
+      8.2220103987002e-11
+ 1.83e+10    
+    8.235216763051265e-11
+   -2.052513211114332e-11
+    8.390131859938427e-11
+   -9.822244797021066e-13
+   -9.783611341218486e-12
+     8.39254772617286e-11
+   -5.810866585997936e-13
+   -9.785282918124315e-13
+   -2.052833103707193e-11
+    8.221665118206341e-11
+ 1.84e+10    
+    8.234873252293367e-11
+   -2.052579669337461e-11
+    8.389939892612018e-11
+   -9.856047004086879e-13
+   -9.784166299757462e-12
+    8.392355144613203e-11
+   -5.852132290176587e-13
+   -9.818990561720295e-13
+   -2.052898902381815e-11
+     8.22132211095232e-11
+ 1.85e+10    
+    8.234531997834435e-11
+    -2.05264733933981e-11
+    8.389751295820068e-11
+   -9.889924414975236e-13
+   -9.784723207970233e-12
+    8.392165952381926e-11
+   -5.893352018642263e-13
+   -9.852773375042729e-13
+   -2.052965913045062e-11
+    8.220981344409025e-11
+ 1.86e+10    
+     8.23419296632376e-11
+   -2.052716220133341e-11
+    8.389566037520162e-11
+    -9.92387459094692e-13
+   -9.785282307409842e-12
+    8.391980117019951e-11
+   -5.934522234118152e-13
+   -9.886628932979745e-13
+   -2.053034134786313e-11
+    8.220642786056289e-11
+ 1.87e+10    
+     8.23385612443152e-11
+   -2.052786311205692e-11
+    8.389384085959936e-11
+   -9.957895130823318e-13
+   -9.785843841773224e-12
+    8.391797606335322e-11
+   -5.975639452285597e-13
+    -9.92055484794628e-13
+   -2.053103567164425e-11
+    8.220306403388334e-11
+ 1.88e+10    
+    8.233521438854891e-11
+   -2.052857612496261e-11
+    8.389205409666614e-11
+   -9.991983671061973e-13
+    -9.78640805643968e-12
+    8.391618388393802e-11
+   -6.016700241276749e-13
+   -9.954548769952909e-13
+   -2.053174210183869e-11
+    8.219972163919204e-11
+ 1.89e+10    
+    8.233188876323961e-11
+   -2.052930124372886e-11
+    8.389029977436722e-11
+   -1.002613788579926e-12
+   -9.786975198030088e-12
+    8.391442431509607e-11
+   -6.057701221165255e-13
+   -9.988608386643003e-13
+   -2.053246064271485e-11
+    8.219640035187969e-11
+ 1.9e+10     
+    8.232858403607443e-11
+   -2.053003847609173e-11
+     8.38885775832604e-11
+   -1.006035548686278e-12
+   -9.787545513986788e-12
+    8.391269704236492e-11
+   -6.098639063455184e-13
+   -1.002273142329797e-12
+   -2.053319130253853e-11
+    8.219309984763839e-11
+ 1.91e+10    
+    8.232529987518317e-11
+   -2.053078783362377e-11
+    8.388688721639713e-11
+   -1.009463422375149e-12
+   -9.788119252173676e-12
+    8.391100175358829e-11
+   -6.139510490568258e-13
+    -1.00569156428129e-12
+   -2.053393409335293e-11
+     8.21898198025124e-11
+ 1.92e+10    
+    8.232203594919199e-11
+   -2.053154933151925e-11
+    8.388522836922669e-11
+   -1.012897188358807e-12
+   -9.788696660496398e-12
+    8.390933813883168e-11
+   -6.180312275329833e-13
+   -1.009115884564209e-12
+   -2.053468903076493e-11
+     8.21865598929472e-11
+ 1.93e+10    
+     8.23187919272772e-11
+   -2.053232298838555e-11
+    8.388360073950189e-11
+   -1.016336629104018e-12
+   -9.789277986541905e-12
+    8.390770589029872e-11
+   -6.221041240453893e-13
+    -1.01254588697156e-12
+   -2.053545613373722e-11
+    8.218331979583691e-11
+ 1.94e+10    
+    8.231556747921539e-11
+   -2.053310882604021e-11
+    8.388200402718778e-11
+    -1.01978153082134e-12
+   -9.789863477237556e-12
+    8.390610470225049e-11
+   -6.261694258027508e-13
+    -1.01598135903265e-12
+   -2.053623542438694e-11
+    8.218009918857141e-11
+ 1.95e+10    
+    8.231236227543401e-11
+   -2.053390686931433e-11
+    8.388043793437271e-11
+   -1.023231683451808e-12
+   -9.790453378528783e-12
+    8.390453427092796e-11
+    -6.30226824899442e-13
+   -1.019422091999211e-12
+    -2.05370269277902e-11
+    8.217689774908195e-11
+ 1.96e+10    
+    8.230917598705944e-11
+   -2.053471714586188e-11
+    8.387890216518249e-11
+   -1.026686880650702e-12
+    -9.79104793507529e-12
+    8.390299429447659e-11
+   -6.342760182638729e-13
+    -1.02286788082872e-12
+   -2.053783067179275e-11
+    8.217371515588563e-11
+ 1.97e+10    
+    8.230600828596376e-11
+   -2.053553968597479e-11
+    8.387739642569624e-11
+   -1.030146919768954e-12
+   -9.791647389965139e-12
+    8.390148447287378e-11
+   -6.383167076068293e-13
+     -1.0263185241652e-12
+   -2.053864668682655e-11
+    8.217055108812856e-11
+ 1.98e+10    
+    8.230285884481026e-11
+   -2.053637452240398e-11
+    8.387592042386637e-11
+   -1.033611601831843e-12
+   -9.792251984446344e-12
+    8.390000450785919e-11
+   -6.423485993698378e-13
+   -1.029773824317563e-12
+   -2.053947500573254e-11
+     8.21674052256285e-11
+ 1.99e+10    
+    8.229972733709704e-11
+   -2.053722169018622e-11
+    8.387447386944006e-11
+   -1.037080731515473e-12
+   -9.792861957675346e-12
+    8.389855410286739e-11
+   -6.463714046735668e-13
+   -1.033233587235517e-12
+   -2.054031566358881e-11
+    8.216427724891561e-11
+ 2e+10       
+    8.229661343720017e-11
+   -2.053808122647679e-11
+    8.387305647388478e-11
+   -1.040554117120871e-12
+   -9.793477546482158e-12
+    8.389713296296473e-11
+   -6.503848392662639e-13
+    -1.03669762248321e-12
+   -2.054116869754532e-11
+     8.21611668392729e-11
+ 2.01e+10    
+    8.229351682041439e-11
+   -2.053895317038765e-11
+    8.387166795031538e-11
+   -1.044031570545842e-12
+   -9.794098985151281e-12
+    8.389574079478703e-11
+   -6.543886234722899e-13
+   -1.040165743210641e-12
+   -2.054203414666343e-11
+    8.215807367877469e-11
+ 2.02e+10    
+    8.229043716299326e-11
+   -2.053983756283139e-11
+    8.387030801342553e-11
+   -1.047512907254796e-12
+   -9.794726505218328e-12
+    8.389437730648203e-11
+   -6.583824821407167e-13
+   -1.043637766123112e-12
+   -2.054291205176209e-11
+    8.215499745032538e-11
+ 2.03e+10    
+    8.228737414218736e-11
+   -2.054073444637045e-11
+    8.386897637942092e-11
+   -1.050997946246547e-12
+   -9.795360335281395e-12
+    8.389304220765338e-11
+    -6.62366144594023e-13
+    -1.04711351144848e-12
+   -2.054380245526864e-11
+    8.215193783769506e-11
+ 2.04e+10    
+    8.228432743628228e-11
+   -2.054164386507219e-11
+    8.386767276595586e-11
+   -1.054486510020266e-12
+   -9.796000700827038e-12
+     8.38917352093083e-11
+   -6.663393445769256e-13
+   -1.050592802902778e-12
+   -2.054470540107595e-11
+    8.214889452555661e-11
+ 2.05e+10    
+    8.228129672463343e-11
+   -2.054256586436882e-11
+    8.386639689207253e-11
+   -1.057978424539541e-12
+   -9.796647824069983e-12
+    8.389045602380739e-11
+   -6.703018202053082e-13
+    -1.05407546765385e-12
+   -2.054562093440426e-11
+    8.214586719951967e-11
+ 2.06e+10    
+    8.227828168770209e-11
+   -2.054350049092289e-11
+    8.386514847814362e-11
+   -1.061473519194785e-12
+   -9.797301923806501e-12
+    8.388920436481813e-11
+   -6.742533139153468e-13
+   -1.057561336283391e-12
+   -2.054654910166876e-11
+    8.214285554616481e-11
+ 2.07e+10    
+    8.227528200708798e-11
+   -2.054444779249792e-11
+    8.386392724581719e-11
+   -1.064971626764173e-12
+    -9.79796321528038e-12
+    8.388797994727014e-11
+   -6.781935724127003e-13
+   -1.061050242747462e-12
+   -2.054748995035215e-11
+    8.213985925307611e-11
+ 2.08e+10    
+    8.227229736556212e-11
+   -2.054540781783401e-11
+    8.386273291796506e-11
+   -1.068472583372904e-12
+   -9.798631910061503e-12
+    8.388678248731425e-11
+   -6.821223466219633e-13
+   -1.064542024335371e-12
+   -2.054844352888251e-11
+    8.213687800887321e-11
+ 2.09e+10    
+     8.22693274470977e-11
+   -2.054638061652842e-11
+    8.386156521863334e-11
+   -1.071976228451183e-12
+   -9.799308215936123e-12
+    8.388561170228338e-11
+   -6.860393916362206e-13
+   -1.068036521627397e-12
+   -2.054940988651585e-11
+     8.21339115032421e-11
+ 2.1e+10     
+    8.226637193690055e-11
+   -2.054736623892118e-11
+    8.386042387299638e-11
+   -1.075482404690934e-12
+   -9.799992336808568e-12
+    8.388446731065695e-11
+   -6.899444666668232e-13
+    -1.07153357845099e-12
+   -2.055038907322389e-11
+    8.213095942696496e-11
+ 2.11e+10    
+    8.226343052143745e-11
+   -2.054836473598516e-11
+    8.385930860731338e-11
+   -1.078990958001185e-12
+   -9.800684472613848e-12
+    8.388334903202699e-11
+   -6.938373349933462e-13
+   -1.075033041836034e-12
+    -2.05513811395863e-11
+    8.212802147194921e-11
+ 2.12e+10    
+     8.22605028884649e-11
+   -2.054937615922121e-11
+    8.385821914888739e-11
+   -1.082501737462526e-12
+   -9.801384819240513e-12
+    8.388225658706782e-11
+   -6.977177639137863e-13
+   -1.078534761968785e-12
+    -2.05523861366879e-11
+    8.212509733125554e-11
+ 2.13e+10    
+    8.225758872705484e-11
+   -2.055040056055751e-11
+    8.385715522602743e-11
+   -1.086014595280417e-12
+   -9.802093568463593e-12
+    8.388118969750791e-11
+   -7.015855246948916e-13
+   -1.082038592144977e-12
+   -2.055340411602034e-11
+    8.212218669912511e-11
+ 2.14e+10    
+    8.225468772762133e-11
+   -2.055143799225342e-11
+    8.385611656801291e-11
+   -1.089529386737654e-12
+   -9.802810907886712e-12
+     8.38801480861038e-11
+   -7.054403925228253e-13
+   -1.085544388721995e-12
+   -2.055443512938808e-11
+    8.211928927100601e-11
+ 2.15e+10    
+    8.225179958194475e-11
+   -2.055248850680801e-11
+    8.385510290506142e-11
+   -1.093045970145984e-12
+   -9.803537020893494e-12
+     8.38791314766172e-11
+   -7.092821464539646e-13
+   -1.089052011070096e-12
+   -2.055547922881893e-11
+    8.211640474357841e-11
+ 2.16e+10    
+    8.224892398319588e-11
+   -2.055355215687246e-11
+    8.385411396829835e-11
+   -1.096564206796904e-12
+   -9.804272086607196e-12
+    8.387813959379405e-11
+   -7.131105693659962e-13
+    -1.09256132152311e-12
+    -2.05565364664787e-11
+    8.211353281477899e-11
+ 2.17e+10    
+    8.224606062595832e-11
+   -2.055462899516665e-11
+    8.385314948972905e-11
+   -1.100083960911958e-12
+   -9.805016279858627e-12
+    8.387717216334605e-11
+    -7.16925447909224e-13
+   -1.096072185328297e-12
+   -2.055760689459007e-11
+    8.211067318382539e-11
+ 2.18e+10    
+    8.224320920625082e-11
+   -2.055571907440005e-11
+    8.385220920221414e-11
+   -1.103605099592259e-12
+   -9.805769771161668e-12
+    8.387622891193468e-11
+   -7.207265724581555e-13
+   -1.099584470595727e-12
+   -2.055869056535541e-11
+    8.210782555123818e-11
+ 2.19e+10    
+    8.224036942154772e-11
+   -2.055682244719615e-11
+    8.385129283944691e-11
+   -1.107127492767639e-12
+   -9.806532726695984e-12
+    8.387530956715689e-11
+   -7.245137370633351e-13
+   -1.103098048247155e-12
+   -2.055978753088346e-11
+    8.210498961886369e-11
+ 2.2e+10     
+    8.223754097079935e-11
+     -2.0557939166021e-11
+    8.385040013593251e-11
+   -1.110651013145295e-12
+   -9.807305308296668e-12
+    8.387441385753343e-11
+   -7.282867394034425e-13
+   -1.106612791964459e-12
+   -2.056089784311993e-11
+    8.210216508989471e-11
+ 2.21e+10    
+     8.22347235544508e-11
+   -2.055906928311541e-11
+    8.384953082697109e-11
+   -1.114175536158105e-12
+   -9.808087673450397e-12
+    8.387354151249928e-11
+   -7.320453807376746e-13
+   -1.110128578137717e-12
+   -2.056202155378165e-11
+    8.209935166889142e-11
+ 2.22e+10    
+    8.223191687446072e-11
+   -2.056021285043063e-11
+    8.384868464864172e-11
+   -1.117700939912622e-12
+   -9.808879975297575e-12
+    8.387269226239598e-11
+   -7.357894658583979e-13
+    -1.11364528581303e-12
+   -2.056315871429448e-11
+     8.20965490618009e-11
+ 2.23e+10    
+      8.2229120634318e-11
+   -2.056136991956758e-11
+    8.384786133778875e-11
+   -1.121227105136895e-12
+   -9.809682362640202e-12
+    8.387186583846564e-11
+   -7.395188030440933e-13
+   -1.117162796640138e-12
+   -2.056430937573439e-11
+    8.209375697597622e-11
+ 2.24e+10    
+     8.22263345390591e-11
+    -2.05625405417196e-11
+    8.384706063201113e-11
+   -1.124753915128072e-12
+   -9.810494979955218e-12
+    8.387106197284769e-11
+   -7.432332040125745e-13
+   -1.120680994819859e-12
+   -2.056547358877226e-11
+    8.209097512019439e-11
+ 2.25e+10    
+    8.222355829528378e-11
+   -2.056372476761848e-11
+    8.384628226965342e-11
+   -1.128281255699898e-12
+   -9.811317967412827e-12
+     8.38702803985763e-11
+   -7.469324838745438e-13
+   -1.124199767051419e-12
+   -2.056665140362155e-11
+    8.208820320467431e-11
+ 2.26e+10    
+    8.222079161116944e-11
+   -2.056492264748331e-11
+    8.384552598979894e-11
+   -1.131809015130257e-12
+   -9.812151460899608e-12
+    8.386952084958102e-11
+    -7.50616461087389e-13
+    -1.12771900247985e-12
+    -2.05678428699896e-11
+    8.208544094109322e-11
+ 2.27e+10    
+    8.221803419648637e-11
+   -2.056613423097309e-11
+    8.384479153226454e-11
+   -1.135337084108599e-12
+   -9.812995592045859e-12
+    8.386878306068751e-11
+   -7.542849574093406e-13
+     -1.1312385926433e-12
+   -2.056904803703139e-11
+    8.208268804260289e-11
+ 2.28e+10    
+    8.221528576261057e-11
+   -2.056735956714175e-11
+    8.384407863759811e-11
+   -1.138865355683499e-12
+   -9.813850488257313e-12
+    8.386806676762113e-11
+    -7.57937797853926e-13
+   -1.134758431420445e-12
+   -2.057026695330671e-11
+     8.20799442238448e-11
+ 2.29e+10    
+    8.221254602253698e-11
+    -2.05685987043964e-11
+    8.384338704707745e-11
+   -1.142393725210355e-12
+   -9.814716272750465e-12
+    8.386737170701247e-11
+   -7.615748106447292e-13
+   -1.138278414978116e-12
+   -2.057149966674008e-11
+    8.207720920096542e-11
+ 2.3e+10     
+    8.220981469089118e-11
+   -2.056985169045815e-11
+    8.384271650271105e-11
+   -1.145922090299158e-12
+   -9.815593064591494e-12
+    8.386669761640198e-11
+   -7.651958271704814e-13
+   -1.141798441718961e-12
+   -2.057274622458306e-11
+    8.207448269162937e-11
+ 2.31e+10    
+    8.220709148394118e-11
+   -2.057111857232586e-11
+    8.384206674724068e-11
+   -1.149450350762615e-12
+   -9.816480978738511e-12
+    8.386604423424914e-11
+   -7.688006819404607e-13
+   -1.145318412229475e-12
+   -2.057400667337974e-11
+    8.207176441503351e-11
+ 2.32e+10    
+    8.220437611960779e-11
+   -2.057239939624236e-11
+    8.384143752414641e-11
+   -1.152978408564314e-12
+   -9.817380126086875e-12
+    8.386541129994126e-11
+   -7.723892125402677e-13
+   -1.148838229228158e-12
+   -2.057528105893446e-11
+    8.206905409191939e-11
+ 2.33e+10    
+    8.220166831747508e-11
+   -2.057369420766324e-11
+    8.384082857765175e-11
+   -1.156506167767393e-12
+   -9.818290613517106e-12
+    8.386479855380358e-11
+   -7.759612595878771e-13
+   -1.152357797514078e-12
+   -2.057656942628195e-11
+     8.20663514445855e-11
+ 2.34e+10    
+     8.21989677987994e-11
+   -2.057500305122807e-11
+    8.384023965273209e-11
+    -1.16003353448338e-12
+   -9.819212543945577e-12
+    8.386420573711109e-11
+    -7.79516666690077e-13
+   -1.155877023915702e-12
+   -2.057787181965997e-11
+    8.206365619689838e-11
+ 2.35e+10    
+    8.219627428651859e-11
+   -2.057632597073386e-11
+    8.383967049512348e-11
+   -1.163560416821491e-12
+   -9.820146016377372e-12
+    8.386363259210192e-11
+   -7.830552803992109e-13
+   -1.159395817240207e-12
+   -2.057918828248423e-11
+    8.206096807430401e-11
+ 2.36e+10    
+    8.219358750525968e-11
+   -2.057766300911103e-11
+    8.383912085133367e-11
+   -1.167086724838227e-12
+   -9.821091125961443e-12
+    8.386307886199043e-11
+   -7.865769501703098e-13
+   -1.162914088223033e-12
+   -2.058051885732526e-11
+    8.205828680383776e-11
+ 2.37e+10    
+    8.219090718134702e-11
+   -2.057901420840112e-11
+    8.383859046865421e-11
+   -1.170612370487517e-12
+   -9.822047964047471e-12
+    8.386254429098317e-11
+    -7.90081528318528e-13
+   -1.166431749478042e-12
+   -2.058186358588772e-11
+    8.205561211413419e-11
+ 2.38e+10    
+    8.218823304280855e-11
+   -2.058037960973709e-11
+    8.383807909517397e-11
+   -1.174137267571171e-12
+   -9.823016618244726e-12
+    8.386202862429438e-11
+   -7.935688699769735e-13
+   -1.169948715448084e-12
+   -2.058322250899139e-11
+    8.205294373543596e-11
+ 2.39e+10    
+    8.218556481938316e-11
+   -2.058175925332526e-11
+    8.383758647979379e-11
+   -1.177661331690012e-12
+   -9.823997172482158e-12
+    8.386153160816277e-11
+   -7.970388330548554e-13
+   -1.173464902356026e-12
+   -2.058459566655424e-11
+    8.205028139960285e-11
+ 2.4e+10     
+    8.218290224252589e-11
+   -2.058315317842921e-11
+    8.383711237224322e-11
+   -1.181184480195288e-12
+    -9.82498970707026e-12
+    8.386105298987004e-11
+   -8.004912781960389e-13
+   -1.176980228156358e-12
+   -2.058598309757744e-11
+    8.204762484011928e-11
+ 2.41e+10    
+     8.21802450454135e-11
+   -2.058456142335566e-11
+    8.383665652309693e-11
+   -1.184706632140777e-12
+   -9.825994298763783e-12
+    8.386059251775878e-11
+   -8.039260687379257e-13
+   -1.180494612487301e-12
+   -2.058738484013178e-11
+    8.204497379210182e-11
+ 2.42e+10    
+    8.217759296294917e-11
+   -2.058598402544215e-11
+    8.383621868379411e-11
+   -1.188227708235391e-12
+   -9.827011020825832e-12
+    8.386014994125236e-11
+    -8.07343070670709e-13
+   -1.184007976623518e-12
+   -2.058880093134623e-11
+    8.204232799230653e-11
+ 2.43e+10    
+    8.217494573176686e-11
+   -2.058742102104596e-11
+    8.383579860665695e-11
+   -1.191747630796327e-12
+   -9.828039943092558e-12
+    8.385972501087446e-11
+   -8.107421525970127e-13
+   -1.187520243429406e-12
+   -2.059023140739775e-11
+    8.203968717913483e-11
+ 2.44e+10    
+    8.217230309023531e-11
+   -2.058887244553534e-11
+    8.383539604491194e-11
+   -1.195266323702895e-12
+   -9.829081132038936e-12
+    8.385931747827009e-11
+   -8.141231856918861e-13
+   -1.191031337312951e-12
+   -2.059167630350271e-11
+    8.203705109263987e-11
+ 2.45e+10    
+    8.216966477846108e-11
+   -2.059033833328176e-11
+    8.383501075271084e-11
+   -1.198783712350782e-12
+   -9.830134650845062e-12
+    8.385892709622636e-11
+   -8.174860436631808e-13
+   -1.194541184180252e-12
+   -2.059313565390985e-11
+    8.203441947453129e-11
+ 2.46e+10    
+    8.216703053829113e-11
+   -2.059181871765362e-11
+    8.383464248515296e-11
+   -1.202299723607139e-12
+   -9.831200559462904e-12
+    8.385855361869453e-11
+   -8.208306027123081e-13
+   -1.198049711390666e-12
+   -2.059460949189464e-11
+    8.203179206818065e-11
+ 2.47e+10    
+    8.216440011331596e-11
+   -2.059331363101183e-11
+    8.383429099830849e-11
+   -1.205814285766152e-12
+   -9.832278914683582e-12
+    8.385819680081163e-11
+   -8.241567414953707e-13
+   -1.201556847712577e-12
+   -2.059609784975482e-11
+    8.202916861862602e-11
+ 2.48e+10    
+    8.216177324887077e-11
+   -2.059482310470624e-11
+    8.383395604924199e-11
+    -1.20932732850533e-12
+   -9.833369770204919e-12
+     8.38578563989234e-11
+    -8.27464341084661e-13
+   -1.205062523279876e-12
+   -2.059760075880728e-11
+    8.202654887257498e-11
+ 2.49e+10    
+    8.215914969203744e-11
+   -2.059634716907359e-11
+    8.383363739603745e-11
+   -1.212838782842432e-12
+   -9.834473176699171e-12
+     8.38575321706065e-11
+   -8.307532849305843e-13
+   -1.208566669549042e-12
+   -2.059911824938615e-11
+    8.202393257840911e-11
+ 2.5e+10     
+    8.215652919164499e-11
+   -2.059788585343637e-11
+    8.383333479782251e-11
+   -1.216348581093019e-12
+   -9.835589181880775e-12
+    8.385722387469179e-11
+   -8.340234588239338e-13
+    -1.21206921925696e-12
+   -2.060065035084184e-11
+    8.202131948618648e-11
+ 2.51e+10    
+    8.215391149827084e-11
+   -2.059943918610337e-11
+    8.383304801479514e-11
+    -1.21985665682876e-12
+   -9.836717830574321e-12
+    8.385693127128756e-11
+   -8.372747508585445e-13
+   -1.215570106379414e-12
+   -2.060219709154149e-11
+    8.201870934764424e-11
+ 2.52e+10    
+    8.215129636424067e-11
+   -2.060100719437069e-11
+    8.383277680824895e-11
+   -1.223362944836371e-12
+   -9.837859164782241e-12
+    8.385665412180263e-11
+   -8.405070513943815e-13
+   -1.219069266090211e-12
+   -2.060375849886999e-11
+    8.201610191620096e-11
+ 2.53e+10    
+    8.214868354362807e-11
+   -2.060258990452415e-11
+    8.383252094060031e-11
+   -1.226867381077223e-12
+    -9.83901322375233e-12
+    8.385639218896973e-11
+   -8.437202530209663e-13
+   -1.222566634721183e-12
+   -2.060533459923226e-11
+    8.201349694695824e-11
+ 2.54e+10    
+    8.214607279225431e-11
+   -2.060418734184265e-11
+    8.383228017541497e-11
+   -1.230369902647639e-12
+   -9.840180044045276e-12
+    8.385614523686904e-11
+   -8.469142505212384e-13
+   -1.226062149722608e-12
+   -2.060692541805621e-11
+    8.201089419670194e-11
+ 2.55e+10    
+    8.214346386768717e-11
+   -2.060579953060212e-11
+    8.383205427743539e-11
+   -1.233870447739984e-12
+   -9.841359659601607e-12
+    8.385591303095167e-11
+   -8.500889408357828e-13
+   -1.229555749624583e-12
+   -2.060853097979685e-11
+    8.200829342390314e-11
+ 2.56e+10    
+    8.214085652923978e-11
+   -2.060742649408083e-11
+    8.383184301260858e-11
+   -1.237368955604287e-12
+   -9.842552101808364e-12
+    8.385569533806256e-11
+   -8.532442230274623e-13
+   -1.233047373999073e-12
+   -2.061015130794061e-11
+    8.200569438871893e-11
+ 2.57e+10    
+    8.213825053796862e-11
+   -2.060906825456499e-11
+    8.383164614811287e-11
+    -1.24086536651071e-12
+   -9.843757399565429e-12
+    8.385549192646405e-11
+   -8.563799982464533e-13
+   -1.236536963422482e-12
+   -2.061178642501103e-11
+    8.200309685299166e-11
+ 2.58e+10    
+    8.213564565667162e-11
+   -2.061072483335531e-11
+    8.383146345238634e-11
+   -1.244359621712644e-12
+   -9.844975579351208e-12
+    8.385530256585878e-11
+   -8.594961696956548e-13
+   -1.240024459439176e-12
+   -2.061343635257465e-11
+     8.20005005802499e-11
+ 2.59e+10    
+    8.213304164988624e-11
+   -2.061239625077452e-11
+    8.383129469515461e-11
+   -1.247851663410499e-12
+   -9.846206665287866e-12
+    8.385512702741233e-11
+   -8.625926425965286e-13
+   -1.243509804525604e-12
+   -2.061510111124779e-11
+    8.199790533570661e-11
+ 2.6e+10     
+    8.213043828388562e-11
+    -2.06140825261749e-11
+     8.38311396474582e-11
+   -1.251341434716239e-12
+   -9.847450679205974e-12
+    8.385496508377559e-11
+   -8.656693241552946e-13
+   -1.246992942055107e-12
+   -2.061678072070372e-11
+    8.199531088625879e-11
+ 2.61e+10    
+    8.212783532667681e-11
+   -2.061578367794711e-11
+     8.38309980816807e-11
+    -1.25482887961859e-12
+   -9.848707640708468e-12
+    8.385481650910748e-11
+   -8.687261235295787e-13
+   -1.250473816263479e-12
+   -2.061847519968067e-11
+    8.199271700048608e-11
+ 2.62e+10    
+    8.212523254799668e-11
+   -2.061749972352909e-11
+    8.383086977157601e-11
+   -1.258313942948948e-12
+   -9.849977567233893e-12
+    8.385468107909596e-11
+   -8.717629517954087e-13
+   -1.253952372215232e-12
+   -2.062018456598988e-11
+    8.199012344864879e-11
+ 2.63e+10    
+    8.212262971930848e-11
+   -2.061923067941565e-11
+    8.383075449229568e-11
+   -1.261796570347988e-12
+   -9.851260474119053e-12
+    8.385455857098028e-11
+   -8.747797219146362e-13
+   -1.257428555770547e-12
+   -2.062190883652464e-11
+    8.198753000268595e-11
+ 2.64e+10    
+    8.212002661379771e-11
+   -2.062097656116852e-11
+    8.383065202041678e-11
+   -1.265276708232917e-12
+   -9.852556374660817e-12
+    8.385444876357112e-11
+   -8.777763487027616e-13
+   -1.260902313552973e-12
+   -2.062364802726923e-11
+    8.198493643621307e-11
+ 2.65e+10    
+    8.211742300636799e-11
+   -2.062273738342674e-11
+    8.383056213396762e-11
+   -1.268754303765544e-12
+    -9.85386528017705e-12
+    8.385435143727166e-11
+   -8.807527487971404e-13
+   -1.264373592917724e-12
+   -2.062540215330856e-11
+    8.198234252451911e-11
+ 2.66e+10    
+    8.211481867363675e-11
+   -2.062451315991769e-11
+    8.383048461245524e-11
+   -1.272229304820863e-12
+    -9.85518720006692e-12
+    8.385426637409703e-11
+    -8.83708840625611e-13
+   -1.267842341920779e-12
+   -2.062717122883819e-11
+    8.197974804456398e-11
+ 2.67e+10    
+    8.211221339392988e-11
+   -2.062630390346802e-11
+    8.383041923689074e-11
+   -1.275701659956469e-12
+   -9.856522141870207e-12
+    8.385419335769409e-11
+   -8.866445443754932e-13
+   -1.271308509288608e-12
+    -2.06289552671743e-11
+    8.197715277497458e-11
+ 2.68e+10    
+    8.210960694727737e-11
+   -2.062810962601539e-11
+    8.383036578981564e-11
+   -1.279171318382584e-12
+   -9.857870111325783e-12
+    8.385413217336004e-11
+   -8.895597819630277e-13
+   -1.274772044388553e-12
+   -2.063075428076437e-11
+    8.197455649604162e-11
+ 2.69e+10    
+     8.21069991154072e-11
+   -2.062993033862006e-11
+    8.383032405532651e-11
+   -1.282638229932674e-12
+   -9.859231112429204e-12
+    8.385408260806028e-11
+   -8.924544770031652e-13
+   -1.278232897200015e-12
+   -2.063256828119765e-11
+    8.197195898971546e-11
+ 2.7e+10     
+    8.210438968174038e-11
+   -2.063176605147696e-11
+     8.38302938190994e-11
+   -1.286102345034933e-12
+   -9.860605147489362e-12
+    8.385404445044654e-11
+   -8.953285547797984e-13
+   -1.281691018286101e-12
+   -2.063439727921635e-11
+    8.196936003960204e-11
+ 2.71e+10    
+    8.210177843138474e-11
+     -2.0633616773928e-11
+     8.38302748684144e-11
+   -1.289563614684192e-12
+   -9.861992217184241e-12
+    8.385401749087264e-11
+   -8.981819422163732e-13
+   -1.285146358766137e-12
+   -2.063624128472647e-11
+    8.196675943095845e-11
+ 2.72e+10    
+    8.209916515112922e-11
+   -2.063548251447427e-11
+     8.38302669921783e-11
+   -1.293021990414691e-12
+   -9.863392320615689e-12
+     8.38540015214118e-11
+   -9.010145678468734e-13
+   -1.288598870288719e-12
+   -2.063810030680925e-11
+     8.19641569506879e-11
+ 2.73e+10    
+    8.209654962943714e-11
+   -2.063736328078871e-11
+    8.383026998094777e-11
+   -1.296477424273364e-12
+   -9.864805455363204e-12
+    8.385399633587065e-11
+    -9.03826361787252e-13
+   -1.292048505005442e-12
+   -2.063997435373229e-11
+    8.196155238733495e-11
+ 2.74e+10    
+    8.209393165643997e-11
+   -2.063925907972871e-11
+    8.383028362695074e-11
+   -1.299929868793745e-12
+   -9.866231617536869e-12
+    8.385400172980458e-11
+   -9.066172557072229e-13
+   -1.295495215545291e-12
+   -2.064186343296117e-11
+    8.195894553108033e-11
+ 2.75e+10    
+    8.209131102393055e-11
+   -2.064116991734877e-11
+    8.383030772410781e-11
+   -1.303379276970656e-12
+   -9.867670801829145e-12
+    8.385401750053154e-11
+   -9.093871828024485e-13
+    -1.29893895498961e-12
+   -2.064376755117099e-11
+    8.195633617373493e-11
+ 2.76e+10    
+    8.208868752535627e-11
+   -2.064309579891352e-11
+    8.383034206805245e-11
+   -1.306825602235382e-12
+   -9.869123001565743e-12
+    8.385404344714428e-11
+   -9.121360777671297e-13
+   -1.302379676847774e-12
+   -2.064568671425778e-11
+    8.195372410873459e-11
+ 2.77e+10    
+    8.208606095581144e-11
+   -2.064503672891016e-11
+    8.383038645615056e-11
+   -1.310268798431487e-12
+   -9.870588208755561e-12
+    8.385407937052304e-11
+    -9.14863876766998e-13
+   -1.305817335033414e-12
+   -2.064762092735025e-11
+    8.195110913113399e-11
+ 2.78e+10    
+    8.208343111203045e-11
+   -2.064699271106155e-11
+    8.383044068751869e-11
+   -1.313708819791304e-12
+   -9.872066414139455e-12
+    8.385412507334636e-11
+   -9.175705174126731e-13
+   -1.309251883841284e-12
+   -2.064957019482129e-11
+    8.194849103760027e-11
+ 2.79e+10    
+       8.208079779238e-11
+     -2.0648963748339e-11
+    8.383050456304198e-11
+    -1.31714562091298e-12
+   -9.873557607238107e-12
+    8.385418036010166e-11
+   -9.202559387334223e-13
+   -1.312683277924713e-12
+    -2.06515345202995e-11
+    8.194586962640643e-11
+ 2.8e+10     
+    8.207816079685149e-11
+   -2.065094984297504e-11
+    8.383057788539102e-11
+   -1.320579156738061e-12
+   -9.875061776398978e-12
+    8.385424503709454e-11
+   -9.229200811513253e-13
+   -1.316111472273666e-12
+   -2.065351390668097e-11
+    8.194324469742546e-11
+ 2.81e+10    
+    8.207551992705293e-11
+    -2.06529509964759e-11
+    8.383066045903674e-11
+   -1.324009382529819e-12
+   -9.876578908841989e-12
+    8.385431891245743e-11
+   -9.255628864557947e-13
+   -1.319536422193367e-12
+   -2.065550835614048e-11
+    8.194061605212247e-11
+ 2.82e+10    
+    8.207287498620106e-11
+   -2.065496720963456e-11
+    8.383075209026623e-11
+   -1.327436253851986e-12
+   -9.878108990704478e-12
+    8.385440179615717e-11
+   -9.281842977784918e-13
+    -1.32295808328351e-12
+   -2.065751787014306e-11
+    8.193798349354831e-11
+ 2.83e+10    
+    8.207022577911293e-11
+   -2.065699848254293e-11
+    8.383085258719592e-11
+    -1.33085972654815e-12
+   -9.879652007084925e-12
+    8.385449350000173e-11
+   -9.307842595686573e-13
+   -1.326376411418024e-12
+   -2.065954244945533e-11
+    8.193534682633219e-11
+ 2.84e+10    
+    8.206757211219777e-11
+   -2.065904481460448e-11
+    8.383096175978393e-11
+   -1.334279756721739e-12
+    -9.88120794208577e-12
+    8.385459383764626e-11
+   -9.333627175687585e-13
+   -1.329791362725441e-12
+   -2.066158209415683e-11
+    8.193270585667423e-11
+ 2.85e+10    
+    8.206491379344793e-11
+   -2.066110620454639e-11
+    8.383107941984214e-11
+   -1.337696300716434e-12
+   -9.882776778855242e-12
+    8.385470262459739e-11
+   -9.359196187905836e-13
+   -1.333202893569722e-12
+   -2.066363680365089e-11
+    8.193006039233758e-11
+ 2.86e+10    
+    8.206225063243089e-11
+   -2.066318265043191e-11
+     8.38312053810466e-11
+   -1.341109315097293e-12
+   -9.884358499628111e-12
+    8.385481967821758e-11
+   -9.384549114916651e-13
+   -1.336610960531722e-12
+   -2.066570657667584e-11
+    8.192741024264132e-11
+ 2.87e+10    
+    8.205958244027958e-11
+   -2.066527414967205e-11
+    8.383133945894696e-11
+   -1.344518756632274e-12
+   -9.885953085765583e-12
+    8.385494481772829e-11
+   -9.409685451520971e-13
+   -1.340015520391103e-12
+    -2.06677914113159e-11
+    8.192475521845175e-11
+ 2.88e+10    
+    8.205690902968427e-11
+   -2.066738069903778e-11
+    8.383148147097461e-11
+   -1.347924582274334e-12
+   -9.887560517793983e-12
+    8.385507786421151e-11
+   -9.434604704517472e-13
+   -1.343416530108826e-12
+   -2.066989130501172e-11
+    8.192209513217476e-11
+ 2.89e+10    
+    8.205423021488254e-11
+   -2.066950229467124e-11
+     8.38316312364502e-11
+    -1.35132674914407e-12
+   -9.889180775442731e-12
+    8.385521864061123e-11
+   -9.459306392477799e-13
+   -1.346813946810105e-12
+   -2.067200625457106e-11
+    8.191942979774742e-11
+ 2.9e+10     
+    8.205154581165089e-11
+   -2.067163893209761e-11
+    8.383178857658961e-11
+   -1.354725214512853e-12
+   -9.890813837681124e-12
+    8.385536697173359e-11
+   -9.483790045526327e-13
+   -1.350207727767931e-12
+   -2.067413625617919e-11
+    8.191675903062963e-11
+ 2.91e+10    
+    8.204885563729465e-11
+   -2.067379060623589e-11
+    8.383195331450886e-11
+   -1.358119935786475e-12
+   -9.892459682754278e-12
+    8.385552268424607e-11
+   -9.508055205122557e-13
+   -1.353597830386992e-12
+   -2.067628130540907e-11
+    8.191408264779543e-11
+ 2.92e+10    
+      8.2046159510639e-11
+    -2.06759573114104e-11
+    8.383212527522835e-11
+   -1.361510870489209e-12
+   -9.894118288218038e-12
+    8.385568560667601e-11
+   -9.532101423848214e-13
+   -1.356984212188212e-12
+    -2.06784413972314e-11
+     8.19114004677246e-11
+ 2.93e+10    
+    8.204345725201915e-11
+   -2.067813904136111e-11
+    8.383230428567463e-11
+     -1.3648979762485e-12
+   -9.895789630973017e-12
+    8.385585556940769e-11
+   -9.555928265197331e-13
+   -1.360366830793585e-12
+   -2.068061652602449e-11
+     8.19087123103934e-11
+ 2.94e+10    
+    8.204074868327063e-11
+   -2.068033578925451e-11
+    8.383249017468329e-11
+   -1.368281210780007e-12
+   -9.897473687297674e-12
+    8.385603240467931e-11
+   -9.579535303369885e-13
+    -1.36374564391168e-12
+   -2.068280668558383e-11
+     8.19060179972662e-11
+ 2.95e+10    
+    8.203803362771953e-11
+   -2.068254754769383e-11
+    8.383268277299851e-11
+   -1.371660531873189e-12
+   -9.899170432880423e-12
+    8.385621594657818e-11
+   -9.602922123069329e-13
+   -1.367120609323421e-12
+    -2.06850118691317e-11
+     8.19033173512858e-11
+ 2.96e+10    
+    8.203531191017265e-11
+   -2.068477430872909e-11
+    8.383288191327307e-11
+   -1.375035897377272e-12
+   -9.900879842850949e-12
+    8.385640603103601e-11
+   -9.626088319303546e-13
+   -1.370491684868467e-12
+   -2.068723206932634e-11
+    8.190061019686495e-11
+ 2.97e+10    
+    8.203258335690737e-11
+   -2.068701606386698e-11
+    8.383308743006596e-11
+   -1.378407265187751e-12
+   -9.902601891810426e-12
+    8.385660249582202e-11
+   -9.649033497189165e-13
+   -1.373858828431915e-12
+   -2.068946727827092e-11
+    8.189789635987653e-11
+ 2.98e+10    
+    8.202984779566181e-11
+   -2.068927280408039e-11
+    8.383329915984012e-11
+   -1.381774593233324e-12
+   -9.904336553861131e-12
+    8.385680518053678e-11
+   -9.671757271759465e-13
+   -1.377221997931508e-12
+   -2.069171748752243e-11
+    8.189517566764415e-11
+ 2.99e+10    
+    8.202710505562449e-11
+   -2.069154451981776e-11
+    8.383351694095822e-11
+    -1.38513783946315e-12
+   -9.906083802634899e-12
+    8.385701392660385e-11
+   -9.694259267775943e-13
+   -1.380581151305231e-12
+   -2.069398268810044e-11
+    8.189244794893339e-11
+ 3e+10       
+    8.202435496742404e-11
+   -2.069383120101216e-11
+    8.383374061367811e-11
+   -1.388496961834697e-12
+   -9.907843611320953e-12
+    8.385722857726146e-11
+   -9.716539119542844e-13
+    -1.38393624649934e-12
+   -2.069626287049524e-11
+    8.188971303394123e-11
+ 3.01e+10    
+    8.202159736311924e-11
+   -2.069613283708992e-11
+    8.383397002014602e-11
+   -1.391851918301911e-12
+   -9.909615952692684e-12
+    8.385744897755282e-11
+   -9.738596470725564e-13
+   -1.387287241456785e-12
+   -2.069855802467626e-11
+    8.188697075428711e-11
+ 3.02e+10    
+     8.20188320761882e-11
+   -2.069844941697943e-11
+    8.383420500439029e-11
+   -1.395202666803736e-12
+   -9.911400799133821e-12
+    8.385767497431596e-11
+   -9.760430974172214e-13
+   -1.390634094106043e-12
+   -2.070086814009987e-11
+    8.188422094300314e-11
+ 3.03e+10    
+    8.201605894151837e-11
+    -2.07007809291192e-11
+    8.383444541231305e-11
+   -1.398549165253251e-12
+    -9.91319812266362e-12
+    8.385790641617332e-11
+   -9.782042291738314e-13
+   -1.393976762350333e-12
+   -2.070319320571728e-11
+    8.188146343452372e-11
+ 3.04e+10    
+    8.201327779539564e-11
+   -2.070312736146591e-11
+     8.38346910916807e-11
+   -1.401891371526923e-12
+   -9.915007894961242e-12
+    8.385814315351879e-11
+   -9.803430094115384e-13
+   -1.397315204057232e-12
+   -2.070553320998193e-11
+    8.187869806467676e-11
+ 3.05e+10    
+    8.201048847549421e-11
+   -2.070548870150216e-11
+     8.38349418921146e-11
+   -1.405229243454459e-12
+   -9.916830087389495e-12
+    8.385838503850621e-11
+   -9.824594060662186e-13
+   -1.400649377048622e-12
+   -2.070788814085686e-11
+    8.187592467067241e-11
+ 3.06e+10    
+    8.200769082086578e-11
+     -2.0707864936244e-11
+    8.383519766507953e-11
+   -1.408562738808927e-12
+    -9.91866467101773e-12
+    8.385863192503631e-11
+    -9.84553387923961e-13
+    -1.40397923909104e-12
+   -2.071025798582188e-11
+     8.18731430910942e-11
+ 3.07e+10    
+    8.200488467192901e-11
+   -2.071025605224804e-11
+    8.383545826387203e-11
+   -1.411891815297301e-12
+   -9.920511616643894e-12
+    8.385888366874217e-11
+    -9.86624924604863e-13
+   -1.407304747886393e-12
+   -2.071264273188034e-11
+    8.187035316588823e-11
+ 3.08e+10    
+    8.200206987045878e-11
+   -2.071266203561844e-11
+    8.383572354360729e-11
+   -1.415216430551328e-12
+   -9.922370894815956e-12
+    8.385914012697508e-11
+   -9.886739865471501e-13
+   -1.410625861062987e-12
+   -2.071504236556583e-11
+    8.186755473635363e-11
+ 3.09e+10    
+    8.199924625957543e-11
+   -2.071508287201364e-11
+    8.383599336120586e-11
+   -1.418536542118759e-12
+   -9.924242475852576e-12
+    8.385940115878943e-11
+   -9.907005449916126e-13
+   -1.413942536166957e-12
+   -2.071745687294862e-11
+    8.186474764513183e-11
+ 3.1e+10     
+    8.199641368373441e-11
+    -2.07175185466527e-11
+    8.383626757537873e-11
+   -1.421852107454985e-12
+   -9.926126329863084e-12
+    8.385966662492716e-11
+   -9.927045719663482e-13
+   -1.417254730653927e-12
+   -2.071988623964196e-11
+     8.18619317361969e-11
+ 3.11e+10    
+    8.199357198871512e-11
+   -2.071996904432165e-11
+     8.38365460466122e-11
+   -1.425163083914888e-12
+   -9.928022426766701e-12
+    8.385993638780076e-11
+   -9.946860402718245e-13
+   -1.420562401881171e-12
+     -2.0722330450808e-11
+    8.185910685484502e-11
+ 3.12e+10    
+    8.199072102161019e-11
+   -2.072243434937919e-11
+    8.383682863715154e-11
+    -1.42846942874516e-12
+   -9.929930736311198e-12
+    8.386021031147742e-11
+    -9.96644923466239e-13
+   -1.423865507099895e-12
+    -2.07247894911638e-11
+     8.18562728476843e-11
+ 3.13e+10    
+    8.198786063081511e-11
+   -2.072491444576275e-11
+    8.383711521098437e-11
+    -1.43177109907686e-12
+    -9.93185122809075e-12
+    8.386048826166069e-11
+   -9.985811958511939e-13
+   -1.427164003447999e-12
+   -2.072726334498674e-11
+    8.185342956262441e-11
+ 3.14e+10    
+    8.198499066601693e-11
+   -2.072740931699351e-11
+    8.383740563382256e-11
+   -1.435068051918324e-12
+   -9.933783871563243e-12
+    8.386077010567284e-11
+   -1.000494832457653e-12
+   -1.430457847943054e-12
+   -2.072975199612004e-11
+    8.185057684886649e-11
+ 3.15e+10    
+    8.198211097818357e-11
+   -2.072991894618192e-11
+    8.383769977308453e-11
+   -1.438360244148377e-12
+   -9.935728636067021e-12
+    8.386105571243696e-11
+   -1.002385809032215e-12
+   -1.433746997475622e-12
+   -2.073225542797811e-11
+    8.184771455689258e-11
+ 3.16e+10    
+     8.19792214195533e-11
+   -2.073244331603262e-11
+    8.383799749787556e-11
+   -1.441647632509837e-12
+   -9.937685490836784e-12
+    8.386134495245725e-11
+   -1.004254102023671e-12
+   -1.437031408802811e-12
+   -2.073477362355137e-11
+    8.184484253845533e-11
+ 3.17e+10    
+    8.197632184362353e-11
+   -2.073498240884906e-11
+     8.38382986789686e-11
+   -1.444930173603367e-12
+   -9.939654405019129e-12
+    8.386163769780055e-11
+   -1.006099688569856e-12
+   -1.440311038542236e-12
+   -2.073730656541125e-11
+    8.184196064656775e-11
+ 3.18e+10    
+    8.197341210514025e-11
+   -2.073753620653833e-11
+    8.383860318878427e-11
+   -1.448207823881537e-12
+   -9.941635347687409e-12
+    8.386193382207594e-11
+   -1.007922546484774e-12
+   -1.443585843166138e-12
+   -2.073985423571481e-11
+    8.183906873549263e-11
+ 3.19e+10    
+    8.197049206008714e-11
+   -2.074010469061521e-11
+    8.383891090136939e-11
+   -1.451480539643241e-12
+   -9.943628287856018e-12
+    8.386223320041542e-11
+   -1.009722654246034e-12
+   -1.446855778995814e-12
+   -2.074241661620931e-11
+    8.183616666073249e-11
+ 3.2e+10     
+    8.196756156567481e-11
+   -2.074268784220641e-11
+    8.383922169237628e-11
+   -1.454748277028367e-12
+   -9.945633194494122e-12
+    8.386253570945271e-11
+   -1.011499990982549e-12
+   -1.450120802196379e-12
+   -2.074499368823633e-11
+    8.183325427901876e-11
+ 3.21e+10    
+    8.196462048032989e-11
+   -2.074528564205454e-11
+    8.383953543904074e-11
+     -1.4580109920127e-12
+   -9.947650036538932e-12
+    8.386284122730334e-11
+   -1.013254536462506e-12
+   -1.453380868771697e-12
+   -2.074758543273616e-11
+    8.183033144830178e-11
+ 3.22e+10    
+    8.196166866368454e-11
+    -2.07478980705217e-11
+    8.383985202015985e-11
+   -1.461268640403193e-12
+   -9.949678782908336e-12
+    8.386314963354279e-11
+   -1.014986271081631e-12
+    -1.45663593455964e-12
+   -2.075019183025158e-11
+    8.182739802774037e-11
+ 3.23e+10    
+     8.19587059765654e-11
+   -2.075052510759308e-11
+    8.384017131606904e-11
+   -1.464521177833352e-12
+   -9.951719402513129e-12
+    8.386346080918599e-11
+   -1.016695175851713e-12
+   -1.459885955227542e-12
+   -2.075281286093181e-11
+     8.18244538776913e-11
+ 3.24e+10    
+    8.195573228098307e-11
+   -2.075316673288038e-11
+    8.384049320861937e-11
+   -1.467768559759027e-12
+   -9.953771864268692e-12
+    8.386377463666526e-11
+   -1.018381232389389e-12
+   -1.463130886267951e-12
+   -2.075544850453609e-11
+    8.182149885969894e-11
+ 3.25e+10    
+    8.195274744012126e-11
+   -2.075582292562481e-11
+    8.384081758115379e-11
+   -1.471010741454315e-12
+   -9.955836137106236e-12
+    8.386409099980852e-11
+   -1.020044422905214e-12
+   -1.466370682994582e-12
+   -2.075809874043718e-11
+    8.181853283648526e-11
+ 3.26e+10    
+    8.194975131832615e-11
+   -2.075849366470016e-11
+    8.384114431848346e-11
+   -1.474247678007781e-12
+   -9.957912189983522e-12
+     8.38644097838177e-11
+    -1.02168473019298e-12
+   -1.469605300538535e-12
+   -2.076076354762485e-11
+     8.18155556719393e-11
+ 3.27e+10    
+    8.194674378109596e-11
+   -2.076117892861577e-11
+    8.384147330686418e-11
+   -1.477479324318927e-12
+   -9.959999991895307e-12
+    8.386473087524632e-11
+   -1.023302137619272e-12
+   -1.472834693844675e-12
+   -2.076344290470893e-11
+    8.181256723110661e-11
+ 3.28e+10    
+    8.194372469507004e-11
+   -2.076387869551887e-11
+    8.384180443397074e-11
+   -1.480705635094828e-12
+   -9.962099511883011e-12
+    8.386505416197734e-11
+   -1.024896629113337e-12
+   -1.476058817668359e-12
+   -2.076613678992251e-11
+    8.180956738017951e-11
+ 3.29e+10    
+    8.194069392801867e-11
+    -2.07665929431975e-11
+    8.384213758887385e-11
+   -1.483926564847023e-12
+     -9.9642107190444e-12
+    8.386537953320069e-11
+   -1.026468189157148e-12
+   -1.479277626572214e-12
+   -2.076884518112485e-11
+    8.180655598648655e-11
+ 3.3e+10     
+    8.193765134883191e-11
+   -2.076932164908253e-11
+    8.384247266201454e-11
+   -1.487142067888655e-12
+   -9.966333582542554e-12
+    8.386570687939059e-11
+   -1.028016802775732e-12
+   -1.482491074923304e-12
+   -2.077156805580419e-11
+    8.180353291848224e-11
+ 3.31e+10    
+    8.193459682750975e-11
+   -2.077206479025007e-11
+    8.384280954517926e-11
+   -1.490352098331761e-12
+   -9.968468071614435e-12
+    8.386603609228361e-11
+   -1.029542455527764e-12
+   -1.485699116890366e-12
+   -2.077430539108047e-11
+    8.180049804573719e-11
+ 3.32e+10    
+     8.19315302351516e-11
+   -2.077482234342354e-11
+    8.384314813147524e-11
+   -1.493556610084834e-12
+   -9.970614155579396e-12
+    8.386636706485497e-11
+   -1.031045133496387e-12
+   -1.488901706441312e-12
+   -2.077705716370787e-11
+    8.179745123892749e-11
+ 3.33e+10    
+    8.192845144394538e-11
+    -2.07775942849756e-11
+    8.384348831530472e-11
+   -1.496755556850527e-12
+   -9.972771803846961e-12
+      8.3866699691297e-11
+   -1.032524823280261e-12
+   -1.492098797340919e-12
+   -2.077982335007736e-11
+    8.179439236982526e-11
+ 3.34e+10    
+    8.192536032715803e-11
+   -2.078038059093012e-11
+    8.384382999234024e-11
+   -1.499948892123621e-12
+   -9.974940985924415e-12
+    8.386703386699575e-11
+   -1.033981511984881e-12
+   -1.495290343148722e-12
+   -2.078260392621899e-11
+    8.179132131128791e-11
+ 3.35e+10    
+     8.19222567591243e-11
+   -2.078318123696369e-11
+    8.384417305949885e-11
+   -1.503136569189124e-12
+   -9.977121671424038e-12
+    8.386736948850825e-11
+   -1.035415187214082e-12
+    -1.49847629721706e-12
+   -2.078539886780413e-11
+    8.178823793724857e-11
+ 3.36e+10    
+    8.191914061523704e-11
+   -2.078599619840736e-11
+    8.384451741491722e-11
+   -1.506318541120597e-12
+    -9.97931383007003e-12
+    8.386770645354054e-11
+   -1.036825837061818e-12
+   -1.501656612689367e-12
+    -2.07882081501477e-11
+    8.178514212270604e-11
+ 3.37e+10    
+    8.191601177193724e-11
+   -2.078882545024828e-11
+    8.384486295792582e-11
+    -1.50949476077863e-12
+   -9.981517431705112e-12
+    8.386804466092417e-11
+   -1.038213450104149e-12
+   -1.504831242498558e-12
+    -2.07910317482101e-11
+    8.178203374371472e-11
+ 3.38e+10    
+    8.191287010670318e-11
+    -2.07916689671309e-11
+    8.384520958902414e-11
+   -1.512665180809544e-12
+   -9.983732446296709e-12
+    8.386838401059445e-11
+   -1.039578015391438e-12
+   -1.508000139365672e-12
+   -2.079386963659933e-11
+    8.177891267737497e-11
+ 3.39e+10    
+    8.190971549804133e-11
+   -2.079452672335846e-11
+    8.384555720985475e-11
+   -1.515829753644247e-12
+   -9.985958843943063e-12
+    8.386872440356752e-11
+   -1.040919522440791e-12
+   -1.511163255798646e-12
+   -2.079672178957282e-11
+    8.177577880182296e-11
+ 3.4e+10     
+    8.190654782547526e-11
+   -2.079739869289407e-11
+      8.3845905723179e-11
+   -1.518988431497195e-12
+   -9.988196594878857e-12
+    8.386906574191812e-11
+   -1.042237961228704e-12
+   -1.514320544091257e-12
+   -2.079958818103908e-11
+    8.177263199622128e-11
+ 3.41e+10    
+    8.190336696953688e-11
+   -2.080028484936215e-11
+    8.384625503285104e-11
+   -1.522141166365644e-12
+   -9.990445669480665e-12
+    8.386940792875743e-11
+   -1.043533322183937e-12
+   -1.517471956322216e-12
+   -2.080246878455966e-11
+    8.176947214074903e-11
+ 3.42e+10    
+    8.190017281175559e-11
+   -2.080318516604916e-11
+    8.384660504379345e-11
+   -1.525287910028954e-12
+   -9.992706038272114e-12
+    8.386975086821071e-11
+   -1.044805596180569e-12
+    -1.52061744435445e-12
+   -2.080536357335061e-11
+    8.176629911659197e-11
+ 3.43e+10    
+    8.189696523464901e-11
+   -2.080609961590485e-11
+    8.384695566197204e-11
+   -1.528428614048087e-12
+   -9.994977671928784e-12
+    8.387009446539585e-11
+   -1.046054774531301e-12
+    -1.52375695983452e-12
+   -2.080827252028416e-11
+    8.176311280593329e-11
+ 3.44e+10    
+    8.189374412171309e-11
+   -2.080902817154314e-11
+    8.384730679437176e-11
+   -1.531563229765285e-12
+   -9.997260541282936e-12
+    8.387043862640074e-11
+   -1.047280848980937e-12
+     -1.5268904541922e-12
+   -2.081119559789015e-11
+    8.175991309194406e-11
+ 3.45e+10    
+    8.189050935741275e-11
+   -2.081197080524304e-11
+    8.384765834897138e-11
+   -1.534691708303857e-12
+   -9.999554617327859e-12
+    8.387078325826252e-11
+   -1.048483811700067e-12
+   -1.530017878640165e-12
+   -2.081413277835744e-11
+    8.175669985877302e-11
+ 3.46e+10    
+    8.188726082717195e-11
+   -2.081492748894943e-11
+    8.384801023472001e-11
+   -1.537814000568103e-12
+   -1.000185987122219e-11
+    8.387112826894584e-11
+   -1.049663655278999e-12
+    -1.53313918417389e-12
+   -2.081708403353557e-11
+    8.175347299153869e-11
+ 3.47e+10    
+    8.188399841736392e-11
+   -2.081789819427383e-11
+    8.384836236151271e-11
+   -1.540930057243448e-12
+   -1.000417627429382e-11
+    8.387147356732126e-11
+   -1.050820372721785e-12
+   -1.536254321571618e-12
+   -2.082004933493562e-11
+    8.175023237631803e-11
+ 3.48e+10    
+    8.188072201530257e-11
+   -2.082088289249516e-11
+    8.384871464016639e-11
+   -1.544039828796616e-12
+   -1.000650379804373e-11
+    8.387181906314478e-11
+   -1.051953957440565e-12
+   -1.539363241394522e-12
+    -2.08230286537319e-11
+     8.17469779001388e-11
+ 3.49e+10    
+    8.187743150923259e-11
+   -2.082388155456052e-11
+    8.384906698239699e-11
+   -1.547143265476008e-12
+   -1.000884241414966e-11
+    8.387216466703684e-11
+   -1.053064403250011e-12
+   -1.542465893986946e-12
+   -2.082602196076304e-11
+     8.17437094509697e-11
+ 3.5e+10     
+    8.187412678831999e-11
+   -2.082689415108562e-11
+     8.38494193007954e-11
+    -1.55024031731218e-12
+   -1.001119209446932e-11
+    8.387251029046135e-11
+   -1.054151704361996e-12
+   -1.545562229476839e-12
+   -2.082902922653297e-11
+    8.174042691771105e-11
+ 3.51e+10    
+    8.187080774264326e-11
+   -2.082992065235556e-11
+    8.384977150880494e-11
+   -1.553330934118469e-12
+   -1.001355281104384e-11
+    8.387285584570645e-11
+   -1.055215855380443e-12
+    -1.54865219777623e-12
+   -2.083205042121242e-11
+    8.173713019018599e-11
+ 3.52e+10    
+     8.18674742631843e-11
+   -2.083296102832541e-11
+    8.385012352069851e-11
+   -1.556415065491708e-12
+   -1.001592453610064e-11
+    8.387320124586314e-11
+   -1.056256851296366e-12
+   -1.551735748581919e-12
+   -2.083508551463971e-11
+    8.173381915913136e-11
+ 3.53e+10    
+    8.186412624181892e-11
+   -2.083601524862062e-11
+    8.385047525155592e-11
+   -1.559492660813075e-12
+   -1.001830724205642e-11
+    8.387354640480665e-11
+   -1.057274687483081e-12
+   -1.554812831376201e-12
+   -2.083813447632202e-11
+    8.173049371618892e-11
+ 3.54e+10    
+    8.186076357130831e-11
+   -2.083908328253773e-11
+    8.385082661724244e-11
+   -1.562563669249068e-12
+   -1.002070090151988e-11
+    8.387389123717607e-11
+   -1.058269359691581e-12
+   -1.557883395427789e-12
+   -2.084119727543621e-11
+    8.172715375389614e-11
+ 3.55e+10    
+    8.185738614529001e-11
+    -2.08421650990448e-11
+    8.385117753438652e-11
+    -1.56562803975259e-12
+   -1.002310548729423e-11
+    8.387423565835569e-11
+   -1.059240864046121e-12
+   -1.560947389792762e-12
+      -2.084427388083e-11
+    8.172379916567757e-11
+ 3.56e+10    
+    8.185399385826901e-11
+   -2.084526066678179e-11
+    8.385152792035814e-11
+   -1.568685721064129e-12
+   -1.002552097237962e-11
+    8.387457958445579e-11
+   -1.060189197039946e-12
+   -1.564004763315697e-12
+   -2.084736426102281e-11
+    8.172042984583617e-11
+ 3.57e+10    
+    8.185058660560917e-11
+   -2.084836995406123e-11
+    8.385187769324846e-11
+   -1.571736661713046e-12
+   -1.002794732997551e-11
+    8.387492293229397e-11
+   -1.061114355531211e-12
+   -1.567055464630871e-12
+   -2.085046838420676e-11
+    8.171704568954489e-11
+ 3.58e+10    
+    8.184716428352455e-11
+   -2.085149292886852e-11
+    8.385222677184867e-11
+   -1.574780810018994e-12
+   -1.003038453348269e-11
+    8.387526561937696e-11
+   -1.062016336739038e-12
+   -1.570099442163566e-12
+   -2.085358621824756e-11
+    8.171364659283746e-11
+ 3.59e+10    
+    8.184372678907076e-11
+   -2.085462955886246e-11
+    8.385257507562961e-11
+   -1.577818114093376e-12
+   -1.003283255650543e-11
+    8.387560756388227e-11
+   -1.062895138239763e-12
+   -1.573136644131499e-12
+   -2.085671773068528e-11
+    8.171023245260032e-11
+ 3.6e+10     
+    8.184027402013647e-11
+   -2.085777981137561e-11
+    8.385292252472173e-11
+   -1.580848521841007e-12
+   -1.003529137285326e-11
+     8.38759486846408e-11
+   -1.063750757963335e-12
+   -1.576167018546323e-12
+   -2.085986288873548e-11
+     8.17068031665643e-11
+ 3.61e+10    
+    8.183680587543546e-11
+   -2.086094365341488e-11
+     8.38532690398959e-11
+   -1.583871980961729e-12
+   -1.003776095654284e-11
+    8.387628890111941e-11
+   -1.064583194189888e-12
+   -1.579190513215228e-12
+   -2.086302165928982e-11
+    8.170335863329581e-11
+ 3.62e+10    
+    8.183332225449752e-11
+   -2.086412105166178e-11
+    8.385361454254372e-11
+   -1.586888438952217e-12
+   -1.004024128179959e-11
+    8.387662813340335e-11
+    -1.06539244554645e-12
+   -1.582207075742656e-12
+     -2.0866194008917e-11
+    8.169989875218906e-11
+ 3.63e+10    
+    8.182982305766088e-11
+   -2.086731197247295e-11
+    8.385395895465876e-11
+   -1.589897843107887e-12
+    -1.00427323230592e-11
+    8.387696630217986e-11
+     -1.0661785110038e-12
+   -1.585216653532091e-12
+   -2.086937990386349e-11
+     8.16964234234576e-11
+ 3.64e+10    
+     8.18263081860638e-11
+   -2.087051638188049e-11
+    8.385430219881825e-11
+   -1.592900140524789e-12
+   -1.004523405496922e-11
+    8.387730332872172e-11
+   -1.066941389873519e-12
+    -1.58821919378793e-12
+    -2.08725793100544e-11
+     8.16929325481259e-11
+ 3.65e+10    
+    8.182277754163668e-11
+   -2.087373424559261e-11
+    8.385464419816516e-11
+   -1.595895278101697e-12
+   -1.004774645239028e-11
+    8.387763913487083e-11
+    -1.06768108180514e-12
+   -1.591214643517454e-12
+   -2.087579219309428e-11
+    8.168942602802211e-11
+ 3.66e+10    
+    8.181923102709383e-11
+   -2.087696552899385e-11
+    8.385498487639003e-11
+    -1.59888320254219e-12
+   -1.005026949039745e-11
+     8.38779736430225e-11
+   -1.068397586783491e-12
+   -1.594202949532865e-12
+    -2.08790185182678e-11
+    8.168590376576931e-11
+ 3.67e+10    
+    8.181566854592584e-11
+   -2.088021019714553e-11
+    8.385532415771417e-11
+   -1.601863860356877e-12
+   -1.005280314428135e-11
+    8.387830677611023e-11
+   -1.069090905126126e-12
+   -1.597184058453421e-12
+   -2.088225825054069e-11
+    8.168236566477803e-11
+ 3.68e+10    
+     8.18120900023915e-11
+   -2.088346821478633e-11
+    8.385566196687254e-11
+   -1.604837197865652e-12
+   -1.005534738954929e-11
+    8.387863845758985e-11
+   -1.069761037480972e-12
+   -1.600157916707635e-12
+   -2.088551135456027e-11
+    8.167881162923818e-11
+ 3.69e+10    
+    8.180849530151061e-11
+   -2.088673954633264e-11
+    8.385599822909713e-11
+   -1.607803161200068e-12
+   -1.005790220192624e-11
+    8.387896861142568e-11
+   -1.070407984824053e-12
+    -1.60312447053556e-12
+   -2.088877779465641e-11
+    8.167524156411158e-11
+ 3.7e+10     
+    8.180488434905559e-11
+   -2.089002415587907e-11
+    8.385633287010128e-11
+   -1.610761696305723e-12
+   -1.006046755735577e-11
+     8.38792971620748e-11
+   -1.071031748457373e-12
+   -1.606083665991145e-12
+   -2.089205753484211e-11
+    8.167165537512407e-11
+ 3.71e+10    
+    8.180125705154452e-11
+   -2.089332200719884e-11
+    8.385666581606377e-11
+   -1.613712748944777e-12
+   -1.006304343200093e-11
+    8.387962403447399e-11
+   -1.071632330006939e-12
+   -1.609035448944638e-12
+   -2.089535053881443e-11
+    8.166805296875813e-11
+ 3.72e+10    
+    8.179761331623363e-11
+   -2.089663306374441e-11
+    8.385699699361344e-11
+   -1.616656264698496e-12
+   -1.006562980224503e-11
+     8.38799491540254e-11
+   -1.072209731420928e-12
+    -1.61197976508511e-12
+   -2.089865676995508e-11
+    8.166443425224521e-11
+ 3.73e+10    
+    8.179395305110951e-11
+   -2.089995728864783e-11
+    8.385732632981446e-11
+   -1.619592188969859e-12
+   -1.006822664469228e-11
+    8.388027244658221e-11
+   -1.072763954967953e-12
+   -1.614916559923003e-12
+   -2.090197619133104e-11
+    8.166079913355815e-11
+ 3.74e+10    
+     8.17902761648822e-11
+   -2.090329464472132e-11
+    8.385765375215185e-11
+   -1.622520466986269e-12
+   -1.007083393616855e-11
+    8.388059383843718e-11
+   -1.073295003235485e-12
+   -1.617845778792739e-12
+   -2.090530876569573e-11
+    8.165714752140453e-11
+ 3.75e+10    
+    8.178658256697791e-11
+   -2.090664509445772e-11
+     8.38579791885168e-11
+   -1.625441043802276e-12
+   -1.007345165372182e-11
+    8.388091325630808e-11
+    -1.07380287912839e-12
+   -1.620767366855417e-12
+   -2.090865445548925e-11
+    8.165347932521836e-11
+ 3.76e+10    
+    8.178287216753174e-11
+   -2.091000860003117e-11
+    8.385830256719402e-11
+   -1.628353864302382e-12
+   -1.007607977462288e-11
+    8.388123062732589e-11
+   -1.074287585867596e-12
+   -1.623681269101582e-12
+   -2.091201322283933e-11
+    8.164979445515376e-11
+ 3.77e+10    
+    8.177914487738072e-11
+   -2.091338512329746e-11
+    8.385862381684729e-11
+   -1.631258873203899e-12
+   -1.007871827636561e-11
+    8.388154587902256e-11
+   -1.074749126988871e-12
+   -1.626587430353982e-12
+    -2.09153850295622e-11
+    8.164609282207752e-11
+ 3.78e+10    
+    8.177540060805679e-11
+   -2.091677462579472e-11
+    8.385894286650721e-11
+   -1.634156015059882e-12
+   -1.008136713666756e-11
+    8.388185893931898e-11
+   -1.075187506341738e-12
+   -1.629485795270474e-12
+   -2.091876983716306e-11
+    8.164237433756184e-11
+ 3.79e+10    
+    8.177163927178023e-11
+   -2.092017706874399e-11
+    8.385925964555805e-11
+   -1.637045234262065e-12
+    -1.00840263334701e-11
+    8.388216973651303e-11
+   -1.075602728088488e-12
+   -1.632376308346934e-12
+    -2.09221676068369e-11
+    8.163863891387764e-11
+ 3.8e+10     
+    8.176786078145222e-11
+   -2.092359241304974e-11
+    8.385957408372665e-11
+   -1.639926475043875e-12
+   -1.008669584493902e-11
+    8.388247819926858e-11
+   -1.075994796703322e-12
+     -1.6352589139202e-12
+   -2.092557829946932e-11
+    8.163488646398757e-11
+ 3.81e+10    
+    8.176406505064875e-11
+   -2.092702061930053e-11
+    8.385988611106882e-11
+   -1.642799681483543e-12
+   -1.008937564946448e-11
+    8.388278425660443e-11
+   -1.076363716971622e-12
+   -1.638133556171125e-12
+   -2.092900187563719e-11
+    8.163111690153941e-11
+ 3.82e+10    
+     8.17602519936133e-11
+   -2.093046164776956e-11
+    8.386019565795926e-11
+    -1.64566479750717e-12
+   -1.009206572566139e-11
+    8.388308783788358e-11
+   -1.076709493989282e-12
+   -1.641000179127626e-12
+   -2.093243829560941e-11
+    8.162733014085879e-11
+ 3.83e+10    
+    8.175642152525122e-11
+   -2.093391545841542e-11
+     8.38605026550801e-11
+   -1.648521766891916e-12
+   -1.009476605236959e-11
+    8.388338887280269e-11
+   -1.077032133162205e-12
+   -1.643858726667814e-12
+    -2.09358875193476e-11
+    8.162352609694321e-11
+ 3.84e+10    
+    8.175257356112228e-11
+   -2.093738201088262e-11
+    8.386080703340978e-11
+   -1.651370533269177e-12
+   -1.009747660865385e-11
+    8.388368729138226e-11
+   -1.077331640205887e-12
+   -1.646709142523145e-12
+   -2.093934950650703e-11
+    8.161970468545502e-11
+ 3.85e+10    
+    8.174870801743503e-11
+   -2.094086126450235e-11
+    8.386110872421299e-11
+   -1.654211040127854e-12
+   -1.010019737380411e-11
+    8.388398302395633e-11
+   -1.077608021145091e-12
+   -1.649551370281633e-12
+   -2.094282421643705e-11
+    8.161586582271488e-11
+ 3.86e+10    
+    8.174482481103951e-11
+     -2.0944353178293e-11
+    8.386140765903025e-11
+   -1.657043230817606e-12
+   -1.010292832733534e-11
+    8.388427600116313e-11
+   -1.077861282313636e-12
+   -1.652385353391107e-12
+   -2.094631160818205e-11
+    8.161200942569542e-11
+ 3.87e+10    
+    8.174092385942218e-11
+   -2.094785771096103e-11
+    8.386170376966862e-11
+   -1.659867048552232e-12
+   -1.010566944898768e-11
+    8.388456615393618e-11
+   -1.078091430354311e-12
+   -1.655211035162481e-12
+   -2.094981164048234e-11
+    8.160813541201519e-11
+ 3.88e+10    
+    8.173700508069892e-11
+   -2.095137482090167e-11
+    8.386199698819191e-11
+   -1.662682436412956e-12
+   -1.010842071872632e-11
+    8.388485341349438e-11
+   -1.078298472218848e-12
+   -1.658028358773112e-12
+   -2.095332427177447e-11
+    8.160424369993164e-11
+ 3.89e+10    
+    8.173306839360899e-11
+   -2.095490446619937e-11
+    8.386228724691152e-11
+   -1.665489337351901e-12
+   -1.011118211674149e-11
+    8.388513771133459e-11
+    -1.07848241516801e-12
+   -1.660837267270131e-12
+   -2.095684946019252e-11
+    8.160033420833553e-11
+ 3.9e+10     
+    8.172911371750955e-11
+   -2.095844660462895e-11
+    8.386257447837815e-11
+   -1.668287694195471e-12
+   -1.011395362344825e-11
+    8.388541897922191e-11
+   -1.078643266771788e-12
+   -1.663637703573885e-12
+   -2.096038716356841e-11
+    8.159640685674458e-11
+ 3.91e+10    
+    8.172514097236889e-11
+     -2.0962001193656e-11
+    8.386285861537281e-11
+   -1.671077449647822e-12
+   -1.011673521948648e-11
+    8.388569714918236e-11
+   -1.078781034909681e-12
+   -1.666429610481342e-12
+   -2.096393733943309e-11
+    8.159246156529751e-11
+ 3.92e+10    
+    8.172115007876147e-11
+   -2.096556819043779e-11
+      8.3863139590899e-11
+   -1.673858546294396e-12
+   -1.011952688572057e-11
+    8.388597215349445e-11
+   -1.078895727771062e-12
+   -1.669212930669578e-12
+   -2.096749994501688e-11
+    8.158849825474763e-11
+ 3.93e+10    
+    8.171714095786102e-11
+   -2.096914755182405e-11
+    8.386341733817476e-11
+   -1.676630926605395e-12
+    -1.01223286032393e-11
+    8.388624392468191e-11
+   -1.078987353855638e-12
+   -1.671987606699284e-12
+   -2.097107493725052e-11
+    8.158451684645718e-11
+ 3.94e+10    
+    8.171311353143589e-11
+   -2.097273923435766e-11
+    8.386369179062492e-11
+   -1.679394532939382e-12
+   -1.012514035335554e-11
+    8.388651239550576e-11
+   -1.079055921974005e-12
+   -1.674753581018267e-12
+   -2.097466227276591e-11
+    8.158051726239169e-11
+ 3.95e+10    
+    8.170906772184261e-11
+   -2.097634319427557e-11
+    8.386396288187409e-11
+   -1.682149307546837e-12
+   -1.012796211760601e-11
+    8.388677749895743e-11
+    -1.07910144124829e-12
+   -1.677510795965075e-12
+   -2.097826190789678e-11
+    8.157649942511369e-11
+ 3.96e+10    
+     8.17050034520209e-11
+   -2.097995938750954e-11
+    8.386423054573976e-11
+   -1.684895192573781e-12
+   -1.013079387775099e-11
+     8.38870391682522e-11
+   -1.079123921112867e-12
+   -1.680259193772516e-12
+   -2.098187379867967e-11
+     8.15724632577774e-11
+ 3.97e+10    
+     8.17009206454875e-11
+   -2.098358776968694e-11
+    8.386449471622488e-11
+   -1.687632130065413e-12
+   -1.013363561577393e-11
+    8.388729733682195e-11
+   -1.079123371315158e-12
+   -1.682998716571306e-12
+   -2.098549790085454e-11
+    8.156840868412285e-11
+ 3.98e+10    
+    8.169681922633133e-11
+   -2.098722829613161e-11
+    8.386475532751249e-11
+   -1.690360061969762e-12
+   -1.013648731388115e-11
+    8.388755193830847e-11
+   -1.079099801916536e-12
+   -1.685729306393718e-12
+   -2.098913416986559e-11
+    8.156433562847027e-11
+ 3.99e+10    
+    8.169269911920758e-11
+   -2.099088092186468e-11
+     8.38650123139585e-11
+   -1.693078930141349e-12
+   -1.013934895450143e-11
+    8.388780290655798e-11
+   -1.079053223293277e-12
+   -1.688450905177239e-12
+   -2.099278256086211e-11
+    8.156024401571474e-11
+ 4e+10       
+    8.168856024933281e-11
+   -2.099454560160547e-11
+    8.386526561008631e-11
+   -1.695788676344943e-12
+   -1.014222052028558e-11
+     8.38880501756144e-11
+   -1.078983646137602e-12
+   -1.691163454768246e-12
+   -2.099644302869928e-11
+    8.155613377132053e-11
+ 4.01e+10    
+    8.168440254247951e-11
+   -2.099822228977222e-11
+    8.386551515058105e-11
+   -1.698489242259243e-12
+   -1.014510199410607e-11
+    8.388829367971424e-11
+   -1.078891081458811e-12
+   -1.693866896925716e-12
+   -2.100011552793891e-11
+    8.155200482131575e-11
+ 4.02e+10    
+    8.168022592497093e-11
+   -2.100191094048315e-11
+    8.386576087028406e-11
+   -1.701180569480613e-12
+   -1.014799335905646e-11
+    8.388853335328023e-11
+    -1.07877554058447e-12
+   -1.696561173324984e-12
+   -2.100380001285037e-11
+    8.154785709228741e-11
+ 4.03e+10    
+    8.167603032367593e-11
+   -2.100561150755716e-11
+    8.386600270418747e-11
+   -1.703862599526877e-12
+   -1.015089459845096e-11
+    8.388876913091614e-11
+   -1.078637035161673e-12
+   -1.699246225561437e-12
+   -2.100749643741104e-11
+    8.154369051137513e-11
+ 4.04e+10    
+    8.167181566600409e-11
+   -2.100932394451478e-11
+    8.386624058742972e-11
+   -1.706535273841074e-12
+   -1.015380569582395e-11
+    8.388900094740221e-11
+   -1.078475577158394e-12
+   -1.701921995154323e-12
+    -2.10112047553077e-11
+    8.153950500626727e-11
+ 4.05e+10    
+    8.166758187990054e-11
+   -2.101304820457911e-11
+    8.386647445529024e-11
+   -1.709198533795243e-12
+   -1.015672663492939e-11
+    8.388922873768904e-11
+   -1.078291178864875e-12
+   -1.704588423550529e-12
+   -2.101492491993671e-11
+    8.153530050519473e-11
+ 4.06e+10    
+     8.16633288938411e-11
+   -2.101678424067659e-11
+      8.3866704243185e-11
+    -1.71185232069426e-12
+   -1.015965739974025e-11
+    8.388945243689377e-11
+   -1.078083852895128e-12
+   -1.707245452128341e-12
+   -2.101865688440537e-11
+    8.153107693692654e-11
+ 4.07e+10    
+    8.165905663682745e-11
+     -2.1020532005438e-11
+    8.386692988666276e-11
+   -1.714496575779624e-12
+   -1.016259797444798e-11
+    8.388967198029501e-11
+   -1.077853612188451e-12
+   -1.709893022201304e-12
+   -2.102240060153236e-11
+     8.15268342307645e-11
+ 4.08e+10    
+    8.165476503838231e-11
+    -2.10242914511994e-11
+    8.386715132139994e-11
+   -1.717131240233323e-12
+   -1.016554834346184e-11
+     8.38898873033281e-11
+   -1.077600470011051e-12
+   -1.712531075022003e-12
+   -2.102615602384864e-11
+    8.152257231653815e-11
+ 4.09e+10    
+     8.16504540285447e-11
+   -2.102806253000285e-11
+    8.386736848319747e-11
+   -1.719756255181645e-12
+   -1.016850849140833e-11
+    8.389009834158145e-11
+   -1.077324439957711e-12
+    -1.71515955178594e-12
+   -2.102992310359839e-11
+    8.151829112460036e-11
+ 4.1e+10     
+     8.16461235378652e-11
+   -2.103184519359757e-11
+    8.386758130797659e-11
+   -1.722371561699077e-12
+   -1.017147840313043e-11
+    8.389030503079178e-11
+     -1.0770255359535e-12
+   -1.717778393635365e-12
+   -2.103370179273958e-11
+    8.151399058582182e-11
+ 4.11e+10    
+    8.164177349740154e-11
+   -2.103563939344067e-11
+    8.386778973177531e-11
+   -1.724977100812135e-12
+   -1.017445806368701e-11
+    8.389050730684081e-11
+   -1.076703772255603e-12
+   -1.720387541663114e-12
+   -2.103749204294506e-11
+    8.150967063158678e-11
+ 4.12e+10    
+    8.163740383871366e-11
+   -2.103944508069822e-11
+     8.38679936907453e-11
+   -1.727572813503259e-12
+   -1.017744745835215e-11
+    8.389070510575107e-11
+   -1.076359163455129e-12
+   -1.722986936916526e-12
+    -2.10412938056033e-11
+    8.150533119378847e-11
+ 4.13e+10    
+    8.163301449385984e-11
+   -2.104326220624606e-11
+     8.38681931211485e-11
+   -1.730158640714678e-12
+   -1.018044657261435e-11
+    8.389089836368224e-11
+    -1.07599172447905e-12
+    -1.72557652040128e-12
+   -2.104510703181893e-11
+    8.150097220482372e-11
+ 4.14e+10    
+    8.162860539539164e-11
+   -2.104709072067087e-11
+    8.386838795935372e-11
+   -1.732734523352327e-12
+   -1.018345539217581e-11
+    8.389108701692809e-11
+   -1.075601470592122e-12
+   -1.728156233085289e-12
+   -2.104893167241405e-11
+    8.149659359758922e-11
+ 4.15e+10    
+    8.162417647634963e-11
+   -2.105093057427083e-11
+    8.386857814183447e-11
+   -1.735300402289714e-12
+   -1.018647390295168e-11
+     8.38912710019124e-11
+   -1.075188417398943e-12
+   -1.730726015902613e-12
+   -2.105276767792851e-11
+    8.149219530547613e-11
+ 4.16e+10    
+    8.161972767025937e-11
+   -2.105478171705692e-11
+    8.386876360516551e-11
+   -1.737856218371854e-12
+   -1.018950209106928e-11
+    8.389145025518672e-11
+    -1.07475258084598e-12
+   -1.733285809757326e-12
+    -2.10566149986212e-11
+    8.148777726236635e-11
+ 4.17e+10    
+    8.161525891112695e-11
+   -2.105864409875358e-11
+    8.386894428602039e-11
+   -1.740401912419138e-12
+   -1.019253994286727e-11
+    8.389162471342643e-11
+   -1.074293977223709e-12
+    -1.73583555552744e-12
+   -2.106047358447051e-11
+    8.148333940262762e-11
+ 4.18e+10    
+    8.161077013343457e-11
+   -2.106251766879971e-11
+    8.386912012116953e-11
+   -1.742937425231284e-12
+   -1.019558744489485e-11
+    8.389179431342848e-11
+   -1.073812623168772e-12
+   -1.738375194068808e-12
+   -2.106434338517534e-11
+    8.147888166110947e-11
+ 4.19e+10    
+    8.160626127213699e-11
+   -2.106640237634977e-11
+    8.386929104747716e-11
+   -1.745462697591215e-12
+   -1.019864458391093e-11
+    8.389195899210834e-11
+   -1.073308535666191e-12
+   -1.740904666219017e-12
+   -2.106822435015587e-11
+    8.147440397313856e-11
+ 4.2e+10     
+    8.160173226265651e-11
+    -2.10702981702744e-11
+     8.38694570018998e-11
+   -1.747977670268999e-12
+    -1.02017113468832e-11
+     8.38921186864972e-11
+   -1.072781732051621e-12
+   -1.743423912801337e-12
+   -2.107211642855436e-11
+    8.146990627451471e-11
+ 4.21e+10    
+    8.159718304087977e-11
+   -2.107420499916171e-11
+    8.386961792148357e-11
+   -1.750482284025748e-12
+   -1.020478772098733e-11
+    8.389227333373965e-11
+   -1.072232230013663e-12
+   -1.745932874628592e-12
+    -2.10760195692359e-11
+    8.146538850150643e-11
+ 4.22e+10    
+    8.159261354315324e-11
+   -2.107812281131792e-11
+    8.386977374336286e-11
+   -1.752976479617558e-12
+   -1.020787369360601e-11
+    8.389242287109121e-11
+   -1.071660047596199e-12
+   -1.748431492507116e-12
+   -2.107993372078933e-11
+    8.146085059084712e-11
+ 4.23e+10    
+    8.158802370627943e-11
+   -2.108205155476848e-11
+    8.386992440475816e-11
+   -1.755460197799398e-12
+   -1.021096925232804e-11
+    8.389256723591598e-11
+   -1.071065203200792e-12
+   -1.750919707240637e-12
+   -2.108385883152795e-11
+     8.14562924797304e-11
+ 4.24e+10    
+    8.158341346751295e-11
+   -2.108599117725898e-11
+    8.387006984297455e-11
+   -1.757933379329058e-12
+   -1.021407438494741e-11
+    8.389270636568447e-11
+   -1.070447715589101e-12
+    -1.75339745963421e-12
+   -2.108779484949043e-11
+    8.145171410580668e-11
+ 4.25e+10    
+    8.157878276455665e-11
+   -2.108994162625597e-11
+    8.387020999539993e-11
+    -1.76039596497102e-12
+   -1.021718907946232e-11
+    8.389284019797155e-11
+   -1.069807603885371e-12
+   -1.755864690498126e-12
+   -2.109174172244146e-11
+    8.144711540717884e-11
+ 4.26e+10    
+    8.157413153555776e-11
+   -2.109390284894799e-11
+    8.387034479950364e-11
+   -1.762847895500453e-12
+    -1.02203133240742e-11
+    8.389296867045433e-11
+     -1.0691448875789e-12
+   -1.758321340651819e-12
+   -2.109569939787277e-11
+    8.144249632239818e-11
+ 4.27e+10    
+    8.156945971910467e-11
+   -2.109787479224662e-11
+    8.387047419283532e-11
+   -1.765289111707028e-12
+   -1.022344710718675e-11
+    8.389309172091046e-11
+   -1.068459586526622e-12
+   -1.760767350927778e-12
+   -2.109966782300361e-11
+    8.143785679046055e-11
+ 4.28e+10    
+    8.156476725422202e-11
+   -2.110185740278712e-11
+    8.387059811302308e-11
+   -1.767719554398871e-12
+   -1.022659041740484e-11
+    8.389320928721614e-11
+   -1.067751720955648e-12
+   -1.763202662175468e-12
+   -2.110364694478193e-11
+    8.143319675080281e-11
+ 4.29e+10    
+    8.156005408036833e-11
+   -2.110585062692951e-11
+    8.387071649777296e-11
+   -1.770139164406488e-12
+   -1.022974324353358e-11
+    8.389332130734461e-11
+   -1.067021311465898e-12
+   -1.765627215265206e-12
+   -2.110763670988488e-11
+    8.142851614329867e-11
+ 4.3e+10     
+    8.155532013743163e-11
+   -2.110985441075956e-11
+     8.38708292848673e-11
+   -1.772547882586625e-12
+   -1.023290557457717e-11
+    8.389342771936445e-11
+   -1.066268379032731e-12
+   -1.768040951092066e-12
+   -2.111163706471967e-11
+    8.142381490825485e-11
+ 4.31e+10    
+    8.155056536572599e-11
+   -2.111386870008964e-11
+    8.387093641216433e-11
+   -1.774945649826179e-12
+   -1.023607739973794e-11
+    8.389352846143782e-11
+   -1.065492945009614e-12
+   -1.770443810579804e-12
+   -2.111564795542449e-11
+    8.141909298640794e-11
+ 4.32e+10    
+    8.154578970598823e-11
+   -2.111789344045956e-11
+    8.387103781759624e-11
+    -1.77733240704608e-12
+   -1.023925870841515e-11
+    8.389362347181967e-11
+   -1.064695031130823e-12
+   -1.772835734684668e-12
+   -2.111966932786915e-11
+    8.141435031891999e-11
+ 4.33e+10    
+    8.154099309937435e-11
+   -2.112192857713761e-11
+    8.387113343916945e-11
+   -1.779708095205186e-12
+   -1.024244949020395e-11
+    8.389371268885547e-11
+   -1.063874659514186e-12
+   -1.775216664399367e-12
+   -2.112370112765585e-11
+     8.14095868473753e-11
+ 4.34e+10    
+    8.153617548745581e-11
+   -2.112597405512139e-11
+     8.38712232149633e-11
+    -1.78207265530413e-12
+    -1.02456497348943e-11
+    8.389379605098072e-11
+   -1.063031852663813e-12
+   -1.777586540756878e-12
+   -2.112774330012012e-11
+    8.140480251377688e-11
+ 4.35e+10    
+     8.15313368122166e-11
+   -2.113002981913879e-11
+     8.38713070831292e-11
+   -1.784426028389207e-12
+   -1.024885943246967e-11
+    8.389387349671918e-11
+   -1.062166633472895e-12
+   -1.779945304834347e-12
+   -2.113179579033139e-11
+    8.139999726054274e-11
+ 4.36e+10    
+    8.152647701604949e-11
+   -2.113409581364879e-11
+    8.387138498189048e-11
+   -1.786768155556237e-12
+   -1.025207857310612e-11
+    8.389394496468222e-11
+   -1.061279025226506e-12
+   -1.782292897756917e-12
+   -2.113585854309399e-11
+    8.139517103050249e-11
+ 4.37e+10    
+     8.15215960417528e-11
+   -2.113817198284241e-11
+    8.387145684954118e-11
+   -1.789098977954398e-12
+   -1.025530714717091e-11
+    8.389401039356736e-11
+   -1.060369051604405e-12
+    -1.78462926070161e-12
+   -2.113993150294772e-11
+    8.139032376689365e-11
+ 4.38e+10    
+    8.151669383252768e-11
+   -2.114225827064365e-11
+    8.387152262444607e-11
+   -1.791418436790071e-12
+   -1.025854514522144e-11
+    8.389406972215726e-11
+   -1.059436736683929e-12
+   -1.786954334901134e-12
+   -2.114401461416871e-11
+    8.138545541335881e-11
+ 4.39e+10    
+    8.151177033197363e-11
+   -2.114635462071021e-11
+    8.387158224504003e-11
+   -1.793726473330666e-12
+   -1.026179255800399e-11
+    8.389412288931892e-11
+   -1.058482104942814e-12
+   -1.789268061647721e-12
+   -2.114810782077017e-11
+    8.138056591394168e-11
+ 4.4e+10     
+    8.150682548408677e-11
+   -2.115046097643469e-11
+    8.387163564982761e-11
+   -1.796023028908469e-12
+   -1.026504937645255e-11
+    8.389416983400297e-11
+   -1.057505181262113e-12
+    -1.79157038229696e-12
+   -2.115221106650323e-11
+    8.137565521308395e-11
+ 4.41e+10    
+    8.150185923325587e-11
+   -2.115457728094505e-11
+    8.387168277738247e-11
+   -1.798308044924422e-12
+    -1.02683155916875e-11
+    8.389421049524233e-11
+   -1.056505990929093e-12
+   -1.793861238271579e-12
+   -2.115632429485751e-11
+    8.137072325562204e-11
+ 4.42e+10    
+    8.149687152425914e-11
+   -2.115870347710592e-11
+    8.387172356634792e-11
+   -1.800581462851919e-12
+   -1.027159119501446e-11
+    8.389424481215181e-11
+   -1.055484559640134e-12
+   -1.796140571065263e-12
+   -2.116044744906213e-11
+     8.13657699867842e-11
+ 4.43e+10    
+    8.149186230226143e-11
+   -2.116283950751907e-11
+    8.387175795543543e-11
+   -1.802843224240615e-12
+   -1.027487617792294e-11
+    8.389427272392741e-11
+   -1.054440913503695e-12
+   -1.798408322246425e-12
+   -2.116458047208615e-11
+    8.136079535218641e-11
+ 4.44e+10    
+    8.148683151281138e-11
+   -2.116698531452454e-11
+    8.387178588342536e-11
+   -1.805093270720197e-12
+   -1.027817053208508e-11
+    8.389429416984525e-11
+   -1.053375079043251e-12
+   -1.800664433462001e-12
+   -2.116872330663964e-11
+    8.135579929783035e-11
+ 4.45e+10    
+    8.148177910183818e-11
+    -2.11711408402015e-11
+     8.38718072891665e-11
+   -1.807331544004126e-12
+   -1.028147424935437e-11
+    8.389430908926142e-11
+   -1.052287083200233e-12
+   -1.802908846441148e-12
+   -2.117287589517418e-11
+    8.135078177009913e-11
+ 4.46e+10    
+    8.147670501564836e-11
+   -2.117530602636888e-11
+    8.387182211157578e-11
+   -1.809557985893397e-12
+   -1.028478732176432e-11
+    8.389431742161127e-11
+   -1.051176953337046e-12
+   -1.805141502999068e-12
+   -2.117703817988381e-11
+    8.134574271575531e-11
+ 4.47e+10    
+    8.147160920092338e-11
+   -2.117948081458652e-11
+    8.387183028963875e-11
+   -1.811772538280291e-12
+   -1.028810974152711e-11
+     8.38943191064084e-11
+       -1.05004471724e-12
+   -1.807362345040696e-12
+   -2.118121010270554e-11
+     8.13406820819369e-11
+ 4.48e+10    
+    8.146649160471628e-11
+   -2.118366514615565e-11
+     8.38718317624085e-11
+   -1.813975143152071e-12
+    -1.02914415010323e-11
+    8.389431408324491e-11
+   -1.048890403122333e-12
+   -1.809571314564414e-12
+   -2.118539160532029e-11
+    8.133559981615495e-11
+ 4.49e+10    
+    8.146135217444946e-11
+   -2.118785896212023e-11
+    8.387182646900702e-11
+   -1.816165742594707e-12
+   -1.029478259284546e-11
+    8.389430229179048e-11
+    -1.04771403962721e-12
+   -1.811768353665786e-12
+   -2.118958262915347e-11
+    8.133049586629033e-11
+ 4.5e+10     
+     8.14561908579109e-11
+   -2.119206220326725e-11
+    8.387181434862385e-11
+   -1.818344278796543e-12
+   -1.029813300970671e-11
+     8.38942836717919e-11
+    -1.04651565583071e-12
+   -1.813953404541211e-12
+   -2.119378311537583e-11
+    8.132537018059085e-11
+ 4.51e+10    
+    8.145100760325224e-11
+   -2.119627481012798e-11
+    8.387179534051704e-11
+   -1.820510694052028e-12
+   -1.030149274452947e-11
+    8.389425816307307e-11
+    -1.04529528124485e-12
+   -1.816126409491621e-12
+   -2.119799300490411e-11
+    8.132022270766825e-11
+ 4.52e+10    
+    8.144580235898551e-11
+   -2.120049672297853e-11
+    8.387176938401287e-11
+   -1.822664930765312e-12
+   -1.030486179039897e-11
+    8.389422570553407e-11
+   -1.044052945820595e-12
+    -1.81828731092614e-12
+   -2.120221223840181e-11
+    8.131505339649552e-11
+ 4.53e+10    
+    8.144057507398083e-11
+   -2.120472788184081e-11
+    8.387173641850592e-11
+    -1.82480693145395e-12
+   -1.030824014057085e-11
+    8.389418623915154e-11
+   -1.042788679950867e-12
+   -1.820436051365693e-12
+   -2.120644075627989e-11
+    8.130986219640385e-11
+ 4.54e+10    
+    8.143532569746321e-11
+    -2.12089682264833e-11
+    8.387169638345926e-11
+   -1.826936638752476e-12
+   -1.031162778846976e-11
+    8.389413970397764e-11
+   -1.041502514473588e-12
+   -1.822572573446689e-12
+   -2.121067849869743e-11
+    8.130464905708014e-11
+ 4.55e+10    
+    8.143005417901042e-11
+   -2.121321769642191e-11
+    8.387164921840466e-11
+    -1.82905399541607e-12
+   -1.031502472768791e-11
+    8.389408604014057e-11
+   -1.040194480674677e-12
+   -1.824696819924556e-12
+   -2.121492540556248e-11
+    8.129941392856377e-11
+ 4.56e+10    
+    8.142476046854976e-11
+   -2.121747623092066e-11
+    8.387159486294265e-11
+   -1.831158944324134e-12
+   -1.031843095198359e-11
+    8.389402518784359e-11
+   -1.038864610291067e-12
+   -1.826808733677421e-12
+   -2.121918141653266e-11
+    8.129415676124428e-11
+ 4.57e+10    
+    8.141944451635613e-11
+   -2.122174376899266e-11
+    8.387153325674274e-11
+   -1.833251428483867e-12
+   -1.032184645527973e-11
+    8.389395708736539e-11
+   -1.037512935513733e-12
+   -1.828908257709594e-12
+   -2.122344647101587e-11
+    8.128887750585813e-11
+ 4.58e+10    
+    8.141410627304896e-11
+   -2.122602024940076e-11
+    8.387146433954339e-11
+   -1.835331391033811e-12
+   -1.032527123166245e-11
+    8.389388167905961e-11
+   -1.036139488990709e-12
+   -1.830995335155185e-12
+   -2.122772050817113e-11
+    8.128357611348703e-11
+ 4.59e+10    
+    8.140874568958984e-11
+   -2.123030561065842e-11
+    8.387138805115271e-11
+   -1.837398775247439e-12
+   -1.032870527537953e-11
+    8.389379890335477e-11
+   -1.034744303830091e-12
+   -1.833069909281634e-12
+   -2.123200346690911e-11
+    8.127825253555422e-11
+ 4.6e+10     
+    8.140336271728019e-11
+   -2.123459979103051e-11
+    8.387130433144825e-11
+   -1.839453524536636e-12
+   -1.033214858083888e-11
+     8.38937087007541e-11
+    -1.03332741360303e-12
+   -1.835131923493211e-12
+   -2.123629528589293e-11
+    8.127290672382234e-11
+ 4.61e+10    
+    8.139795730775853e-11
+   -2.123890272853408e-11
+    8.387121312037724e-11
+   -1.841495582455261e-12
+   -1.033560114260708e-11
+    8.389361101183542e-11
+   -1.031888852346756e-12
+   -1.837181321334526e-12
+   -2.124059590353884e-11
+     8.12675386303908e-11
+ 4.62e+10    
+    8.139252941299787e-11
+   -2.124321436093903e-11
+    8.387111435795724e-11
+   -1.843524892702558e-12
+   -1.033906295540787e-11
+    8.389350577725111e-11
+   -1.030428654567547e-12
+   -1.839218046494024e-12
+   -2.124490525801694e-11
+    8.126214820769337e-11
+ 4.63e+10    
+    8.138707898530385e-11
+    -2.12475346257691e-11
+     8.38710079842761e-11
+   -1.845541399126704e-12
+   -1.034253401412056e-11
+    8.389339293772789e-11
+   -1.028946855243724e-12
+    -1.84124204280744e-12
+   -2.124922328725178e-11
+    8.125673540849523e-11
+ 4.64e+10    
+    8.138160597731202e-11
+   -2.125186346030255e-11
+    8.387089393949209e-11
+   -1.847545045728206e-12
+   -1.034601431377847e-11
+    8.389327243406708e-11
+   -1.027443489828621e-12
+   -1.843253254261234e-12
+   -2.125354992892326e-11
+    8.125130018589109e-11
+ 4.65e+10    
+    8.137611034198514e-11
+   -2.125620080157282e-11
+    8.387077216383458e-11
+   -1.849535776663371e-12
+   -1.034950384956747e-11
+    8.389314420714413e-11
+   -1.025918594253538e-12
+   -1.845251624996026e-12
+   -2.125788512046714e-11
+    8.124584249330231e-11
+ 4.66e+10    
+    8.137059203261164e-11
+   -2.126054658636944e-11
+    8.387064259760372e-11
+   -1.851513536247688e-12
+   -1.035300261682429e-11
+    8.389300819790889e-11
+   -1.024372204930711e-12
+   -1.847237099309994e-12
+   -2.126222879907572e-11
+     8.12403622844743e-11
+ 4.67e+10    
+    8.136505100280226e-11
+   -2.126490075123873e-11
+    8.387050518117145e-11
+   -1.853478268959221e-12
+   -1.035651061103503e-11
+    8.389286434738553e-11
+   -1.022804358756226e-12
+    -1.84920962166227e-12
+   -2.126658090169865e-11
+    8.123485951347457e-11
+ 4.68e+10    
+    8.135948720648893e-11
+   -2.126926323248461e-11
+    8.387035985498143e-11
+   -1.855429919442015e-12
+   -1.036002782783351e-11
+     8.38927125966724e-11
+   -1.021215093112966e-12
+    -1.85116913667629e-12
+   -2.127094136504364e-11
+    8.122933413469021e-11
+ 4.69e+10    
+    8.135390059792144e-11
+   -2.127363396616932e-11
+     8.38702065595493e-11
+   -1.857368432509388e-12
+   -1.036355426299974e-11
+    8.389255288694226e-11
+   -1.019604445873504e-12
+   -1.853115589143137e-12
+   -2.127531012557692e-11
+    8.122378610282513e-11
+ 4.7e+10     
+    8.134829113166595e-11
+   -2.127801288811418e-11
+    8.387004523546305e-11
+   -1.859293753147329e-12
+   -1.036708991245821e-11
+    8.389238515944215e-11
+   -1.017972455402995e-12
+   -1.855048924024877e-12
+   -2.127968711952418e-11
+    8.121821537289842e-11
+ 4.71e+10    
+    8.134265876260223e-11
+   -2.128239993390027e-11
+    8.386987582338326e-11
+   -1.861205826517729e-12
+   -1.037063477227638e-11
+    8.389220935549345e-11
+    -1.01631916056207e-12
+   -1.856969086457841e-12
+   -2.128407228287111e-11
+    8.121262190024153e-11
+ 4.72e+10    
+    8.133700344592194e-11
+   -2.128679503886938e-11
+    8.386969826404358e-11
+   -1.863104597961742e-12
+   -1.037418883866297e-11
+    8.389202541649214e-11
+   -1.014644600709677e-12
+   -1.858876021755907e-12
+   -2.128846555136421e-11
+    8.120700564049605e-11
+ 4.73e+10    
+    8.133132513712606e-11
+   -2.129119813812447e-11
+    8.386951249825084e-11
+   -1.864990013003001e-12
+   -1.037775210796636e-11
+    8.389183328390828e-11
+   -1.012948815705919e-12
+   -1.860769675413786e-12
+   -2.129286686051125e-11
+     8.12013665496116e-11
+ 4.74e+10    
+    8.132562379202321e-11
+   -2.129560916653073e-11
+    8.386931846688558e-11
+   -1.866862017350896e-12
+   -1.038132457667296e-11
+    8.389163289928671e-11
+   -1.011231845914885e-12
+   -1.862649993110204e-12
+    -2.12972761455822e-11
+     8.11957045838436e-11
+ 4.75e+10    
+    8.131989936672685e-11
+   -2.130002805871605e-11
+    8.386911611090217e-11
+   -1.868720556903762e-12
+    -1.03849062414055e-11
+    8.389142420424687e-11
+   -1.009493732207443e-12
+   -1.864516920711163e-12
+   -2.130169334160981e-11
+    8.119001969975105e-11
+ 4.76e+10    
+    8.131415181765386e-11
+    -2.13044547490719e-11
+    8.386890537132923e-11
+   -1.870565577752103e-12
+   -1.038849709892144e-11
+    8.389120714048264e-11
+   -1.007734515964005e-12
+   -1.866370404273124e-12
+   -2.130611838339022e-11
+    8.118431185419424e-11
+ 4.77e+10    
+    8.130838110152199e-11
+   -2.130888917175409e-11
+    8.386868618926985e-11
+    -1.87239702618176e-12
+   -1.039209714611122e-11
+     8.38909816497628e-11
+   -1.005954239077299e-12
+   -1.868210390046144e-12
+   -2.131055120548374e-11
+    8.117858100433249e-11
+ 4.78e+10    
+    8.130258717534804e-11
+   -2.131333126068338e-11
+    8.386845850590191e-11
+    -1.87421484867709e-12
+   -1.039570637999667e-11
+    8.389074767393097e-11
+   -1.004152943955073e-12
+   -1.870036824477063e-12
+   -2.131499174221554e-11
+    8.117282710762243e-11
+ 4.79e+10    
+    8.129676999644592e-11
+   -2.131778094954639e-11
+    8.386822226247866e-11
+   -1.876018991924052e-12
+   -1.039932479772925e-11
+    8.389050515490558e-11
+   -1.002330673522833e-12
+   -1.871849654212598e-12
+   -2.131943992767633e-11
+    8.116705012181569e-11
+ 4.8e+10     
+    8.129092952242406e-11
+   -2.132223817179613e-11
+    8.386797740032867e-11
+   -1.877809402813359e-12
+    -1.04029523965884e-11
+     8.38902540346801e-11
+    -1.00048747122648e-12
+   -1.873648826102478e-12
+    -2.13238956957229e-11
+    8.116125000495657e-11
+ 4.81e+10    
+    8.128506571118416e-11
+   -2.132670286065289e-11
+    8.386772386085611e-11
+   -1.879586028443553e-12
+   -1.040658917397983e-11
+    8.388999425532314e-11
+   -9.986233810349898e-13
+   -1.875434287202469e-12
+   -2.132835897997896e-11
+    8.115542671538003e-11
+ 4.82e+10    
+      8.1279178520919e-11
+   -2.133117494910504e-11
+    8.386746158554149e-11
+   -1.881348816124055e-12
+    -1.04102351274338e-11
+     8.38897257589785e-11
+   -9.967384474430306e-13
+   -1.877205984777478e-12
+   -2.133282971383588e-11
+    8.114958021171028e-11
+ 4.83e+10    
+    8.127326791010981e-11
+    -2.13356543699094e-11
+    8.386719051594144e-11
+   -1.883097713378226e-12
+   -1.041389025460342e-11
+    8.388944848786517e-11
+   -9.948327154735415e-13
+   -1.878963866304563e-12
+   -2.133730783045316e-11
+    8.114371045285772e-11
+ 4.84e+10    
+    8.126733383752544e-11
+   -2.134014105559242e-11
+    8.386691059368933e-11
+   -1.884832667946376e-12
+   -1.041755455326294e-11
+    8.388916238427779e-11
+   -9.929062306803198e-13
+   -1.880707879475934e-12
+    -2.13417932627593e-11
+    8.113781739801781e-11
+ 4.85e+10    
+     8.12613762622195e-11
+   -2.134463493845065e-11
+    8.386662176049553e-11
+   -1.886553627788745e-12
+     -1.0421228021306e-11
+    8.388886739058646e-11
+   -9.909590391505261e-13
+   -1.882437972201968e-12
+   -2.134628594345236e-11
+    8.113190100666846e-11
+ 4.86e+10    
+    8.125539514352918e-11
+   -2.134913595055155e-11
+    8.386632395814747e-11
+   -1.888260541088512e-12
+   -1.042491065674393e-11
+    8.388856344923664e-11
+   -9.889911875072236e-13
+   -1.884154092614121e-12
+    -2.13507858050008e-11
+    8.112596123856863e-11
+ 4.87e+10    
+    8.124939044107288e-11
+   -2.135364402373417e-11
+     8.38660171285103e-11
+   -1.889953356254691e-12
+   -1.042860245770398e-11
+    8.388825050275007e-11
+   -9.870027229118044e-13
+   -1.885856189067913e-12
+   -2.135529277964406e-11
+    8.111999805375604e-11
+ 4.88e+10    
+    8.124336211474837e-11
+   -2.135815908960991e-11
+    8.386570121352667e-11
+   -1.891632021925087e-12
+   -1.043230342242763e-11
+    8.388792849372398e-11
+    -9.84993693066464e-13
+   -1.887544210145791e-12
+   -2.135980679939329e-11
+    8.111401141254515e-11
+ 4.89e+10    
+    8.123731012473111e-11
+   -2.136268107956326e-11
+    8.386537615521738e-11
+    -1.89329648696919e-12
+   -1.043601354926875e-11
+    8.388759736483152e-11
+    -9.82964146216568e-13
+   -1.889218104660066e-12
+   -2.136432779603192e-11
+    8.110800127552543e-11
+ 4.9e+10     
+    8.123123443147279e-11
+   -2.136720992475259e-11
+    8.386504189568158e-11
+   -1.894946700491036e-12
+   -1.043973283669194e-11
+    8.388725705882224e-11
+   -9.809141311530519e-13
+   -1.890877821655762e-12
+   -2.136885570111667e-11
+    8.110196760355973e-11
+ 4.91e+10    
+    8.122513499569848e-11
+   -2.137174555611078e-11
+    8.386469837709702e-11
+   -1.896582611832073e-12
+   -1.044346128327076e-11
+    8.388690751852167e-11
+   -9.788436972147159e-13
+    -1.89252331041343e-12
+   -2.137339044597791e-11
+    8.109591035778168e-11
+ 4.92e+10    
+    8.121901177840593e-11
+   -2.137628790434597e-11
+     8.38643455417202e-11
+   -1.898204170573981e-12
+   -1.044719888768595e-11
+     8.38865486868319e-11
+   -9.767528942905564e-13
+   -1.894154520451989e-12
+   -2.137793196172053e-11
+    8.108982949959467e-11
+ 4.93e+10    
+    8.121286474086317e-11
+   -2.138083689994235e-11
+    8.386398333188655e-11
+   -1.899811326541464e-12
+   -1.045094564872357e-11
+    8.388618050673123e-11
+   -9.746417728219842e-13
+   -1.895771401531517e-12
+   -2.138248017922474e-11
+    8.108372499066955e-11
+ 4.94e+10    
+    8.120669384460692e-11
+    -2.13853924731609e-11
+    8.386361169001104e-11
+   -1.901404029805044e-12
+   -1.045470156527348e-11
+    8.388580292127461e-11
+   -9.725103838050675e-13
+   -1.897373903656004e-12
+   -2.138703502914647e-11
+    8.107759679294279e-11
+ 4.95e+10    
+    8.120049905144097e-11
+   -2.138995455404013e-11
+      8.3863230558588e-11
+   -1.902982230683806e-12
+   -1.045846663632729e-11
+    8.388541587359367e-11
+     -9.7035877879269e-13
+   -1.898961977076115e-12
+   -2.139159644191838e-11
+    8.107144486861487e-11
+ 4.96e+10    
+    8.119428032343401e-11
+   -2.139452307239668e-11
+    8.386283988019166e-11
+   -1.904545879748105e-12
+   -1.046224086097678e-11
+    8.388501930689671e-11
+   -9.681870098967106e-13
+   -1.900535572291869e-12
+   -2.139616434775049e-11
+    8.106526918014851e-11
+ 4.97e+10    
+    8.118803762291864e-11
+   -2.139909795782629e-11
+    8.386243959747593e-11
+   -1.906094927822313e-12
+   -1.046602423841199e-11
+    8.388461316446923e-11
+   -9.659951297900292e-13
+   -1.902094640055378e-12
+   -2.140073867663085e-11
+    8.105906969026678e-11
+ 4.98e+10    
+    8.118177091248895e-11
+   -2.140367913970444e-11
+    8.386202965317539e-11
+   -1.907629325987464e-12
+   -1.046981676791957e-11
+    8.388419738967337e-11
+     -9.6378319170866e-13
+   -1.903639131373484e-12
+   -2.140531935832625e-11
+    8.105284636195111e-11
+ 4.99e+10    
+    8.117548015499929e-11
+   -2.140826654718702e-11
+    8.386160999010461e-11
+   -1.909149025583911e-12
+   -1.047361844888085e-11
+    8.388377192594855e-11
+   -9.615512494537455e-13
+   -1.905168997510418e-12
+   -2.140990632238299e-11
+    8.104659915844035e-11
+ 5e+10       
+    8.116916531356227e-11
+    -2.14128601092112e-11
+    8.386118055115904e-11
+   -1.910653978213946e-12
+   -1.047742928077019e-11
+     8.38833367168113e-11
+   -9.592993573935002e-13
+    -1.90668418999039e-12
+   -2.141449949812763e-11
+    8.104032804322814e-11
+ 5.01e+10    
+    8.116282635154761e-11
+   -2.141745975449616e-11
+    8.386074127931488e-11
+   -1.912144135744433e-12
+   -1.048124926315307e-11
+    8.388289170585563e-11
+   -9.570275704651647e-13
+   -1.908184660600226e-12
+   -2.141909881466773e-11
+    8.103403298006196e-11
+ 5.02e+10    
+     8.11564632325798e-11
+   -2.142206541154381e-11
+    8.386029211762901e-11
+   -1.913619450309362e-12
+   -1.048507839568439e-11
+    8.388243683675287e-11
+   -9.547359441768479e-13
+   -1.909670361391881e-12
+   -2.142370420089242e-11
+     8.10277139329406e-11
+ 5.03e+10    
+    8.115007592053731e-11
+   -2.142667700863964e-11
+    8.385983300924002e-11
+   -1.915079874312403e-12
+   -1.048891667810663e-11
+    8.388197205325173e-11
+     -9.5242453460939e-13
+   -1.911141244685034e-12
+   -2.142831558547343e-11
+    8.102137086611358e-11
+ 5.04e+10    
+    8.114366437954995e-11
+   -2.143129447385327e-11
+    8.385936389736737e-11
+   -1.916525360429444e-12
+   -1.049276411024807e-11
+    8.388149729917889e-11
+   -9.500933984181304e-13
+   -1.912597263069568e-12
+   -2.143293289686558e-11
+    8.101500374407854e-11
+ 5.05e+10    
+    8.113722857399833e-11
+   -2.143591773503948e-11
+    8.385888472531232e-11
+   -1.917955861611081e-12
+   -1.049662069202095e-11
+    8.388101251843818e-11
+   -9.477425928346375e-13
+   -1.914038369408097e-12
+   -2.143755606330761e-11
+    8.100861253157988e-11
+ 5.06e+10    
+    8.113076846851144e-11
+   -2.144054671983889e-11
+    8.385839543645767e-11
+   -1.919371331085092e-12
+   -1.050048642341979e-11
+    8.388051765501175e-11
+   -9.453721756684252e-13
+   -1.915464516838379e-12
+   -2.144218501282307e-11
+    8.100219719360763e-11
+ 5.07e+10    
+    8.112428402796582e-11
+   -2.144518135567863e-11
+    8.385789597426823e-11
+   -1.920771722358931e-12
+   -1.050436130451946e-11
+    8.388001265295935e-11
+   -9.429822053085563e-13
+   -1.916875658775819e-12
+    -2.14468196732209e-11
+    8.099575769539509e-11
+ 5.08e+10    
+    8.111777521748317e-11
+   -2.144982156977332e-11
+    8.385738628229053e-11
+   -1.922156989222082e-12
+   -1.050824533547343e-11
+    8.387949745641877e-11
+   -9.405727407252673e-13
+   -1.918271748915829e-12
+   -2.145145997209624e-11
+    8.098929400241762e-11
+ 5.09e+10    
+     8.11112420024294e-11
+    -2.14544672891256e-11
+    8.385686630415351e-11
+   -1.923527085748525e-12
+   -1.051213851651198e-11
+    8.387897200960583e-11
+     -9.3814384147148e-13
+   -1.919652741236279e-12
+   -2.145610583683126e-11
+    8.098280608039104e-11
+ 5.1e+10     
+    8.110468434841304e-11
+   -2.145911844052721e-11
+    8.385633598356819e-11
+   -1.924881966299062e-12
+   -1.051604084794041e-11
+     8.38784362568144e-11
+   -9.356955676843117e-13
+   -1.921018589999796e-12
+    -2.14607571945959e-11
+    8.097629389527001e-11
+ 5.11e+10    
+    8.109810222128329e-11
+   -2.146377495055954e-11
+    8.385579526432799e-11
+   -1.926221585523716e-12
+   -1.051995233013717e-11
+     8.38778901424167e-11
+   -9.332279800864904e-13
+   -1.922369249756173e-12
+   -2.146541397234869e-11
+    8.096975741324667e-11
+ 5.12e+10    
+    8.109149558712925e-11
+   -2.146843674559458e-11
+    8.385524409030895e-11
+   -1.927545898364014e-12
+    -1.05238729635522e-11
+    8.387733361086308e-11
+   -9.307411399877665e-13
+   -1.923704675344614e-12
+   -2.147007609683742e-11
+    8.096319660074843e-11
+ 5.13e+10    
+    8.108486441227759e-11
+   -2.147310375179563e-11
+    8.385468240546964e-11
+    -1.92885486005531e-12
+   -1.052780274870495e-11
+    8.387676660668244e-11
+   -9.282351092862164e-13
+    -1.92502482189608e-12
+   -2.147474349460013e-11
+    8.095661142443745e-11
+ 5.14e+10    
+    8.107820866329156e-11
+   -2.147777589511822e-11
+    8.385411015385144e-11
+    -1.93014842612905e-12
+   -1.053174168618273e-11
+    8.387618907448181e-11
+   -9.257099504695357e-13
+   -1.926329644835529e-12
+   -2.147941609196571e-11
+     8.09500018512082e-11
+ 5.15e+10    
+    8.107152830696963e-11
+   -2.148245310131085e-11
+    8.385352727957874e-11
+    -1.93142655241501e-12
+   -1.053568977663884e-11
+     8.38756009589469e-11
+   -9.231657266162578e-13
+   -1.927619099884155e-12
+   -2.148409381505489e-11
+    8.094336784818659e-11
+ 5.16e+10    
+    8.106482331034348e-11
+   -2.148713529591578e-11
+    8.385293372685854e-11
+   -1.932689195043565e-12
+   -1.053964702079074e-11
+    8.387500220484206e-11
+   -9.206025013969232e-13
+   -1.928893143061604e-12
+   -2.148877658978091e-11
+    8.093670938272794e-11
+ 5.17e+10    
+    8.105809364067707e-11
+   -2.149182240426994e-11
+    8.385232943998105e-11
+   -1.933936310447816e-12
+   -1.054361341941835e-11
+    8.387439275700988e-11
+   -9.180203390751932e-13
+   -1.930151730688164e-12
+    -2.14934643418504e-11
+    8.093002642241617e-11
+ 5.18e+10    
+    8.105133926546472e-11
+   -2.149651435150568e-11
+    8.385171436331969e-11
+   -1.935167855365821e-12
+   -1.054758897336216e-11
+     8.38737725603719e-11
+   -9.154193045088874e-13
+   -1.931394819386941e-12
+    -2.14981569967642e-11
+    8.092331893506136e-11
+ 5.19e+10    
+    8.104456015243027e-11
+   -2.150121106255175e-11
+    8.385108844133103e-11
+   -1.936383786842715e-12
+   -1.055157368352151e-11
+    8.387314155992835e-11
+    -9.12799463151021e-13
+   -1.932622366085949e-12
+   -2.150285447981828e-11
+    8.091658688869953e-11
+ 5.2e+10     
+    8.103775626952524e-11
+   -2.150591246213403e-11
+    8.385045161855503e-11
+   -1.937584062232829e-12
+   -1.055556755085274e-11
+    8.387249970075816e-11
+   -9.101608810507017e-13
+   -1.933834328020289e-12
+   -2.150755671610438e-11
+    8.090983025158992e-11
+ 5.21e+10    
+    8.103092758492742e-11
+   -2.151061847477631e-11
+    8.384980383961463e-11
+   -1.938768639201817e-12
+    -1.05595705763674e-11
+    8.387184692801907e-11
+   -9.075036248540426e-13
+   -1.935030662734191e-12
+   -2.151226363051106e-11
+    8.090304899221449e-11
+ 5.22e+10    
+    8.102407406703949e-11
+   -2.151532902480142e-11
+    8.384914504921676e-11
+   -1.939937475728673e-12
+   -1.056358276113053e-11
+    8.387118318694765e-11
+   -9.048277618049731e-13
+   -1.936211328083094e-12
+   -2.151697514772448e-11
+    8.089624307927612e-11
+ 5.23e+10    
+    8.101719568448781e-11
+    -2.15200440363318e-11
+    8.384847519215153e-11
+    -1.94109053010782e-12
+    -1.05676041062588e-11
+    8.387050842285952e-11
+   -9.021333597460091e-13
+   -1.937376282235658e-12
+   -2.152169119222925e-11
+    8.088941248169702e-11
+ 5.24e+10    
+    8.101029240612087e-11
+   -2.152476343329055e-11
+    8.384779421329255e-11
+   -1.942227760951135e-12
+   -1.057163461291869e-11
+    8.386982258114894e-11
+   -8.994204871189489e-13
+   -1.938525483675824e-12
+   -2.152641168830926e-11
+     8.08825571686177e-11
+ 5.25e+10    
+    8.100336420100796e-11
+   -2.152948713940231e-11
+    8.384710205759717e-11
+   -1.943349127189896e-12
+   -1.057567428232486e-11
+    8.386912560728947e-11
+   -8.966892129655314e-13
+   -1.939658891204757e-12
+   -2.153113656004874e-11
+    8.087567710939548e-11
+ 5.26e+10    
+    8.099641103843762e-11
+   -2.153421507819397e-11
+    8.384639867010623e-11
+   -1.944454588076799e-12
+   -1.057972311573825e-11
+     8.38684174468336e-11
+   -8.939396069280114e-13
+   -1.940776463942809e-12
+   -2.153586573133293e-11
+     8.08687722736027e-11
+ 5.27e+10    
+    8.098943288791674e-11
+   -2.153894717299588e-11
+    8.384568399594457e-11
+   -1.945544103187875e-12
+   -1.058378111446429e-11
+    8.386769804541261e-11
+   -8.911717392496764e-13
+   -1.941878161331491e-12
+   -2.154059912584906e-11
+    8.086184263102597e-11
+ 5.28e+10    
+     8.09824297191688e-11
+   -2.154368334694246e-11
+    8.384495798032019e-11
+   -1.946617632424446e-12
+   -1.058784827985116e-11
+    8.386696734873713e-11
+   -8.883856807753138e-13
+    -1.94296394313536e-12
+   -2.154533666708735e-11
+    8.085488815166441e-11
+ 5.29e+10    
+    8.097540150213256e-11
+   -2.154842352297328e-11
+    8.384422056852551e-11
+   -1.947675136014943e-12
+   -1.059192461328814e-11
+     8.38662253025968e-11
+   -8.855815029516076e-13
+   -1.944033769443894e-12
+   -2.155007827834171e-11
+    8.084790880572817e-11
+ 5.3e+10     
+    8.096834820696104e-11
+   -2.155316762383394e-11
+    8.384347170593629e-11
+   -1.948716574516871e-12
+   -1.059601011620358e-11
+    8.386547185286048e-11
+   -8.827592778274738e-13
+   -1.945087600673369e-12
+   -2.155482388271098e-11
+    8.084090456363777e-11
+ 5.31e+10    
+    8.096126980401961e-11
+   -2.155791557207687e-11
+    8.384271133801194e-11
+   -1.949741908818577e-12
+   -1.060010479006333e-11
+    8.386470694547588e-11
+   -8.799190780543267e-13
+   -1.946125397568707e-12
+   -2.155957340309941e-11
+    8.083387539602178e-11
+ 5.32e+10    
+     8.09541662638856e-11
+   -2.156266729006262e-11
+    8.384193941029632e-11
+   -1.950751100141114e-12
+     -1.0604208636369e-11
+    8.386393052647014e-11
+   -8.770609768862858e-13
+    -1.94714712120526e-12
+   -2.156432676221809e-11
+    8.082682127371629e-11
+ 5.33e+10    
+    8.094703755734587e-11
+   -2.156742269996032e-11
+    8.384115586841653e-11
+    -1.95174411004001e-12
+   -1.060832165665607e-11
+     8.38631425419496e-11
+    -8.74185048180318e-13
+   -1.948152732990619e-12
+   -2.156908388258555e-11
+    8.081974216776315e-11
+ 5.34e+10    
+    8.093988365539656e-11
+    -2.15721817237491e-11
+    8.384036065808378e-11
+    -1.95272090040705e-12
+   -1.061244385249223e-11
+    8.386234293809949e-11
+   -8.712913663963268e-13
+    -1.94914219466636e-12
+   -2.157384468652882e-11
+    8.081263804940895e-11
+ 5.35e+10    
+    8.093270452924107e-11
+   -2.157694428321868e-11
+    8.383955372509295e-11
+   -1.953681433472017e-12
+   -1.061657522547557e-11
+    8.386153166118457e-11
+   -8.683800065971484e-13
+   -1.950115468309809e-12
+   -2.157860909618444e-11
+    8.080550889010347e-11
+ 5.36e+10    
+    8.092550015028911e-11
+   -2.158171029997064e-11
+    8.383873501532322e-11
+   -1.954625671804397e-12
+   -1.062071577723296e-11
+    8.386070865754871e-11
+   -8.654510444485067e-13
+   -1.951072516335722e-12
+   -2.158337703349939e-11
+    8.079835466149851e-11
+ 5.37e+10    
+     8.09182704901554e-11
+   -2.158647969541918e-11
+    8.383790447473723e-11
+   -1.955553578315107e-12
+   -1.062486550941817e-11
+    8.385987387361493e-11
+   -8.625045562188929e-13
+   -1.952013301497993e-12
+   -2.158814842023211e-11
+    8.079117533544655e-11
+ 5.38e+10    
+    8.091101552065832e-11
+   -2.159125239079216e-11
+    8.383706204938135e-11
+   -1.956465116258148e-12
+   -1.062902442371018e-11
+    8.385902725588562e-11
+   -8.595406187793775e-13
+    -1.95293778689131e-12
+   -2.159292317795339e-11
+    8.078397088399957e-11
+ 5.39e+10    
+     8.09037352138187e-11
+   -2.159602830713222e-11
+     8.38362076853862e-11
+   -1.957360249232225e-12
+    -1.06331925218115e-11
+    8.385816875094233e-11
+   -8.565593096033615e-13
+   -1.953845935952794e-12
+   -2.159770122804756e-11
+    8.077674127940785e-11
+ 5.4e+10     
+    8.089642954185852e-11
+   -2.160080736529767e-11
+    8.383534132896608e-11
+   -1.958238941182408e-12
+   -1.063736980544638e-11
+    8.385729830544581e-11
+   -8.535607067662486e-13
+   -1.954737712463649e-12
+   -2.160248249171326e-11
+     8.07694864941183e-11
+ 5.41e+10    
+    8.088909847719982e-11
+   -2.160558948596352e-11
+    8.383446292641911e-11
+   -1.959101156401707e-12
+   -1.064155627635912e-11
+    8.385641586613614e-11
+   -8.505448889450743e-13
+   -1.955613080550685e-12
+   -2.160726688996473e-11
+    8.076220650077374e-11
+ 5.42e+10    
+    8.088174199246342e-11
+   -2.161037458962252e-11
+    8.383357242412705e-11
+   -1.959946859532667e-12
+    -1.06457519363124e-11
+    8.385552137983269e-11
+   -8.475119354180241e-13
+   -1.956472004687941e-12
+   -2.161205434363264e-11
+    8.075490127221131e-11
+ 5.43e+10    
+     8.08743600604673e-11
+   -2.161516259658621e-11
+    8.383266976855572e-11
+   -1.960776015568858e-12
+   -1.064995678708545e-11
+    8.385461479343374e-11
+   -8.444619260639383e-13
+   -1.957314449698214e-12
+   -2.161684477336508e-11
+    8.074757078146129e-11
+ 5.44e+10    
+    8.086695265422628e-11
+   -2.161995342698601e-11
+    8.383175490625456e-11
+   -1.961588589856487e-12
+   -1.065417083047247e-11
+    8.385369605391744e-11
+    -8.41394941361697e-13
+   -1.958140380754574e-12
+   -2.162163809962903e-11
+    8.074021500174624e-11
+ 5.45e+10    
+    8.085951974694968e-11
+   -2.162474700077416e-11
+    8.383082778385694e-11
+   -1.962384548095812e-12
+   -1.065839406828093e-11
+    8.385276510834055e-11
+   -8.383110623895644e-13
+   -1.958949763381851e-12
+   -2.162643424271081e-11
+    8.073283390647896e-11
+ 5.46e+10    
+    8.085206131204098e-11
+   -2.162954323772488e-11
+    8.382988834807987e-11
+   -1.963163856342673e-12
+   -1.066262650232974e-11
+    8.385182190383948e-11
+   -8.352103708244676e-13
+   -1.959742563458134e-12
+   -2.163123312271762e-11
+    8.072542746926216e-11
+ 5.47e+10    
+    8.084457732309633e-11
+   -2.163434205743539e-11
+    8.382893654572396e-11
+   -1.963926481009923e-12
+   -1.066686813444772e-11
+    8.385086638762963e-11
+   -8.320929489411951e-13
+   -1.960518747216178e-12
+   -2.163603465957845e-11
+    8.071799566388676e-11
+ 5.48e+10    
+    8.083706775390328e-11
+   -2.163914337932707e-11
+    8.382797232367351e-11
+   -1.964672388868864e-12
+   -1.067111896647183e-11
+    8.384989850700567e-11
+   -8.289588796115097e-13
+   -1.961278281244861e-12
+   -2.164083877304516e-11
+    8.071053846433088e-11
+ 5.49e+10    
+    8.082953257843969e-11
+   -2.164394712264651e-11
+    8.382699562889659e-11
+   -1.965401547050628e-12
+   -1.067537900024556e-11
+    8.384891820934168e-11
+   -8.258082463032254e-13
+   -1.962021132490583e-12
+   -2.164564538269369e-11
+    8.070305584475863e-11
+ 5.5e+10     
+    8.082197177087248e-11
+   -2.164875320646656e-11
+    8.382600640844483e-11
+   -1.966113923047588e-12
+   -1.067964823761718e-11
+    8.384792544209075e-11
+    -8.22641133079202e-13
+   -1.962747268258605e-12
+   -2.165045440792499e-11
+     8.06955477795187e-11
+ 5.51e+10    
+    8.081438530555662e-11
+   -2.165356154968756e-11
+    8.382500460945341e-11
+   -1.966809484714709e-12
+   -1.068392668043816e-11
+    8.384692015278506e-11
+   -8.194576245962368e-13
+   -1.963456656214477e-12
+   -2.165526576796627e-11
+    8.068801424314348e-11
+ 5.52e+10    
+    8.080677315703386e-11
+   -2.165837207103844e-11
+    8.382399017914115e-11
+   -1.967488200270851e-12
+    -1.06882143305615e-11
+    8.384590228903627e-11
+   -8.162578061039507e-13
+   -1.964149264385267e-12
+   -2.166007938187217e-11
+    8.068045521034777e-11
+ 5.53e+10    
+    8.079913530003138e-11
+   -2.166318468907776e-11
+    8.382296306481026e-11
+   -1.968150038300116e-12
+   -1.069251118984003e-11
+    8.384487179853502e-11
+   -8.130417634435397e-13
+   -1.964825061160964e-12
+   -2.166489516852585e-11
+    8.067287065602779e-11
+ 5.54e+10    
+    8.079147170946114e-11
+   -2.166799932219499e-11
+    8.382192321384649e-11
+   -1.968794967753112e-12
+   -1.069681726012482e-11
+    8.384382862905105e-11
+   -8.098095830464936e-13
+   -1.965484015295706e-12
+   -2.166971304664006e-11
+    8.066526055525974e-11
+ 5.55e+10    
+    8.078378236041825e-11
+   -2.167281588861161e-11
+     8.38208705737189e-11
+   -1.969422957948228e-12
+   -1.070113254326353e-11
+    8.384277272843367e-11
+   -8.065613519332179e-13
+   -1.966126095909054e-12
+   -2.167453293475854e-11
+    8.065762488329888e-11
+ 5.56e+10    
+     8.07760672281798e-11
+   -2.167763430638223e-11
+    8.381980509198023e-11
+   -1.970033978572863e-12
+    -1.07054570410988e-11
+    8.384170404461076e-11
+   -8.032971577116174e-13
+    -1.96675127248724e-12
+   -2.167935475125695e-11
+    8.064996361557818e-11
+ 5.57e+10    
+    8.076832628820445e-11
+   -2.168245449339592e-11
+    8.381872671626628e-11
+   -1.970627999684648e-12
+   -1.070979075546659e-11
+    8.384062252558967e-11
+    -8.00017088575581e-13
+   -1.967359514884362e-12
+   -2.168417841434414e-11
+     8.06422767277075e-11
+ 5.58e+10    
+    8.076055951613032e-11
+   -2.168727636737723e-11
+    8.381763539429628e-11
+   -1.971204991712637e-12
+   -1.071413368819464e-11
+     8.38395281194568e-11
+   -7.967212333033945e-13
+   -1.967950793323595e-12
+   -2.168900384206348e-11
+    8.063456419547217e-11
+ 5.59e+10    
+    8.075276688777476e-11
+   -2.169209984588755e-11
+    8.381653107387276e-11
+   -1.971764925458481e-12
+   -1.071848584110074e-11
+     8.38384207743775e-11
+   -7.934096812560996e-13
+   -1.968525078398353e-12
+   -2.169383095229385e-11
+    8.062682599483197e-11
+ 5.6e+10     
+    8.074494837913245e-11
+   -2.169692484632615e-11
+    8.381541370288148e-11
+   -1.972307772097591e-12
+   -1.072284721599132e-11
+    8.383730043859672e-11
+   -7.900825223757681e-13
+   -1.969082341073439e-12
+   -2.169865966275115e-11
+    8.061906210192024e-11
+ 5.61e+10    
+    8.073710396637498e-11
+    -2.17017512859316e-11
+    8.381428322929119e-11
+    -1.97283350318022e-12
+   -1.072721781465964e-11
+     8.38361670604377e-11
+    -7.86739847183706e-13
+   -1.969622552686164e-12
+   -2.170348989098913e-11
+    8.061127249304238e-11
+ 5.62e+10    
+    8.072923362584917e-11
+   -2.170657908178285e-11
+    8.381313960115403e-11
+   -1.973342090632609e-12
+   -1.073159763888442e-11
+    8.383502058830341e-11
+   -7.833817467785861e-13
+   -1.970145684947449e-12
+   -2.170832155440108e-11
+    8.060345714467502e-11
+ 5.63e+10    
+    8.072133733407662e-11
+   -2.171140815080065e-11
+    8.381198276660532e-11
+    -1.97383350675804e-12
+    -1.07359866904281e-11
+    8.383386097067553e-11
+   -7.800083128345194e-13
+   -1.970651709942924e-12
+   -2.171315457022074e-11
+    8.059561603346495e-11
+ 5.64e+10    
+    8.071341506775192e-11
+   -2.171623840974852e-11
+    8.381081267386301e-11
+   -1.974307724237927e-12
+   -1.074038497103539e-11
+    8.383268815611492e-11
+   -7.766196375990243e-13
+   -1.971140600133951e-12
+   -2.171798885552376e-11
+    8.058774913622771e-11
+ 5.65e+10    
+    8.070546680374211e-11
+   -2.172106977523437e-11
+    8.380962927122843e-11
+    -1.97476471613281e-12
+   -1.074479248243161e-11
+    8.383150209326138e-11
+   -7.732158138909589e-13
+   -1.971612328358703e-12
+   -2.172282432722891e-11
+    8.057985642994707e-11
+ 5.66e+10    
+    8.069749251908524e-11
+    -2.17259021637115e-11
+    8.380843250708575e-11
+   -1.975204455883387e-12
+   -1.074920922632124e-11
+    8.383030273083381e-11
+   -7.697969350983587e-13
+   -1.972066867833138e-12
+   -2.172766090209941e-11
+    8.057193789177349e-11
+ 5.67e+10    
+    8.068949219098968e-11
+   -2.173073549148014e-11
+    8.380722232990229e-11
+   -1.975626917311519e-12
+   -1.075363520438635e-11
+    8.382909001763021e-11
+   -7.663630951762094e-13
+   -1.972504192152017e-12
+    -2.17324984967442e-11
+    8.056399349902333e-11
+ 5.68e+10    
+    8.068146579683265e-11
+   -2.173556967468849e-11
+    8.380599868822781e-11
+   -1.976032074621175e-12
+   -1.075807041828497e-11
+    8.382786390252723e-11
+    -7.62914388644155e-13
+   -1.972924275289871e-12
+   -2.173733702761923e-11
+    8.055602322917751e-11
+ 5.69e+10    
+    8.067341331415958e-11
+   -2.174040462933426e-11
+    8.380476153069529e-11
+   -1.976419902399403e-12
+   -1.076251486964971e-11
+    8.382662433448082e-11
+   -7.594509105841022e-13
+   -1.973327091601941e-12
+   -2.174217641102883e-11
+    8.054802705988083e-11
+ 5.7e+10     
+     8.06653347206827e-11
+   -2.174524027126589e-11
+    8.380351080602032e-11
+   -1.976790375617228e-12
+   -1.076696856008614e-11
+    8.382537126252588e-11
+   -7.559727566378094e-13
+   -1.973712615825104e-12
+     -2.1747016563127e-11
+    8.054000496894049e-11
+ 5.71e+10    
+    8.065722999428008e-11
+   -2.175007651618387e-11
+    8.380224646300136e-11
+   -1.977143469630596e-12
+   -1.077143149117138e-11
+    8.382410463577623e-11
+   -7.524800230043308e-13
+   -1.974080823078808e-12
+   -2.175185739991893e-11
+    8.053195693432573e-11
+ 5.72e+10    
+    8.064909911299493e-11
+   -2.175491327964226e-11
+     8.38009684505196e-11
+    -1.97747916018121e-12
+   -1.077590366445246e-11
+     8.38228244034246e-11
+   -7.489728064374623e-13
+   -1.974431688865911e-12
+   -2.175669883726203e-11
+    8.052388293416571e-11
+ 5.73e+10    
+    8.064094205503399e-11
+   -2.175975047704978e-11
+    8.379967671753893e-11
+   -1.977797423397428e-12
+   -1.078038508144499e-11
+    8.382153051474279e-11
+   -7.454512042430614e-13
+   -1.974765189073598e-12
+   -2.176154079086765e-11
+    8.051578294674991e-11
+ 5.74e+10    
+    8.063275879876705e-11
+   -2.176458802367146e-11
+    8.379837121310573e-11
+   -1.978098235795091e-12
+   -1.078487574363154e-11
+    8.382022291908157e-11
+   -7.419153142763101e-13
+   -1.975081299974171e-12
+    -2.17663831763022e-11
+    8.050765695052575e-11
+ 5.75e+10    
+    8.062454932272559e-11
+   -2.176942583462978e-11
+    8.379705188634913e-11
+   -1.978381574278341e-12
+   -1.078937565246024e-11
+    8.381890156587044e-11
+   -7.383652349389308e-13
+   -1.975379998225913e-12
+   -2.177122590898869e-11
+    8.049950492409846e-11
+ 5.76e+10    
+    8.061631360560188e-11
+    -2.17742638249063e-11
+    8.379571868648088e-11
+    -1.97864741614041e-12
+   -1.079388480934333e-11
+    8.381756640461817e-11
+   -7.348010651762825e-13
+    -1.97566126087387e-12
+   -2.177606890420818e-11
+    8.049132684622986e-11
+ 5.77e+10    
+     8.06080516262481e-11
+   -2.177910190934293e-11
+    8.379437156279513e-11
+    -1.97889573906441e-12
+   -1.079840321565565e-11
+    8.381621738491223e-11
+   -7.312229044744343e-13
+    -1.97592506535062e-12
+   -2.178091207710096e-11
+    8.048312269583701e-11
+ 5.78e+10    
+    8.059976336367502e-11
+   -2.178394000264331e-11
+    8.379301046466856e-11
+   -1.979126521124097e-12
+   -1.080293087273326e-11
+    8.381485445641932e-11
+   -7.276308528571354e-13
+   -1.976171389477072e-12
+   -2.178575534266828e-11
+    8.047489245199188e-11
+ 5.79e+10    
+    8.059144879705123e-11
+   -2.178877801937444e-11
+    8.379163534156056e-11
+   -1.979339740784575e-12
+   -1.080746778187194e-11
+    8.381347756888478e-11
+    -7.24025010882715e-13
+   -1.976400211463172e-12
+   -2.179059861577358e-11
+    8.046663609391971e-11
+ 5.8e+10     
+    8.058310790570231e-11
+   -2.179361587396792e-11
+    8.379024614301278e-11
+   -1.979535376903046e-12
+    -1.08120139443258e-11
+     8.38120866721332e-11
+   -7.204054796409404e-13
+   -1.976611509908624e-12
+   -2.179544181114405e-11
+    8.045835360099846e-11
+ 5.81e+10    
+    8.057474066910961e-11
+    -2.17984534807215e-11
+    8.378884281864905e-11
+   -1.979713408729492e-12
+   -1.081656936130582e-11
+     8.38106817160679e-11
+   -7.167723607497687e-13
+   -1.976805263803608e-12
+   -2.180028484337207e-11
+    8.045004495275783e-11
+ 5.82e+10    
+    8.056634706690903e-11
+   -2.180329075380055e-11
+    8.378742531817609e-11
+   -1.979873815907325e-12
+   -1.082113403397857e-11
+    8.380926265067128e-11
+   -7.131257563520415e-13
+   -1.976981452529457e-12
+   -2.180512762691656e-11
+    8.044171012887776e-11
+ 5.83e+10    
+    8.055792707889098e-11
+   -2.180812760723963e-11
+    8.378599359138275e-11
+   -1.980016578474087e-12
+   -1.082570796346464e-11
+    8.380782942600477e-11
+   -7.094657691121189e-13
+   -1.977140055859288e-12
+   -2.180997007610474e-11
+    8.043334910918829e-11
+ 5.84e+10    
+    8.054948068499813e-11
+   -2.181296395494369e-11
+    8.378454758814013e-11
+   -1.980141676862048e-12
+   -1.083029115083736e-11
+    8.380638199220876e-11
+   -7.057925022124193e-13
+   -1.977281053958686e-12
+   -2.181481210513346e-11
+    8.042496187366821e-11
+ 5.85e+10    
+    8.054100786532551e-11
+   -2.181779971068992e-11
+    8.378308725840189e-11
+   -1.980249091898818e-12
+   -1.083488359712139e-11
+    8.380492029950255e-11
+   -7.021060593499296e-13
+   -1.977404427386281e-12
+   -2.181965362807062e-11
+    8.041654840244373e-11
+ 5.86e+10    
+    8.053250860011909e-11
+   -2.182263478812905e-11
+    8.378161255220376e-11
+   -1.980338804807976e-12
+   -1.083948530329133e-11
+    8.380344429818461e-11
+   -6.984065447325895e-13
+   -1.977510157094372e-12
+   -2.182449455885685e-11
+    8.040810867578826e-11
+ 5.87e+10    
+    8.052398286977494e-11
+   -2.182746910078698e-11
+    8.378012341966384e-11
+   -1.980410797209623e-12
+   -1.084409627027044e-11
+    8.380195393863248e-11
+    -6.94694063075649e-13
+   -1.977598224429506e-12
+   -2.182933481130708e-11
+    8.039964267412097e-11
+ 5.88e+10    
+    8.051543065483817e-11
+   -2.183230256206629e-11
+     8.37786198109827e-11
+   -1.980465051120904e-12
+   -1.084871649892921e-11
+    8.380044917130253e-11
+   -6.909687195979534e-13
+   -1.977668611133047e-12
+   -2.183417429911194e-11
+    8.039115037800634e-11
+ 5.89e+10    
+    8.050685193600223e-11
+   -2.183713508524771e-11
+    8.377710167644288e-11
+   -1.980501548956608e-12
+   -1.085334599008402e-11
+    8.379892994673046e-11
+   -6.872306200181351e-13
+   -1.977721299341677e-12
+   -2.183901293583938e-11
+    8.038263176815254e-11
+ 5.9e+10     
+    8.049824669410788e-11
+   -2.184196658349187e-11
+    8.377556896640948e-11
+   -1.980520273529628e-12
+    -1.08579847444959e-11
+    8.379739621553088e-11
+   -6.834798705507557e-13
+   -1.977756271587977e-12
+   -2.184385063493628e-11
+    8.037408682541114e-11
+ 5.91e+10    
+    8.048961491014195e-11
+   -2.184679696984065e-11
+    8.377402163132956e-11
+   -1.980521208051487e-12
+   -1.086263276286909e-11
+    8.379584792839762e-11
+   -6.797165779023773e-13
+   -1.977773510800898e-12
+   -2.184868730972994e-11
+    8.036551553077584e-11
+ 5.92e+10    
+    8.048095656523734e-11
+   -2.185162615721903e-11
+    8.377245962173241e-11
+   -1.980504336132806e-12
+    -1.08672900458498e-11
+    8.379428503610373e-11
+    -6.75940849267566e-13
+   -1.977773000306228e-12
+    -2.18535228734298e-11
+      8.0356917865382e-11
+ 5.93e+10    
+    8.047227164067088e-11
+   -2.185645405843636e-11
+    8.377088288822989e-11
+   -1.980469641783761e-12
+   -1.087195659402492e-11
+    8.379270748950113e-11
+   -6.721527923248169e-13
+   -1.977754723827121e-12
+    -2.18583572391289e-11
+    8.034829381050522e-11
+ 5.94e+10    
+    8.046356011786348e-11
+   -2.186128058618832e-11
+    8.376929138151582e-11
+   -1.980417109414526e-12
+   -1.087663240792074e-11
+    8.379111523952167e-11
+   -6.683525152324223e-13
+   -1.977718665484457e-12
+   -2.186319031980573e-11
+    8.033964334756075e-11
+ 5.95e+10    
+    8.045482197837866e-11
+   -2.186610565305826e-11
+    8.376768505236648e-11
+   -1.980346723835684e-12
+    -1.08813174880016e-11
+    8.378950823717554e-11
+   -6.645401266242738e-13
+    -1.97766480979736e-12
+   -2.186802202832548e-11
+    8.033096645810266e-11
+ 5.96e+10    
+    8.044605720392186e-11
+   -2.187092917151897e-11
+    8.376606385164021e-11
+   -1.980258470258637e-12
+   -1.088601183466869e-11
+    8.378788643355286e-11
+   -6.607157356055955e-13
+   -1.977593141683542e-12
+   -2.187285227744212e-11
+    8.032226312382282e-11
+ 5.97e+10    
+    8.043726577633961e-11
+   -2.187575105393433e-11
+    8.376442773027748e-11
+   -1.980152334295991e-12
+   -1.089071544825875e-11
+    8.378624977982288e-11
+   -6.568794517486071e-13
+   -1.977503646459733e-12
+   -2.187768097979967e-11
+    8.031353332655022e-11
+ 5.98e+10    
+    8.042844767761837e-11
+   -2.188057121256086e-11
+    8.376277663930135e-11
+   -1.980028301961911e-12
+   -1.089542832904288e-11
+    8.378459822723418e-11
+   -6.530313850881149e-13
+   -1.977396309842017e-12
+   -2.188250804793411e-11
+    8.030477704824974e-11
+ 5.99e+10    
+    8.041960288988439e-11
+   -2.188538955954962e-11
+    8.376111052981708e-11
+   -1.979886359672478e-12
+   -1.090015047722524e-11
+    8.378293172711482e-11
+   -6.491716461170658e-13
+   -1.977271117946242e-12
+   -2.188733339427494e-11
+    8.029599427102177e-11
+ 6e+10       
+    8.041073139540161e-11
+   -2.189020600694757e-11
+    8.375942935301216e-11
+   -1.979726494245987e-12
+   -1.090488189294189e-11
+    8.378125023087241e-11
+   -6.453003457819977e-13
+   -1.977128057288314e-12
+   -2.189215693114695e-11
+    8.028718497710108e-11
+ 6.01e+10    
+    8.040183317657222e-11
+   -2.189502046669947e-11
+    8.375773306015624e-11
+    -1.97954869290331e-12
+   -1.090962257625949e-11
+    8.377955368999385e-11
+   -6.414175954784574e-13
+   -1.976967114784524e-12
+   -2.189697857077174e-11
+      8.0278349148856e-11
+ 6.02e+10    
+    8.039290821593472e-11
+   -2.189983285064954e-11
+    8.375602160260146e-11
+   -1.979352943268139e-12
+   -1.091437252717416e-11
+    8.377784205604571e-11
+   -6.375235070463339e-13
+   -1.976788277751863e-12
+   -2.190179822526965e-11
+    8.026948676878775e-11
+ 6.03e+10    
+     8.03839564961639e-11
+   -2.190464307054325e-11
+    8.375429493178271e-11
+   -1.979139233367284e-12
+   -1.091913174561032e-11
+    8.377611528067447e-11
+   -6.336181927651349e-13
+   -1.976591533908301e-12
+   -2.190661580666141e-11
+    8.026059781952955e-11
+ 6.04e+10    
+    8.037497800006918e-11
+    -2.19094510380288e-11
+    8.375255299921648e-11
+   -1.978907551630914e-12
+   -1.092390023141937e-11
+    8.377437331560571e-11
+   -6.297017653492105e-13
+   -1.976376871373051e-12
+   -2.191143122686973e-11
+    8.025168228384572e-11
+ 6.05e+10    
+    8.036597271059458e-11
+   -2.191425666465914e-11
+    8.375079575650225e-11
+   -1.978657886892803e-12
+   -1.092867798437865e-11
+    8.377261611264527e-11
+   -6.257743379428946e-13
+   -1.976144278666831e-12
+   -2.191624439772117e-11
+    8.024274014463084e-11
+ 6.06e+10    
+     8.03569406108174e-11
+   -2.191905986189351e-11
+    8.374902315532189e-11
+   -1.978390228390567e-12
+    -1.09334650041903e-11
+    8.377084362367869e-11
+   -6.218360241155913e-13
+   -1.975893744712048e-12
+   -2.192105523094798e-11
+    8.023377138490915e-11
+ 6.07e+10    
+    8.034788168394766e-11
+   -2.192386054109944e-11
+    8.374723514743976e-11
+   -1.978104565765823e-12
+   -1.093826129047993e-11
+    8.376905580067116e-11
+   -6.178869378568184e-13
+   -1.975625258833106e-12
+   -2.192586363818961e-11
+    8.022477598783381e-11
+ 6.08e+10    
+    8.033879591332712e-11
+   -2.192865861355414e-11
+    8.374543168470238e-11
+   -1.977800889064425e-12
+   -1.094306684279566e-11
+    8.376725259566814e-11
+   -6.139271935711566e-13
+   -1.975338810756496e-12
+   -2.193066953099471e-11
+    8.021575393668557e-11
+ 6.09e+10    
+    8.032968328242863e-11
+   -2.193345399044661e-11
+    8.374361271903939e-11
+   -1.977479188736593e-12
+   -1.094788166060692e-11
+    8.376543396079483e-11
+   -6.099569060731684e-13
+   -1.975034390611056e-12
+   -2.193547282082275e-11
+    8.020670521487269e-11
+ 6.1e+10     
+    8.032054377485539e-11
+   -2.193824658287935e-11
+    8.374177820246289e-11
+   -1.977139455637089e-12
+   -1.095270574330334e-11
+    8.376359984825675e-11
+   -6.059761905822343e-13
+   -1.974711988928104e-12
+   -2.194027341904605e-11
+     8.01976298059298e-11
+ 6.11e+10    
+    8.031137737433998e-11
+   -2.194303630187007e-11
+     8.37399280870674e-11
+    -1.97678168102534e-12
+   -1.095753909019364e-11
+    8.376175021033951e-11
+   -6.019851627173438e-13
+   -1.974371596641579e-12
+   -2.194507123695123e-11
+    8.018852769351707e-11
+ 6.12e+10    
+    8.030218406474355e-11
+   -2.194782305835352e-11
+    8.373806232503056e-11
+    -1.97640585656555e-12
+   -1.096238170050454e-11
+    8.375988499940899e-11
+   -5.979839384918228e-13
+   -1.974013205088189e-12
+   -2.194986618574139e-11
+    8.017939886141983e-11
+ 6.13e+10    
+    8.029296383005558e-11
+   -2.195260676318349e-11
+    8.373618086861274e-11
+   -1.976011974326813e-12
+    -1.09672335733797e-11
+    8.375800416791144e-11
+   -5.939726343080096e-13
+   -1.973636806007516e-12
+   -2.195465817653768e-11
+    8.017024329354736e-11
+ 6.14e+10    
+    8.028371665439237e-11
+   -2.195738732713443e-11
+    8.373428367015691e-11
+   -1.975600026783191e-12
+   -1.097209470787857e-11
+    8.375610766837353e-11
+   -5.899513669518506e-13
+   -1.973242391542118e-12
+    -2.19594471203813e-11
+    8.016106097393252e-11
+ 6.15e+10    
+    8.027444252199688e-11
+   -2.196216466090332e-11
+    8.373237068208913e-11
+    -1.97517000681378e-12
+   -1.097696510297542e-11
+    8.375419545340244e-11
+   -5.859202535874711e-13
+   -1.972829954237589e-12
+   -2.196423292823511e-11
+    8.015185188673065e-11
+ 6.16e+10    
+     8.02651414172376e-11
+   -2.196693867511161e-11
+    8.373044185691846e-11
+   -1.974721907702757e-12
+   -1.098184475755827e-11
+    8.375226747568613e-11
+   -5.818794117516706e-13
+   -1.972399487042653e-12
+   -2.196901551098591e-11
+    8.014261601621935e-11
+ 6.17e+10    
+    8.025581332460826e-11
+   -2.197170928030714e-11
+     8.37284971472372e-11
+   -1.974255723139423e-12
+   -1.098673367042778e-11
+    8.375032368799314e-11
+   -5.778289593483549e-13
+   -1.971950983309211e-12
+   -2.197379477944591e-11
+    8.013335334679743e-11
+ 6.18e+10    
+     8.02464582287266e-11
+   -2.197647638696574e-11
+     8.37265365057205e-11
+   -1.973771447218219e-12
+   -1.099163184029631e-11
+    8.374836404317302e-11
+   -5.737690146429395e-13
+   -1.971484436792343e-12
+   -2.197857064435475e-11
+    8.012406386298412e-11
+ 6.19e+10    
+    8.023707611433399e-11
+   -2.198123990549346e-11
+    8.372455988512693e-11
+   -1.973269074438715e-12
+   -1.099653926578685e-11
+    8.374638849415587e-11
+   -5.696996962566726e-13
+   -1.970999841650362e-12
+   -2.198334301638131e-11
+    8.011474754941848e-11
+ 6.2e+10     
+    8.022766696629467e-11
+   -2.198599974622822e-11
+    8.372256723829825e-11
+   -1.972748599705619e-12
+   -1.100145594543204e-11
+    8.374439699395342e-11
+   -5.656211231609158e-13
+   -1.970497192444773e-12
+   -2.198811180612592e-11
+    8.010540439085891e-11
+ 6.21e+10    
+    8.021823076959476e-11
+   -2.199075581944178e-11
+    8.372055851815971e-11
+   -1.972210018328719e-12
+   -1.100638187767318e-11
+    8.374238949565815e-11
+   -5.615334146713762e-13
+   -1.969976484140316e-12
+   -2.199287692412181e-11
+     8.00960343721822e-11
+ 6.22e+10    
+    8.020876750934222e-11
+   -2.199550803534175e-11
+    8.371853367772007e-11
+   -1.971653326022852e-12
+   -1.101131706085924e-11
+    8.374036595244393e-11
+   -5.574366904422735e-13
+   -1.969437712104871e-12
+   -2.199763828083736e-11
+    8.008663747838298e-11
+ 6.23e+10    
+    8.019927717076527e-11
+   -2.200025630407333e-11
+    8.371649267007154e-11
+   -1.971078518907851e-12
+   -1.101626149324585e-11
+    8.373832631756607e-11
+   -5.533310704604655e-13
+   -1.968880872109465e-12
+    -2.20023957866779e-11
+    8.007721369457297e-11
+ 6.24e+10    
+    8.018975973921262e-11
+   -2.200500053572143e-11
+     8.37144354483902e-11
+   -1.970485593508454e-12
+   -1.102121517299439e-11
+    8.373627054436144e-11
+    -5.49216675039519e-13
+   -1.968305960328175e-12
+   -2.200714935198764e-11
+    8.006776300598034e-11
+ 6.25e+10    
+    8.018021520015221e-11
+   -2.200974064031252e-11
+     8.37123619659357e-11
+   -1.969874546754204e-12
+   -1.102617809817105e-11
+    8.373419858624859e-11
+   -5.450936248137402e-13
+   -1.967712973338072e-12
+   -2.201189888705172e-11
+     8.00582853979492e-11
+ 6.26e+10    
+    8.017064353917077e-11
+   -2.201447652781661e-11
+    8.371027217605194e-11
+   -1.969245375979354e-12
+    -1.10311502667459e-11
+    8.373211039672775e-11
+   -5.409620407321226e-13
+   -1.967101908119124e-12
+   -2.201664430209797e-11
+    8.004878085593875e-11
+ 6.27e+10    
+    8.016104474197287e-11
+    -2.20192081081491e-11
+    8.370816603216645e-11
+   -1.968598078922739e-12
+   -1.103613167659182e-11
+    8.373000592938092e-11
+   -5.368220440522981e-13
+   -1.966472762054077e-12
+   -2.202138550729906e-11
+    8.003924936552275e-11
+ 6.28e+10    
+     8.01514187943809e-11
+   -2.202393529117296e-11
+    8.370604348779099e-11
+    -1.96793265372764e-12
+   -1.104112232548382e-11
+    8.372788513787262e-11
+   -5.326737563343945e-13
+   -1.965825532928341e-12
+   -2.202612241277442e-11
+    8.002969091238886e-11
+ 6.29e+10    
+    8.014176568233382e-11
+   -2.202865798670053e-11
+    8.370390449652151e-11
+   -1.967249098941624e-12
+   -1.104612221109795e-11
+    8.372574797594925e-11
+   -5.285172994348668e-13
+   -1.965160218929867e-12
+   -2.203085492859222e-11
+    8.002010548233821e-11
+ 6.3e+10     
+    8.013208539188683e-11
+   -2.203337610449573e-11
+    8.370174901203881e-11
+   -1.966547413516358e-12
+   -1.105113133101057e-11
+    8.372359439743963e-11
+   -5.243527955002761e-13
+   -1.964476818648975e-12
+   -2.203558296477129e-11
+    8.001049306128431e-11
+ 6.31e+10    
+    8.012237790921069e-11
+   -2.203808955427568e-11
+    8.369957698810751e-11
+    -1.96582759680747e-12
+   -1.105614968269724e-11
+     8.37214243562551e-11
+   -5.201803669610366e-13
+   -1.963775331078183e-12
+   -2.204030643128324e-11
+    8.000085363525309e-11
+ 6.32e+10    
+     8.01126432205912e-11
+   -2.204279824571314e-11
+    8.369738837857712e-11
+   -1.965089648574301e-12
+   -1.106117726353215e-11
+    8.371923780638978e-11
+   -5.160001365250919e-13
+   -1.963055755612045e-12
+   -2.204502523805445e-11
+    7.999118719038185e-11
+ 6.33e+10    
+    8.010288131242827e-11
+   -2.204750208843818e-11
+    8.369518313738203e-11
+   -1.964333568979714e-12
+     -1.1066214070787e-11
+    8.371703470192016e-11
+   -5.118122271715703e-13
+   -1.962318092046954e-12
+   -2.204973929496787e-11
+    7.998149371291867e-11
+ 6.34e+10    
+    8.009309217123587e-11
+   -2.205220099204052e-11
+    8.369296121854136e-11
+    -1.96355935858986e-12
+   -1.107126010163031e-11
+    8.371481499700626e-11
+   -5.076167621443843e-13
+   -1.961562340580911e-12
+   -2.205444851186548e-11
+    7.997177318922227e-11
+ 6.35e+10    
+    8.008327578364084e-11
+   -2.205689486607123e-11
+    8.369072257615932e-11
+   -1.962767018373948e-12
+   -1.107631535312652e-11
+    8.371257864589084e-11
+   -5.034138649457835e-13
+   -1.960788501813316e-12
+   -2.205915279854988e-11
+    7.996202560576083e-11
+ 6.36e+10    
+    8.007343213638301e-11
+   -2.206158362004511e-11
+    8.368846716442531e-11
+   -1.961956549703951e-12
+    -1.10813798222352e-11
+    8.371032560290021e-11
+   -4.992036593298977e-13
+   -1.959996576744722e-12
+   -2.206385206478668e-11
+      7.9952250949112e-11
+ 6.37e+10    
+    8.006356121631374e-11
+   -2.206626716344237e-11
+    8.368619493761409e-11
+   -1.961127954354375e-12
+   -1.108645350581025e-11
+    8.370805582244389e-11
+   -4.949862692961841e-13
+   -1.959186566776592e-12
+   -2.206854622030624e-11
+    7.994244920596198e-11
+ 6.38e+10    
+    8.005366301039632e-11
+   -2.207094540571112e-11
+    8.368390585008585e-11
+    -1.96028123450194e-12
+    -1.10915364005991e-11
+    8.370576925901546e-11
+   -4.907618190828913e-13
+   -1.958358473711013e-12
+   -2.207323517480608e-11
+    7.993262036310507e-11
+ 6.39e+10    
+    8.004373750570462e-11
+   -2.207561825626903e-11
+    8.368159985628644e-11
+   -1.959416392725303e-12
+   -1.109662850324185e-11
+    8.370346586719197e-11
+   -4.865304331604385e-13
+   -1.957512299750419e-12
+   -2.207791883795261e-11
+    7.992276440744331e-11
+ 6.4e+10     
+    8.003378468942312e-11
+    -2.20802856245057e-11
+     8.36792769107476e-11
+   -1.958533432004719e-12
+   -1.110172981027058e-11
+    8.370114560163434e-11
+   -4.822922362247906e-13
+   -1.956648047497326e-12
+   -2.208259711938337e-11
+    7.991288132598569e-11
+ 6.41e+10    
+    8.002380454884612e-11
+   -2.208494741978459e-11
+    8.367693696808701e-11
+   -1.957632355721735e-12
+    -1.11068403181086e-11
+    8.369880841708837e-11
+   -4.780473531907718e-13
+   -1.955765719953969e-12
+   -2.208726992870924e-11
+    7.990297110584776e-11
+ 6.42e+10    
+    8.001379707137723e-11
+   -2.208960355144517e-11
+    8.367457998300833e-11
+   -1.956713167658814e-12
+   -1.111196002306964e-11
+    8.369645426838358e-11
+   -4.737959091853613e-13
+    -1.95486532052201e-12
+   -2.209193717551621e-11
+     7.98930337342512e-11
+ 6.43e+10    
+    8.000376224452878e-11
+   -2.209425392880501e-11
+    8.367220591030187e-11
+   -1.955775871999021e-12
+   -1.111708892135712e-11
+    8.369408311043427e-11
+   -4.695380295409257e-13
+    -1.95394685300222e-12
+   -2.209659876936775e-11
+    7.988306919852324e-11
+ 6.44e+10    
+    7.999370005592143e-11
+   -2.209889846116183e-11
+    8.366981470484413e-11
+   -1.954820473325606e-12
+   -1.112222700906346e-11
+    8.369169489823969e-11
+   -4.652738397884619e-13
+   -1.953010321594064e-12
+   -2.210125461980688e-11
+    7.987307748609612e-11
+ 6.45e+10    
+     7.99836104932838e-11
+   -2.210353705779568e-11
+    8.366740632159846e-11
+   -1.953846976621646e-12
+   -1.112737428216931e-11
+    8.368928958688389e-11
+   -4.610034656507597e-13
+   -1.952055730895415e-12
+   -2.210590463635811e-11
+    7.986305858450679e-11
+ 6.46e+10    
+    7.997349354445187e-11
+   -2.210816962797117e-11
+    8.366498071561512e-11
+   -1.952855387269656e-12
+   -1.113253073654292e-11
+    8.368686713153622e-11
+   -4.567270330355485e-13
+   -1.951083085902114e-12
+    -2.21105487285298e-11
+    7.985301248139623e-11
+ 6.47e+10    
+    7.996334919736814e-11
+   -2.211279608093931e-11
+     8.36625378420314e-11
+   -1.951845711051132e-12
+   -1.113769636793939e-11
+     8.36844274874511e-11
+   -4.524446680286272e-13
+   -1.950092392007615e-12
+   -2.211518680581604e-11
+    7.984293916450923e-11
+ 6.48e+10    
+     7.99531774400819e-11
+   -2.211741632593989e-11
+    8.366007765607175e-11
+   -1.950817954146178e-12
+   -1.114287117200002e-11
+    8.368197060996925e-11
+   -4.481564968869466e-13
+   -1.949083655002555e-12
+   -2.211981877769911e-11
+    7.983283862169373e-11
+ 6.49e+10    
+    7.994297826074812e-11
+   -2.212203027220355e-11
+    8.365760011304804e-11
+   -1.949772123133018e-12
+   -1.114805514425157e-11
+    8.367949645451651e-11
+   -4.438626460316582e-13
+   -1.948056881074347e-12
+   -2.212444455365124e-11
+    7.982271084090035e-11
+ 6.5e+10     
+     7.99327516476275e-11
+   -2.212663782895393e-11
+    8.365510516836016e-11
+   -1.948708224987584e-12
+   -1.115324828010575e-11
+    8.367700497660513e-11
+   -4.395632420411382e-13
+   -1.947012076806769e-12
+     -2.2129064043137e-11
+    7.981255581018225e-11
+ 6.51e+10    
+    7.992249758908538e-11
+   -2.213123890540971e-11
+    8.365259277749541e-11
+   -1.947626267083024e-12
+   -1.115845057485842e-11
+    8.367449613183361e-11
+   -4.352584116439993e-13
+   -1.945949249179481e-12
+   -2.213367715561549e-11
+    7.980237351769456e-11
+ 6.52e+10    
+    7.991221607359196e-11
+   -2.213583341078703e-11
+    8.365006289602938e-11
+    -1.94652625718923e-12
+   -1.116366202368904e-11
+    8.367196987588669e-11
+   -4.309482817120374e-13
+   -1.944868405567585e-12
+   -2.213828380054223e-11
+    7.979216395169359e-11
+ 6.53e+10    
+    7.990190708972185e-11
+    -2.21404212543015e-11
+    8.364751547962615e-11
+   -1.945408203472335e-12
+   -1.116888262166009e-11
+    8.366942616453624e-11
+      -4.266329792532e-13
+   -1.943769553741168e-12
+   -2.214288388737166e-11
+    7.978192710053714e-11
+ 6.54e+10    
+    7.989157062615314e-11
+   -2.214500234517034e-11
+    8.364495048403799e-11
+   -1.944272114494232e-12
+   -1.117411236371631e-11
+    8.366686495364074e-11
+   -4.223126314044851e-13
+   -1.942652701864795e-12
+   -2.214747732555912e-11
+    7.977166295268364e-11
+ 6.55e+10    
+    7.988120667166733e-11
+   -2.214957659261452e-11
+    8.364236786510601e-11
+   -1.943117999212037e-12
+   -1.117935124468427e-11
+    8.366428619914624e-11
+   -4.179873654248377e-13
+   -1.941517858497032e-12
+   -2.215206402456312e-11
+    7.976137149669182e-11
+ 6.56e+10    
+    7.987081521514898e-11
+   -2.215414390586121e-11
+    8.363976757876043e-11
+   -1.941945866977545e-12
+   -1.118459925927168e-11
+    8.366168985708577e-11
+   -4.136573086880204e-13
+   -1.940365032589921e-12
+   -2.215664389384729e-11
+     7.97510527212203e-11
+ 6.57e+10    
+    7.986039624558537e-11
+   -2.215870419414571e-11
+    8.363714958102053e-11
+    -1.94075572753672e-12
+   -1.118985640206682e-11
+     8.36590758835805e-11
+   -4.093225886754641e-13
+   -1.939194233488473e-12
+   -2.216121684288298e-11
+    7.974070661502764e-11
+ 6.58e+10    
+    7.984994975206573e-11
+   -2.216325736671375e-11
+    8.363451382799505e-11
+   -1.939547591029094e-12
+   -1.119512266753809e-11
+     8.36564442348393e-11
+   -4.049833329690776e-13
+   -1.938005470930115e-12
+   -2.216578278115109e-11
+    7.973033316697121e-11
+ 6.59e+10    
+    7.983947572378152e-11
+    -2.21678033328237e-11
+    8.363186027588243e-11
+   -1.938321467987252e-12
+   -1.120039805003327e-11
+    8.365379486715919e-11
+   -4.006396692440607e-13
+   -1.936798755044168e-12
+   -2.217034161814445e-11
+    7.971993236600751e-11
+ 6.6e+10     
+    7.982897415002542e-11
+   -2.217234200174868e-11
+    8.362918888097095e-11
+   -1.937077369336177e-12
+   -1.120568254377915e-11
+    8.365112773692586e-11
+   -3.962917252616949e-13
+   -1.935574096351263e-12
+   -2.217489326337002e-11
+    7.970950420119193e-11
+ 6.61e+10    
+     7.98184450201913e-11
+   -2.217687328277895e-11
+    8.362649959963915e-11
+   -1.935815306392727e-12
+    -1.12109761428809e-11
+    8.364844280061354e-11
+   -3.919396288620813e-13
+   -1.934331505762776e-12
+   -2.217943762635103e-11
+    7.969904866167753e-11
+ 6.62e+10    
+    7.980788832377443e-11
+   -2.218139708522405e-11
+    8.362379238835593e-11
+   -1.934535290864987e-12
+   -1.121627884132163e-11
+    8.364574001478557e-11
+   -3.875835079569101e-13
+   -1.933070994580264e-12
+   -2.218397461662927e-11
+    7.968856573671571e-11
+ 6.63e+10    
+     7.97973040503698e-11
+   -2.218591331841493e-11
+    8.362106720368097e-11
+   -1.933237334851633e-12
+   -1.122159063296183e-11
+    8.364301933609439e-11
+   -3.832234905221817e-13
+   -1.931792574494826e-12
+   -2.218850414376723e-11
+    7.967805541565519e-11
+ 6.64e+10    
+      7.9786692189673e-11
+   -2.219042189170631e-11
+    8.361832400226474e-11
+   -1.931921450841342e-12
+   -1.122691151153887e-11
+    8.364028072128198e-11
+   -3.788597045909193e-13
+   -1.930496257586558e-12
+   -2.219302611735038e-11
+    7.966751768794254e-11
+ 6.65e+10    
+    7.977605273147964e-11
+   -2.219492271447884e-11
+    8.361556274084898e-11
+   -1.930587651712129e-12
+   -1.123224147066661e-11
+    8.363752412718035e-11
+   -3.744922782458554e-13
+   -1.929182056323839e-12
+   -2.219754044698948e-11
+    7.965695254312074e-11
+ 6.66e+10    
+    7.976538566568481e-11
+   -2.219941569614141e-11
+    8.361278337626682e-11
+   -1.929235950730676e-12
+    -1.12375805038348e-11
+    8.363474951071139e-11
+   -3.701213396121355e-13
+    -1.92784998356279e-12
+   -2.220204704232267e-11
+    7.964635997083004e-11
+ 6.67e+10    
+    7.975469098228291e-11
+   -2.220390074613335e-11
+    8.360998586544327e-11
+   -1.927866361551668e-12
+   -1.124292860440872e-11
+    8.363195682888725e-11
+   -3.657470168499654e-13
+   -1.926500052546597e-12
+   -2.220654581301774e-11
+    7.963573996080705e-11
+ 6.68e+10    
+    7.974396867136738e-11
+   -2.220837777392657e-11
+    8.360717016539521e-11
+   -1.926478898217126e-12
+    -1.12482857656287e-11
+    8.362914603881098e-11
+   -3.613694381472909e-13
+   -1.925132276904803e-12
+   -2.221103666877441e-11
+    7.962509250288444e-11
+ 6.69e+10    
+    7.973321872313056e-11
+   -2.221284668902806e-11
+    8.360433623323193e-11
+   -1.925073575155689e-12
+   -1.125365198060973e-11
+    8.362631709767639e-11
+   -3.569887317124214e-13
+   -1.923746670652721e-12
+    -2.22155195193266e-11
+    7.961441758699118e-11
+ 6.7e+10     
+    7.972244112786326e-11
+   -2.221730740098191e-11
+    8.360148402615511e-11
+   -1.923650407181934e-12
+   -1.125902724234092e-11
+     8.36234699627687e-11
+   -3.526050257666838e-13
+   -1.922343248190702e-12
+   -2.221999427444473e-11
+    7.960371520315188e-11
+ 6.71e+10    
+     7.97116358759546e-11
+   -2.222175981937168e-11
+    8.359861350145942e-11
+   -1.922209409495636e-12
+   -1.126441154368522e-11
+    8.362060459146435e-11
+   -3.482184485370402e-13
+   -1.920922024303453e-12
+   -2.222446084393772e-11
+    7.959298534148668e-11
+ 6.72e+10    
+    7.970080295789162e-11
+   -2.222620385382264e-11
+    8.359572461653265e-11
+   -1.920750597681046e-12
+   -1.126980487737902e-11
+    8.361772094123192e-11
+   -3.438291282487044e-13
+   -1.919483014159316e-12
+   -2.222891913765552e-11
+    7.958222799221092e-11
+ 6.73e+10    
+    7.968994236425948e-11
+   -2.223063941400409e-11
+    8.359281732885603e-11
+   -1.919273987706153e-12
+   -1.127520723603161e-11
+    8.361481896963205e-11
+   -3.394371931177591e-13
+   -1.918026233309603e-12
+   -2.223336906549127e-11
+    7.957144314563535e-11
+ 6.74e+10    
+    7.967905408574082e-11
+   -2.223506640963152e-11
+    8.358989159600458e-11
+   -1.917779595921916e-12
+   -1.128061861212497e-11
+    8.361189863431758e-11
+   -3.350427713437608e-13
+   -1.916551697687802e-12
+   -2.223781053738355e-11
+    7.956063079216542e-11
+ 6.75e+10    
+    7.966813811311549e-11
+   -2.223948475046892e-11
+     8.35869473756472e-11
+   -1.916267439061522e-12
+   -1.128603899801333e-11
+    8.360895989303445e-11
+   -3.306459911023298e-13
+   -1.915059423608878e-12
+   -2.224224346331869e-11
+    7.954979092230139e-11
+ 6.76e+10    
+    7.965719443726098e-11
+   -2.224389434633118e-11
+    8.358398462554731e-11
+   -1.914737534239588e-12
+   -1.129146838592286e-11
+    8.360600270362162e-11
+   -3.262469805377514e-13
+   -1.913549427768499e-12
+   -2.224666775333304e-11
+    7.953892352663803e-11
+ 6.77e+10    
+    7.964622304915149e-11
+    -2.22482951070862e-11
+    8.358100330356283e-11
+   -1.913189898951366e-12
+    -1.12969067679513e-11
+    8.360302702401119e-11
+   -3.218458677555776e-13
+   -1.912021727242303e-12
+    -2.22510833175151e-11
+    7.952802859586462e-11
+ 6.78e+10    
+    7.963522393985815e-11
+    -2.22526869426572e-11
+    8.357800336764689e-11
+    -1.91162455107198e-12
+   -1.130235413606757e-11
+    8.360003281222911e-11
+   -3.174427808151854e-13
+   -1.910476339485105e-12
+   -2.225549006600803e-11
+    7.951710612076448e-11
+ 6.79e+10    
+    7.962419710054877e-11
+   -2.225706976302504e-11
+    8.357498477584737e-11
+   -1.910041508855582e-12
+    -1.13078104821116e-11
+    8.359702002639551e-11
+   -3.130378477224003e-13
+   -1.908913282330071e-12
+    -2.22598879090118e-11
+    7.950615609221507e-11
+ 6.8e+10     
+    7.961314252248795e-11
+   -2.226144347823066e-11
+    8.357194748630854e-11
+    -1.90844079093452e-12
+   -1.131327579779389e-11
+    8.359398862472464e-11
+   -3.086311964220653e-13
+   -1.907332573988005e-12
+   -2.226427675678543e-11
+    7.949517850118801e-11
+ 6.81e+10    
+     7.96020601970365e-11
+   -2.226580799837706e-11
+    8.356889145726999e-11
+   -1.906822416318526e-12
+   -1.131875007469531e-11
+    8.359093856552558e-11
+   -3.042229547906289e-13
+   -1.905734233046478e-12
+   -2.226865651964936e-11
+    7.948417333874853e-11
+ 6.82e+10    
+    7.959095011565126e-11
+   -2.227016323363169e-11
+    8.356581664706767e-11
+   -1.905186404393874e-12
+   -1.132423330426672e-11
+    8.358786980720243e-11
+   -2.998132506287307e-13
+   -1.904118278469019e-12
+   -2.227302710798765e-11
+    7.947314059605549e-11
+ 6.83e+10    
+    7.957981226988561e-11
+   -2.227450909422898e-11
+    8.356272301413428e-11
+   -1.903532774922497e-12
+   -1.132972547782878e-11
+    8.358478230825466e-11
+   -2.954022116538093e-13
+   -1.902484729594303e-12
+   -2.227738843225041e-11
+    7.946208026436168e-11
+ 6.84e+10    
+    7.956864665138879e-11
+    -2.22788454904723e-11
+    8.355961051699919e-11
+   -1.901861548041132e-12
+   -1.133522658657166e-11
+    8.358167602727737e-11
+   -2.909899654926814e-13
+   -1.900833606135264e-12
+   -2.228174040295584e-11
+    7.945099233501284e-11
+ 6.85e+10    
+    7.955745325190598e-11
+    -2.22831723327365e-11
+    8.355647911428927e-11
+   -1.900172744260453e-12
+    -1.13407366215548e-11
+     8.35785509229619e-11
+   -2.865766396741453e-13
+    -1.89916492817831e-12
+   -2.228608293069285e-11
+    7.943987679944878e-11
+ 6.86e+10    
+    7.954623206327811e-11
+   -2.228748953147001e-11
+    8.355332876472884e-11
+   -1.898466384464135e-12
+   -1.134625557370668e-11
+    8.357540695409563e-11
+   -2.821623616215933e-13
+   -1.897478716182394e-12
+   -2.229041592612293e-11
+    7.942873364920198e-11
+ 6.87e+10    
+    7.953498307744199e-11
+   -2.229179699719733e-11
+    8.355015942714014e-11
+   -1.896742489908016e-12
+   -1.135178343382455e-11
+     8.35722440795632e-11
+    -2.77747258645613e-13
+   -1.895774990978168e-12
+   -2.229473929998296e-11
+    7.941756287589872e-11
+ 6.88e+10    
+    7.952370628642998e-11
+   -2.229609464052118e-11
+    8.354697106044372e-11
+   -1.895001082219127e-12
+   -1.135732019257423e-11
+    8.356906225834605e-11
+   -2.733314579366179e-13
+   -1.894053773767104e-12
+   -2.229905296308703e-11
+    7.940636447125823e-11
+ 6.89e+10    
+    7.951240168237003e-11
+   -2.230038237212484e-11
+    8.354376362365889e-11
+   -1.893242183394787e-12
+   -1.136286584048999e-11
+    8.356586144952291e-11
+   -2.689150865574608e-13
+   -1.892315086120569e-12
+   -2.230335682632892e-11
+    7.939513842709282e-11
+ 6.9e+10     
+     7.95010692574857e-11
+   -2.230466010277454e-11
+    8.354053707590376e-11
+   -1.891465815801686e-12
+   -1.136842036797426e-11
+    8.356264161227077e-11
+   -2.644982714360784e-13
+   -1.890558949978939e-12
+   -2.230765080068447e-11
+    7.938388473530807e-11
+ 6.91e+10    
+    7.948970900409625e-11
+   -2.230892774332164e-11
+    8.353729137639575e-11
+   -1.889672002174909e-12
+   -1.137398376529745e-11
+    8.355940270586453e-11
+   -2.600811393581468e-13
+   -1.888785387650666e-12
+   -2.231193479721379e-11
+    7.937260338790271e-11
+ 6.92e+10    
+    7.947832091461595e-11
+   -2.231318520470495e-11
+    8.353402648445217e-11
+   -1.887860765617001e-12
+   -1.137955602259786e-11
+    8.355614468967783e-11
+   -2.556638169597183e-13
+   -1.886994421811358e-12
+   -2.231620872706356e-11
+    7.936129437696828e-11
+ 6.93e+10    
+    7.946690498155482e-11
+   -2.231743239795309e-11
+     8.35307423594904e-11
+    -1.88603212959696e-12
+   -1.138513712988146e-11
+    8.355286752318295e-11
+   -2.512464307199198e-13
+   -1.885186075502826e-12
+   -2.232047250146928e-11
+    7.934995769468962e-11
+ 6.94e+10    
+    7.945546119751822e-11
+   -2.232166923418674e-11
+    8.352743896102798e-11
+   -1.884186117949329e-12
+   -1.139072707702171e-11
+    8.354957116595161e-11
+   -2.468291069535992e-13
+   -1.883360372132154e-12
+   -2.232472603175763e-11
+    7.933859333334432e-11
+ 6.95e+10    
+    7.944398955520707e-11
+   -2.232589562462098e-11
+    8.352411624868356e-11
+   -1.882322754873126e-12
+   -1.139632585375955e-11
+     8.35462555776554e-11
+   -2.424119718040634e-13
+   -1.881517335470707e-12
+    -2.23289692293488e-11
+    7.932720128530352e-11
+ 6.96e+10    
+    7.943249004741763e-11
+   -2.233011148056766e-11
+    8.352077418217684e-11
+   -1.880442064930901e-12
+   -1.140193344970315e-11
+    8.354292071806571e-11
+   -2.379951512357636e-13
+   -1.879656989653164e-12
+   -2.233320200575862e-11
+    7.931578154303097e-11
+ 6.97e+10    
+     7.94209626670414e-11
+   -2.233431671343738e-11
+    8.351741272132899e-11
+    -1.87854407304769e-12
+   -1.140754985432786e-11
+    8.353956654705441e-11
+   -2.335787710270343e-13
+   -1.877779359176563e-12
+   -2.233742427260108e-11
+    7.930433409908381e-11
+ 6.98e+10    
+    7.940940740706561e-11
+   -2.233851123474226e-11
+    8.351403182606332e-11
+   -1.876628804510014e-12
+   -1.141317505697611e-11
+     8.35361930245944e-11
+   -2.291629567628386e-13
+   -1.875884468899261e-12
+   -2.234163594159042e-11
+    7.929285894611214e-11
+ 6.99e+10    
+    7.939782426057275e-11
+   -2.234269495609785e-11
+     8.35106314564051e-11
+    -1.87469628496484e-12
+   -1.141880904685725e-11
+    8.353280011075949e-11
+   -2.247478338275295e-13
+   -1.873972344039975e-12
+   -2.234583692454357e-11
+    7.928135607685955e-11
+ 7e+10       
+    7.938621322074103e-11
+   -2.234686778922564e-11
+    8.350721157248263e-11
+   -1.872746540418529e-12
+   -1.142445181304755e-11
+    8.352938776572516e-11
+   -2.203335273976321e-13
+   -1.872043010176729e-12
+   -2.235002713338225e-11
+     7.92698254841625e-11
* NOTE: Solution at 1e+08 Hz used as DC point.

.ends
