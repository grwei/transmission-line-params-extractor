* BEGIN ANSOFT HEADER
* node 1    1:trace_p_0_T1_A
* node 2    1:trace_n_0_T1_A
* node 3    1:trace_n_1_T1_A
* node 4    1:trace_p_1_T1_A
* node 5    Ground_A
* node 6    1:trace_p_0_T1_B
* node 7    1:trace_n_0_T1_B
* node 8    1:trace_n_1_T1_B
* node 9    1:trace_p_1_T1_B
* node 10   Ground_B
*  Project: 4lines
*   Design: 2-diff-pairs
*   Length: 5
*   Format: HSPICE
*  Creator: Ansoft HFSS
*     Date: Sat Jun 06 09:41:10 2020
* END ANSOFT HEADER

.subckt ckt_m4lines_port_W 1 2 3 4 inref 5 6 7 8 outref length=5.08M

.model m4lines_port_1 W MODELTYPE=table N=4 RMODEL=r_m4lines_port_1
+ LMODEL=l_m4lines_port_1 GMODEL=g_m4lines_port_1 CMODEL=c_m4lines_port_1

* Example usage:
W1 1 2 3 4 inref 5 6 7 8 outref N=4 L=length TABLEMODEL=m4lines_port_1

.model r_m4lines_port_1 sp N=4 SPACING=nonuniform VALTYPE=real
+ INTERPOLATION=spline
+ DATA = 700
+ 0           
+        7.125307581499241
+       0.6582573515222506
+        7.240611774399657
+       0.2632193777876676
+       0.9049689635842689
+        7.260698002125167
+      0.09583671641050204
+       0.2621687410268075
+       0.6381229697293089
+        7.123771171105417
+ 2e+08       
+        10.68201877115167
+       0.9946157371956403
+        10.81326330563095
+       0.3660339899515054
+        1.320626901512357
+        10.84730515947828
+       0.1294697305661216
+       0.3661100477548065
+       0.9619272712194548
+        10.68189060635637
+ 3e+08       
+        13.16803574153734
+        1.109954178989794
+        13.31046467609029
+       0.4219424955503647
+        1.585340516285568
+        13.35992152634004
+       0.1371198524336372
+       0.4225134002200347
+        1.069513144822761
+         13.1731876910728
+ 4e+08       
+        15.28931954253306
+        1.211161828205024
+        15.44485497542442
+       0.4615168841120507
+        1.810674229586082
+        15.51017825065585
+       0.1359146478887154
+       0.4621682891876723
+         1.16235258523667
+        15.30074569927285
+ 5e+08       
+        17.23827617060569
+        1.328149939031001
+        17.40287737113308
+       0.4984667968397924
+        2.018927854728304
+        17.48331042521506
+       0.1360167967970909
+       0.4992193370844184
+        1.271377188946144
+        17.25676113958263
+ 6e+08       
+        19.04053167131416
+        1.443688958021776
+        19.20826104488582
+       0.5344540644259039
+        2.210319212211583
+        19.30219922821312
+       0.1386519144449953
+       0.5354208454114844
+         1.37958808187008
+        19.06654865669796
+ 7e+08       
+        20.70445273123923
+        1.547240858004157
+         20.8708051510677
+        0.568647662247094
+          2.3850664757079
+        20.97654761982336
+       0.1425967315598275
+       0.5699046269442996
+        1.476292492398342
+        20.73818714333684
+ 8e+08       
+        22.24954237385164
+        1.639105672495061
+        22.41253133208093
+       0.6004411260143098
+        2.545906463109019
+         22.5288944092346
+       0.1465951712684085
+        0.602004122360006
+        1.561657633027426
+        22.29101695159466
+ 9e+08       
+        23.70406164368878
+        1.725396003225525
+        23.86365921771039
+       0.6298366535482756
+         2.69686650676344
+        23.99027107056513
+       0.1499098254081976
+       0.6316713990684375
+        1.641752357260546
+        23.75323760055377
+ 1e+09       
+        25.09881826889098
+        1.813812297971196
+         25.2555603810553
+       0.6572543727972335
+          2.8420576047071
+        25.39289332211205
+       0.1522719100559825
+       0.6592920546841539
+        1.724287576546017
+        25.15564670310066
+ 1.1e+09     
+        26.61064338580676
+        1.814247308517565
+         26.7946911284368
+       0.6397067901361019
+        2.968027014749377
+        26.95174280859415
+      0.09851101010940977
+       0.6426017260987825
+        1.721815523818056
+        26.67716583630504
+ 1.2e+09     
+        28.01603059080271
+        1.827339551655135
+        28.22767815453798
+       0.6287430067869149
+         3.09483431692426
+        28.40365202004607
+      0.04743746778408298
+       0.6324690871160593
+        1.732276761178209
+        28.09214772749482
+ 1.3e+09     
+        29.32225138975703
+        1.851001501568814
+        29.56020288138691
+       0.6241277227041446
+        3.220558578919787
+        29.75406351243931
+    0.0007324942406624901
+       0.6286123723671675
+        1.753397916245522
+        29.40772209571553
+ 1.4e+09     
+        30.53998343686792
+        1.883595494956915
+        30.80167860903124
+       0.6255025708135089
+        3.343932621460317
+        31.01221487002466
+      -0.0401238759735858
+       0.6306424244063351
+         1.78339427046146
+        30.63446860786138
+ 1.5e+09     
+        31.68127745959096
+        1.923871392735085
+        31.96322629230881
+       0.6324295873516875
+        3.464212136037881
+        32.18910716663267
+     -0.07393650324965861
+       0.6381047816798847
+        1.820907292238576
+         31.7843773412217
+ 1.6e+09     
+        32.75820504901645
+         1.97087125062971
+        33.05629695964056
+       0.6444206051759355
+        3.581042735478322
+        33.29611933336269
+     -0.09985152036851919
+       0.6505066087867775
+        1.864905203358586
+        32.86948924466887
+ 1.7e+09     
+        33.78203155110806
+        2.023835524646624
+        34.09180169213004
+       0.6609577944223872
+         3.69434320752572
+        34.34412996886095
+      -0.1173827764479888
+        0.667334450166742
+         1.91458354063016
+        33.90106196935354
+ 1.8e+09     
+        34.76276836554231
+         2.08212612270099
+        35.07961482465616
+       0.6815090402905255
+        3.804211561457782
+        35.34301279431811
+      -0.1264093396113209
+       0.6880669456554092
+        1.969282404205717
+        34.88911594626562
+ 1.9e+09     
+        35.70898473278334
+        2.145170492796838
+        36.02833753067396
+       0.7055404827738911
+        3.910854047871867
+        36.30139333060818
+      -0.1271478348612377
+       0.7121850559777035
+        2.028425272094096
+        35.84224100498983
+ 2e+09       
+         36.6277875189646
+        2.212425348526148
+        36.94523427965078
+       0.7325274786707239
+        4.014534342426679
+        37.22657955361237
+      -0.1201052898028345
+       0.7391811368724082
+        2.091478257296104
+        36.76757205216198
+ 2.1e+09     
+        37.52490278189876
+        2.283356366726134
+        37.83627782669812
+       0.7619645028551718
+          4.1155390727449
+        38.12460230784745
+      -0.1060191275056606
+       0.7685673744724063
+        2.157926190127184
+        37.67086749699634
+ 2.2e+09     
+        38.40481316159279
+        2.357429718233585
+         38.7062573063932
+       0.7933740506318374
+        4.214155880533366
+        39.00032004431139
+      -0.0857910290778563
+       0.7998835987083629
+        2.227261320665004
+        38.55664432716682
+ 2.3e+09     
+        39.27092040621169
+        2.434111668645648
+          39.558918456001
+         0.82631437839914
+        4.310660679992262
+         39.8575568032572
+     -0.06042073394800729
+       0.8327042518487164
+        2.298980764317327
+        39.42833899625085
+ 2.4e+09     
+        40.12571337386681
+        2.512873181880424
+        40.39711556724625
+       0.8603858604538619
+        4.405311387565559
+        40.69925286752114
+     -0.03094467485360264
+       0.8666442290014178
+        2.372589497030607
+        40.28847432179537
+ 2.5e+09     
+        40.97092956344301
+         2.59319720216322
+        41.22296225584404
+       0.8952357834446096
+        4.498346001943302
+        41.52761495946508
+     0.001617090570133595
+       0.9013633570627171
+        2.447606454849213
+        41.13882032255019
+ 2.6e+09     
+        41.80770346989358
+        2.674586955170286
+        42.03797330349713
+        0.930561494634403
+        4.589983440269053
+        42.34425799936312
+      0.03630365357710885
+       0.9365693818526653
+        2.523571970754486
+        41.98054218493232
+ 2.7e+09     
+        42.63669852176349
+        2.756574151960449
+        42.84319330151177
+       0.9661119270619937
+        4.680425966877555
+        43.15033391418539
+       0.0722450454440634
+       0.9720194490291736
+        2.600055340240486
+        42.81433203007306
+ 2.8e+09     
+        43.45822157075133
+        2.838726395876862
+        43.63931010150771
+         1.00168761901827
+        4.769862387546594
+        43.94664527256977
+       0.1086834009245546
+        1.007520166824703
+        2.676661739272815
+        43.64052338201492
+ 2.9e+09     
+        44.27232025560054
+        2.920653396863294
+        44.42675252487236
+        1.037139414225644
+        4.858471437774086
+         44.7337429897692
+       0.1449845801858739
+        1.042926414486769
+        2.753038037177604
+        44.45918860491278
+ 3e+09       
+         45.0788643363556
+        3.002011810090047
+         45.2057726658884
+        1.072366069210203
+         4.94642498332084
+        45.51200826115459
+        0.180641764611488
+        1.078139105893338
+         2.82887727286556
+        45.27022036324011
+ 3.1e+09     
+        45.87761248805042
+        3.082508657381571
+         45.9765136341538
+        1.107311008117669
+        5.033890789959847
+        46.28171943359432
+       0.2152727145417269
+        1.113102135735039
+        2.903921716689141
+         46.0733985621949
+ 3.2e+09     
+        46.66826619256321
+        3.161903379401085
+        46.73906385327989
+         1.14195845834657
+        5.121034719840747
+        47.04310484291642
+        0.248612355533581
+        1.147798731737491
+        2.977964541095383
+        46.86844438341758
+ 3.3e+09     
+        47.45051236751126
+        3.240008619330088
+        47.49349915667518
+        1.176329179533593
+        5.208022284500801
+        47.79638282294052
+       0.2805022085308289
+        1.182247417486619
+        3.050850186701604
+         47.6550630379302
+ 3.4e+09     
+         48.2240562847073
+        3.316689866942373
+        48.23991395933938
+        1.210475969851904
+        5.295019537361936
+        48.54179018689911
+       0.3108779554887593
+        1.216497762933185
+        3.122473548601738
+        48.43297677724763
+ 3.5e+09     
+        48.98864619938064
+        3.391864104473797
+        48.97844277736944
+        1.244479102281984
+        5.382193327462362
+        49.27960053271968
+       0.3397561803615896
+        1.250626068810728
+        3.192778129472754
+        49.20194957671158
+ 3.6e+09     
+        49.74409096175835
+        3.465497598856514
+        49.70927333922869
+        1.278441813033446
+        5.469710965307538
+        50.01013375064242
+       0.3672210775839713
+         1.28473110077106
+        3.261753317484545
+        49.96180475915108
+ 3.7e+09     
+        50.49027173122987
+        3.537602982929803
+        50.43265249864542
+        1.312485936788484
+        5.557739373762775
+        50.73375812447916
+       0.3934116959501228
+         1.31892996140483
+        3.329430951987851
+        50.71243667871722
+ 3.8e+09     
+        51.22714876990895
+        3.608235763730383
+        51.14888612434964
+        1.346747759914019
+         5.64644381339915
+        51.45088641801328
+       0.4185100952282705
+        1.353354164696035
+        3.395881340643041
+        51.45381744400794
+ 3.9e+09     
+        51.95476416214334
+        3.677490390273309
+        51.85833410742467
+        1.381374143423342
+        5.735986283382815
+        52.16196732235723
+       0.4427306391304815
+        1.388145958221314
+        3.461208889060377
+        52.18599953168088
+ 4e+09       
+        52.67324119165523
+        3.745496006893201
+        52.56140159017504
+        1.416518951897545
+        5.826523706081401
+        52.86747360301926
+       0.4663105300626444
+        1.423454923326888
+        3.525547498419938
+        52.90911502894075
+ 4.1e+09     
+        53.38278100891387
+        3.812412011232751
+         53.2585274766359
+        1.452339812161944
+         5.91820600600103
+        53.56788822142843
+       0.4895016045059064
+        1.459434872039583
+        3.589055877837819
+        53.62337214597506
+ 4.2e+09     
+        54.08365713725552
+        3.878423528072871
+        53.95017122934495
+        1.488995215532846
+        6.011174191378968
+        54.26368961088204
+       0.5125633478725358
+         1.49624105087953
+        3.651912906297969
+        54.32904955680735
+ 4.3e+09     
+        54.77620829575589
+        3.943736901056725
+        54.63679888564771
+        1.526641969241127
+        6.105558539788296
+        54.95533716028115
+       0.5357570489629999
+        1.534027655313603
+        3.714313163782199
+        55.02648905766144
+ 4.4e+09     
+        55.46082995810708
+        4.008575293700223
+        55.31886913708465
+        1.565432995674454
+        6.201476977763425
+        55.64325780307535
+       0.5593409918033252
+        1.572945653662674
+        3.776462733082661
+        55.71608697393474
+ 4.5e+09     
+        56.13796501781964
+        4.073174478805456
+        55.99682020688515
+        1.605515472003147
+        6.299033729335405
+        56.32783442941933
+       0.5835665723749215
+        1.613140915320876
+        3.838575353271164
+        56.39828469825344
+ 4.6e+09     
+         56.8080938889998
+        4.137778881630218
+        56.67105813516702
+        1.647029297377546
+        6.398318290369872
+        57.00939664536891
+        0.608675226015952
+        1.654752634774348
+        3.900868983798663
+        57.07355870083046
+ 4.7e+09     
+        57.47172433688065
+        4.202637927258955
+        57.34194694317511
+        1.690105870155452
+        6.499404765858337
+        57.68821420454953
+       0.6348960552556697
+        1.697912039880555
+        3.963562815775108
+        57.74241031755745
+ 4.8e+09     
+        58.12938130149065
+        4.268002727108806
+        58.00980100258663
+        1.734867153582697
+        6.602351587075514
+        58.36449324623878
+       0.6624440553811286
+        1.742741370071551
+        4.026874745257533
+        58.40535558920247
+ 4.9e+09     
+         58.7815969498301
+        4.334123124049253
+         58.6748797904545
+        1.781425005096767
+        6.707201606037532
+         59.0383752996096
+       0.6915188445281535
+        1.789353107564129
+        4.091019303420691
+        59.06291539526773
+ 5e+09       
+        59.42890116542048
+        4.401245100923241
+        59.33738507192263
+          1.8298807420483
+        6.813982547112167
+        59.70993886557795
+       0.7223038153901566
+        1.837849442347283
+         4.15620602117537
+        59.71560609724655
+ 5.1e+09     
+        60.07181265809823
+        4.469608544004088
+        59.99746042812683
+        1.880324915198573
+        6.922707780858378
+         60.3792032712624
+       0.7549656359633286
+        1.888321949762664
+         4.22263819175831
+        60.36393087729714
+ 5.2e+09     
+        60.71083085074016
+        4.539445341669852
+        60.65519294122812
+        1.932837260863839
+        7.033377373831102
+        61.04613441050103
+       0.7896540365825628
+        1.940851457986536
+        4.290511984355954
+        61.00837192910392
+ 5.3e+09     
+        61.34642867278809
+        4.610977789727905
+         61.3106167661926
+         1.98748680298964
+        7.145979360485458
+        61.71065193720658
+       0.8265018295430187
+        1.995508081738445
+        4.360015854963132
+        61.64938362762875
+ 5.4e+09     
+        61.97904636286248
+        4.684417268590816
+        61.96371826170574
+        2.044332077646006
+        7.260491179444415
+        62.37263746401296
+        0.865625115689213
+        2.052351398124013
+        4.431330197172062
+        62.28738677357827
+ 5.5e+09     
+        62.60908635450802
+        4.759963153909562
+        62.61444232055013
+        2.103421454290442
+        7.376881215980352
+        63.03194333212052
+       0.9071236394339106
+        2.111430740670075
+        4.504627175000945
+        62.92276397697992
+ 5.6e+09     
+        63.23690929054745
+        4.837801921158742
+        63.26269953121715
+        2.164793530480633
+        7.495110395121931
+        63.68840155366892
+       0.9510812597623346
+        2.172785588297306
+        4.580070681653375
+        63.55585621278696
+ 5.7e+09     
+        63.86283118313612
+        4.918106405741702
+         63.9083738144102
+        2.228477579353757
+        7.615133774715739
+        64.34183257901427
+       0.9975665099473585
+        2.236446027130619
+        4.657816371644729
+        64.18696055055452
+ 5.8e+09     
+        64.48712170905596
+         5.00103518305597
+        64.55133020649875
+        2.294494031959722
+        7.736902094374924
+        64.99205360174466
+        1.046633223042202
+        2.302433264586015
+         4.73801171847545
+        64.81632903073054
+ 5.9e+09     
+        65.11000360375309
+        5.086732037186938
+        65.19142250245577
+        2.362854979295624
+        7.860363243867806
+        65.63888617852378
+        1.098321203833946
+        2.370760176993413
+        4.820796055457706
+        65.44416863277063
+ 6e+09       
+        65.73165309383265
+        5.175325492031656
+        65.82850051891752
+        2.433564681525442
+          7.9854636225282
+        66.28216300425687
+        1.152656930944391
+        2.441431874019831
+        4.906300563015118
+        66.07064225588749
+ 6.1e+09     
+        66.35220128682029
+        5.266928384279259
+        66.46241678963888
+        2.506620074300433
+        8.112149369196352
+        66.92173374207687
+        1.209654275261021
+        2.514446265252985
+        4.994648171475374
+        66.69587061246607
+ 6.2e+09     
+        66.97173641955506
+        5.361637463409295
+        67.09303255719983
+        2.582011264272664
+        8.240367449621514
+        67.55746985981847
+        1.269315222967879
+         2.58979461641332
+        5.085953353878368
+        67.31993491754368
+ 6.3e+09     
+        67.59030685299726
+        5.459533009421231
+        67.72022297357162
+        2.659722007794363
+        8.370066594893625
+        68.18926846861085
+        1.331630593211335
+        2.667462084718887
+        5.180321788534064
+        67.94288024564709
+ 6.4e+09     
+        68.20792469177057
+        5.560678464126952
+        68.34388146597375
+        2.739730168419144
+        8.501198090150313
+        68.81705519444476
+        1.396580741952658
+         2.74742822488647
+        5.277849875959385
+         68.5647194188391
+ 6.5e+09     
+        68.82456990149298
+        5.665120076368447
+        68.96392326209545
+        2.822008150183405
+        8.633716417451106
+         69.4407861402497
+        1.464136244888501
+        2.829667459084224
+         5.37862409943783
+        69.18543728705667
+ 6.6e+09     
+        69.44019479575364
+        5.772886565344131
+        69.58028809953326
+        2.906523304771962
+        8.767579760326443
+        70.06044901480344
+        1.534258553508986
+         2.91414950583851
+        5.482720222828252
+        69.80499526345383
+ 6.7e+09     
+        70.05472876721556
+         5.88398880928919
+        70.19294216814762
+        2.993238311591556
+        8.902750380154544
+        70.67606351666345
+        1.606900619445454
+        3.000839764435097
+        5.590202323474759
+        70.42333598313087
+ 6.8e+09     
+         70.6680831433352
+        5.998419569037541
+        70.80187935128355
+        3.082111530519364
+         9.03919487629555
+        71.28768106739142
+        1.682007483260815
+        3.089699652744067
+        5.701121662196217
+        71.04038796279531
+ 6.9e+09     
+        71.28015605607217
+        6.116153257508798
+        71.40712184305383
+        3.173097327689229
+        9.176884342939774
+        71.89538398978608
+        1.759516824768566
+        3.180686897644484
+        5.815515396411252
+        71.65607015092023
+ 7e+09       
+        71.89083722612679
+        6.237145766951547
+        72.00872022494424
+        3.266146375150806
+        9.315794436036818
+        72.49928422476799
+        1.839359472840651
+         3.27375577833835
+        5.933405146512042
+          72.270296272171
+ 7.1e+09     
+        72.50001257504557
+        6.361334365886286
+         72.6067530867474
+        3.361205925606408
+        9.455905363593523
+        73.09952167596533
+        1.921459873480185
+        3.368857323832716
+        6.054795429638706
+         72.8829788855419
+ 7.2e+09     
+         73.1075685923566
+         6.48863767719511
+        73.20132627514619
+        3.458220063713571
+        9.597201812179874
+        73.69626226478491
+        2.005736515691938
+        3.465939466741762
+        6.179671979007892
+        73.49403309209484
+ 7.3e+09     
+        73.71339639913357
+        6.618955747774667
+        73.79257184898773
+        3.557129935649674
+        9.739672821769728
+        74.28969577152868
+        2.092102315377286
+        3.564947156326522
+        6.307999970874404
+        74.10337984479784
+ 7.4e+09     
+        74.31739546349684
+        6.752170218683012
+        74.38064681416688
+        3.657873958779306
+        9.883311620158342
+        74.88003353048362
+        2.180464958105526
+        3.665822434351169
+        6.439722184985984
+        74.71094882912749
+ 7.5e+09     
+        74.91947693708214
+        6.888144602860366
+          74.965731703719
+        3.760388013351596
+        10.02811542721234
+        75.46750603927421
+        2.270727202166538
+        3.768504477898193
+        6.574757127961361
+        75.31668089838418
+ 7.6e+09     
+        75.51956659405533
+        7.026724675370773
+        75.54802906077154
+        3.864605618190319
+         10.1740852381815
+        76.05236053542322
+        2.362787143785297
+        3.872929613749846
+        6.712997152279964
+        75.92053006164868
+ 7.7e+09     
+        76.11760736556221
+        7.167738978788487
+        76.12776187382002
+        3.970458092329363
+        10.32122559427424
+        76.63485858618868
+        2.456538446775206
+        3.979031309312719
+         6.85430660643157
+        76.52246503474666
+ 7.8e+09     
+        76.71356147235949
+        7.310999443931451
+        76.70517200576545
+        4.077874704494772
+        10.46954434770408
+        77.21527373143812
+        2.551870539222169
+        4.086740145333888
+        6.998520054123161
+        77.12247037524321
+ 7.9e+09     
+        77.30741216669277
+        7.456302123699527
+        77.28051865046493
+        4.186782812248233
+        10.61905242747104
+        77.79388921362045
+        2.648668780025345
+        4.195983775831738
+        7.145440602184552
+         77.7205472313066
+ 8e+09       
+        77.89916510124154
+        7.603428035403426
+        77.85407684344888
+        4.297107992489215
+        10.76976361125981
+        78.37099582377955
+        2.746814598275617
+        4.306686880739518
+        7.294838377848523
+        78.31671374120054
+ 8.1e+09     
+        78.48884934816147
+        7.752144104729648
+        78.42613604698447
+        4.408774164870209
+        10.92169430802207
+        78.94688988797449
+        2.846185608530278
+        4.418771116733483
+        7.446449196316323
+        78.91100512523407
+ 8.2e+09     
+        79.07651809503822
+        7.902204202453627
+         78.9969988239409
+        4.521703709516552
+        11.07486335506146
+        79.52187141436805
+        2.946655705048142
+        4.532155071591651
+        7.599973458877646
+        79.50347351531205
+ 8.3e+09     
+        79.66224904702966
+        8.053350263234544
+        79.56697960991661
+        4.635817580264339
+        11.22929183275286
+        80.09624241751997
+        3.048095137986031
+        4.646754227200043
+        7.755075320269967
+        80.09418756889589
+ 8.4e+09     
+         80.2461445657854
+         8.20531347434782
+        80.13640358882888
+        4.751035414441191
+        11.38500289939646
+        80.67030543301502
+        3.150370574432372
+        4.762480935995724
+        7.911382161398715
+        80.68323191437391
+ 8.5e+09     
+        80.82833157604793
+        8.357815521060834
+        80.70560567361328
+        4.867275640020183
+        11.54202164812412
+        81.24436223236638
+        3.253345146971129
+         4.87924441521033
+        8.068484399976846
+        81.27070647371144
+ 8.6e+09     
+        81.40896127035417
+        8.510569874552653
+        81.27492959077846
+        4.984455580780766
+        11.70037498723392
+        81.81871274511197
+        3.356878492237352
+        4.996950762760457
+        8.225935667098417
+          81.856725705991
+ 8.7e+09     
+        81.98820864110486
+        8.663283107825114
+        81.84472706527329
+        5.102491559915527
+        11.86009154482208
+        82.39365419210819
+        3.460826781649661
+        5.115502998028163
+        8.383253372278322
+        82.44141781224243
+ 8.8e+09     
+        82.56627186764226
+        8.815656224939064
+        82.41535710036042
+        5.221299002330656
+        12.02120159810199
+        82.96948043116831
+        3.565042746193711
+        5.234801130097082
+        8.539919673151905
+         83.0249239379891
+ 8.9e+09     
+        83.14337158399709
+        8.967385989119789
+        82.98718534591599
+        5.340792535705089
+        12.18373702734765
+        83.54648151339561
+        3.669375696790379
+        5.354742255266917
+        8.695382858947657
+        83.60739740537191
+ 9e+09       
+        83.71975005076642
+         9.11816623578563
+        83.56058354771598
+        5.460886090198797
+         12.3477312939678
+        84.12494344579007
+        3.773671541422305
+        5.475220684879424
+        8.849059149174154
+        84.18900300174192
+ 9.1e+09     
+        84.29567025227129
+        9.267689157322096
+        84.13592906975211
+        5.581492996538023
+        12.51321944180787
+        84.70514815299505
+        3.877772799819287
+        5.596128103665365
+        9.000334900876215
+        84.76991634638384
+ 9.2e+09     
+        84.87141493780564
+        9.415646547420291
+        84.71360448141264
+        5.702526082056561
+        12.68023812039311
+        85.28737362841527
+        3.981518616127047
+        5.717353757987443
+        9.148569209526103
+        85.35032335171408
+ 9.3e+09     
+        85.44728562349026
+        9.561730993970547
+        85.29399720138764
+        5.823897764136971
+        12.84882562846712
+        85.87189426240953
+        4.084744769611375
+        5.838784672526113
+         9.29309688034478
+        85.93041979002429
+ 9.4e+09     
+        86.02360156905358
+         9.70563701081611
+        85.87749919038045
+        5.945520140378954
+        13.01902197585333
+        86.45898133290018
+        4.187283683091433
+        5.960305893156823
+        9.433231738836444
+        86.51041097174267
+ 9.5e+09     
+        86.60069874179824
+        9.847062100074666
+        86.46450668507555
+        6.067305074722393
+        13.19086896137532
+        87.04890364159189
+         4.28896442845814
+        6.081800753019429
+        9.568270241812556
+        87.09051153639192
+ 9.6e+09     
+         87.1789287781081
+        9.985707738191149
+        87.05541996629881
+        6.189164278673196
+        13.36441026432296
+        87.64192827710868
+        4.389612728325017
+        6.203151158104932
+        9.697495343404647
+        87.67094535301604
+ 9.7e+09     
+        87.75865795112909
+        10.12128028035409
+        87.65064315485678
+        6.311009386721768
+          13.539691546748
+        88.23832148479728
+        4.489050952586055
+        6.324237888097972
+        9.820180564744604
+        88.25194552293681
+ 9.8e+09     
+         88.3402661517127
+        10.25349177935061
+        88.25058402916065
+         6.43275202500781
+        13.71676056372544
+        88.83834962175378
+        4.587098108424439
+        6.444940907737758
+        9.935594211311852
+        88.83375447434047
+ 9.9e+09     
+        88.92414588834043
+        10.38206071632772
+        88.85565385935926
+        6.554303872271262
+        13.89566727862136
+        89.44228017484008
+        4.683569822131056
+        6.565139683601735
+        10.04300367856163
+        89.41662413543753
+ 1e+10       
+        89.51070131055647
+        10.50671264223988
+        89.46626725335871
+        6.675576712139464
+        14.07646398037794
+         90.0503828191132
+        4.778278310957319
+        6.684713500991911
+        10.14167978447373
+        90.00081617082745
+ 1.01e+10    
+        89.76656630779395
+        10.48716020733756
+        89.77402248218526
+        6.715248657370281
+        14.14391881647264
+         90.3593360577789
+        4.818268850797589
+        6.724327181117335
+        10.11877366730872
+        90.26086269559036
+ 1.02e+10    
+        90.03445911212593
+        10.47578074797125
+         90.0930127065532
+        6.758554595860923
+        14.21649392243604
+        90.67955748419723
+        4.860620945394539
+        6.767577359511954
+        10.10409564299223
+        90.53288909469485
+ 1.03e+10    
+        90.31425124435104
+         10.4724687508715
+        90.42301194820696
+        6.805440630908059
+        14.29408185420827
+        91.01082543804399
+        4.905298735421717
+         6.81440997162216
+        10.09753981194692
+        90.81676653641972
+ 1.04e+10    
+        90.60580783266555
+        10.47711457043487
+        90.76379022536085
+        6.855850912836999
+        14.37657388235862
+        91.35291392033201
+        4.952264876924592
+        6.864769007473097
+        10.09899609085548
+         91.1123599052539
+ 1.05e+10    
+        90.90898784810777
+        10.48960467051912
+        91.11511391451673
+        6.909727745941586
+        14.46386017034329
+        91.70559295518561
+        5.001480599568018
+        6.918596618690227
+        10.10835045654342
+        91.41952803718925
+ 1.06e+10    
+        91.22364433803151
+         10.5098218621387
+        91.47674610457605
+        6.967011694118374
+        14.55582994675469
+        92.06862894489784
+        5.052905764551594
+        6.975833224184081
+        10.12548518577537
+        91.73812395285069
+ 1.07e+10    
+        91.54962465748233
+        10.53764553689708
+        91.84844694314411
+        7.027641685102743
+        14.65237167158327
+        92.44178501813923
+        5.106498922145836
+        7.036417614405762
+        10.15027909079637
+        92.06799508833831
+ 1.08e+10    
+        91.88677069837843
+        10.57295189601362
+        92.22997397493936
+        7.091555113218681
+        14.75337319652364
+        92.82482137119091
+        5.162217368807626
+         7.10028705408665
+         10.1826077504749
+         92.4089835236848
+ 1.09e+10    
+        92.23491911641349
+        10.61561417481875
+        92.62108247224958
+        7.158687940564132
+        14.85872191936975
+        93.21749560209625
+        5.220017203835996
+        7.167377383385624
+        10.22234373691585
+         92.7609262088389
+ 1.1e+10     
+        92.59390155560875
+        10.66550286260705
+        93.02152575737614
+        7.228974796558719
+        14.96830493255328
+        93.61956303764093
+        5.279853385531087
+        7.237623117369841
+        10.26935683743122
+        93.12365518711297
+ 1.11e+10    
+        92.96354487047071
+        10.72248591775582
+        93.43105551703135
+        7.302349075788147
+        15.08200916588854
+        94.03077705307879
+        5.341679786824118
+         7.31095754376663
+        10.32351427177267
+        93.49699781603812
+ 1.12e+10    
+        93.34367134571279
+        10.78642897802894
+        93.84942210866387
+        7.378743034086434
+          15.199721523596
+        94.45088938454288
+        5.405449250346227
+        7.387312818926723
+        10.38468090454301
+         93.8807769855959
+ 1.13e+10    
+        93.73409891352199
+        10.85719556600307
+        94.27637485869836
+         7.45808788280138
+         15.3213290156839
+        94.87965043407726
+         5.47111364290793
+        7.466620061946276
+        10.45271945271942
+         94.2748113338031
+ 1.14e+10    
+        94.13464136835928
+        10.93464728956235
+        94.71166235268156
+        7.540313881197116
+        15.44671888377367
+        95.31680956725167
+        5.538623909363997
+        7.548809446902762
+        10.52749068823336
+        94.67891545964073
+ 1.15e+10    
+        94.54510857929918
+        11.01864403742421
+        95.15503271734511
+        7.625350426951217
+        15.57577872146092
+        95.76211540331678
+        5.607930125838866
+        7.633810293162201
+         10.6088536355666
+         95.0929001333292
+ 1.16e+10    
+        94.96530669991589
+        11.10904416966816
+        95.60623389459404
+         7.71312614470923
+        15.70839658930895
+         96.2153160978702
+        5.678981552290953
+        7.721551153722617
+        10.69666576433001
+        95.51657250396644
+ 1.17e+10    
+        95.39503837574793
+        11.20570470325069
+        96.06501390744272
+        7.803568972665216
+        15.84446112457531
+         96.6761596180141
+        5.751726684396541
+        7.811959901563569
+         10.7907831768089
+        95.94973630455185
+ 1.18e+10    
+        95.83410294936196
+        11.30848149249891
+        96.53112111792213
+        7.896606247142922
+        15.98386164577701
+        97.14439400998587
+        5.826113304735085
+        7.904963813975669
+        10.89106079046281
+        96.39219205442569
+ 1.19e+10    
+         96.2822966630654
+        11.41722940458771
+        97.00430447699507
+        7.992164785152529
+        16.12648825220219
+        97.61976765925317
+        5.902088533259587
+        8.000489654848849
+        10.99735251538096
+        96.84373725917139
+ 1.2e+10     
+        96.73941285930522
+        11.53180249000845
+        97.48431376651079
+        8.090170964906365
+        16.27223191847735
+        98.10202954306413
+        5.979598877037471
+        8.098463754902419
+         11.1095114267026
+        97.30416660802352
+ 1.21e+10    
+        97.20524217881153
+        11.65205414805221
+        97.97089983324433
+        8.190550804281459
+        16.42098458430473
+        98.59092947545997
+        6.058590279249822
+        8.198812089843841
+        11.22738993201597
+        97.77327216883481
+ 1.22e+10    
+        97.67957275653703
+        11.77783728733141
+        98.46381481506445
+          8.2932300372141
+        16.57263923948237
+        99.08621834474303
+        6.139008167436807
+        8.301460356448313
+        11.35083993376522
+        98.25084358066665
+ 1.23e+10    
+        98.16219041545398
+         11.9090044813743
+        98.96281235927719
+        8.398134188024752
+        16.72709000432215
+        99.58764834341946
+         6.22079750097857
+        8.406334046551546
+        11.47971298669028
+        98.73666824406098
+ 1.24e+10    
+         98.6528788582778
+        12.04540811933235
+        99.46764783319855
+        8.505188643667028
+        16.88423220558175
+        100.0949731906144
+        6.303902817804789
+        8.513358518955787
+        11.61386045034189
+        99.23053150906091
+ 1.25e+10    
+        99.15141985717128
+        12.18690055184502
+        99.97807852700969
+        8.614318723901478
+        17.04396244802752
+        100.6079483469856
+        6.388268280322741
+        8.622459069248992
+         11.7531336367113
+        99.73221686105343
+ 1.26e+10    
+        99.65759344150484
+        12.33333423211226
+        100.4938638489504
+        8.725449749397198
+         17.2061786817425
+        101.1263312221416
+        6.473837720559825
+        8.733560997541858
+        11.89738395302449
+        100.2415061044988
+ 1.27e+10    
+        100.1711780837387
+        12.48456185223028
+        101.0147655129106
+        8.838507107767384
+        17.37078026529734
+        101.6498813745921
+        6.560554684513278
+         8.84658967412852
+        12.04646303975221
+        100.7581795446217
+ 1.28e+10    
+        100.6919508834868
+        12.64043647484729
+        101.5405477184782
+        8.953416317546052
+         17.5376680248987
+        102.1783607042484
+        6.648362475702941
+         8.96147060308191
+        12.20022290389436
+        101.2820161671359
+ 1.29e+10    
+        101.2196877498383
+        12.80081166020551
+        102.0709773235095
+        9.070103090116843
+        17.70674430962914
+        102.7115336374961
+        6.737204197924404
+        9.078129483793592
+         12.3585160475967
+        101.8127938160719
+ 1.3e+10     
+        101.7541635819876
+        12.96554158863086
+        102.6058240092806
+        9.188493389607904
+        17.87791304289333
+        103.2491673048746
+        6.827022797198461
+        9.196492270474172
+        12.52119559216628
+        102.3502893697745
+ 1.31e+10    
+        102.2951524482433
+        13.13448117854103
+        103.1448604382885
+        9.308513490765009
+        18.05107977018139
+        103.7910317113832
+        6.917761102915671
+        9.316485229628642
+        12.68811539755002
+         102.894278915145
+ 1.32e+10    
+        102.8424277634661
+        13.30748620004293
+        103.6878624047701
+         9.43009003482358
+        18.22615170326187
+         104.336899899453
+        7.009361868173507
+         9.43803499552493
+        12.85913017734705
+        103.4445379201813
+ 1.33e+10    
+        103.3957624649931
+        13.48441338419091
+        104.2346089780019
+        9.553150083393803
+        18.40303776091268
+         104.886548104616
+        7.101767809307429
+         9.56106862367664
+        13.03409560942551
+        104.0008414048864
+ 1.34e+10    
+        103.9549291870933
+        13.66512052798122
+        104.7848826384574
+        9.677621170382107
+        18.58164860629885
+         105.439755903906
+        7.194921644612995
+        9.685513642358927
+        13.21286844221642
+        104.5629641105959
+ 1.35e+10    
+        104.5197004339957
+        13.84946659515761
+        105.3384694068866
+        9.803431351968861
+        18.76189668110233
+        105.9963063570347
+        7.288766132261054
+        9.811298102181873
+        13.39530659675984
+        105.1306806677767
+ 1.36e+10    
+        105.0898487515333
+        14.03731181290531
+         105.895158966395
+        9.930509254665475
+         18.9436962365095
+        106.5559861403832
+        7.383244107406228
+        9.938350623744228
+        13.58126926457838
+        105.7037657623459
+ 1.37e+10    
+        105.6651468974247
+        14.22851776451168
+        106.4547447775957
+        10.05878412147454
+        19.12696336115771
+         107.118585673852
+        7.478298518489901
+        10.06660044339432
+        13.77061700145551
+         106.281994300547
+ 1.38e+10    
+        106.2453680102201
+        14.42294747806952
+        107.0170241869091
+        10.18818585617861
+        19.31161600614278
+        107.6838992406212
+        7.573872462738817
+        10.19597745712086
+        13.96321181719458
+        106.8651415724194
+ 1.39e+10    
+        106.8302857769303
+        14.62046551130255
+        107.5817985280885
+        10.31864506578296
+        19.49757400718465
+        108.2517250998688
+        7.669909220860884
+        10.32641226260454
+        14.15891726143759
+        107.4529834138878
+ 1.4e+10     
+        107.4196745993419
+        14.82093803259275
+        108.1488732170548
+        10.45009310113834
+        19.68475910405022
+        108.8218655925022
+        7.766352290941196
+        10.45783619945541
+        14.35759850562044
+        108.0452963674914
+ 1.41e+10    
+        108.0133097590194
+        15.02423289828283
+        108.7180578401146
+        10.58246209577293
+        19.87309495732521
+        109.3941272399615
+         7.86314542153938
+        10.59018138766602
+        14.55912242114284
+         108.641857841764
+ 1.42e+10    
+        108.6109675809898
+        15.23021972633841
+        109.2891662356548
+        10.71568500296009
+        20.06250716263099
+        109.9683208361534
+        7.960232643990436
+        10.72338076430833
+        14.76335765383108
+        109.2424462692727
+ 1.43e+10    
+        109.2124255960833
+        15.43876996644015
+        109.8620165693922
+         10.8496956310497
+         20.2529232623749
+        110.5442615325867
+         8.05755830391309
+        10.85736811850537
+        14.97017469477024
+        109.8468412633076
+ 1.44e+10    
+        109.8174627019147
+        15.64975696658706
+        110.4364314032691
+        10.98442867709491
+        20.44427275512354
+         111.121768916765
+        8.155067091926133
+        10.99207812470567
+         15.1794459475818
+        110.4548237732108
+ 1.45e+10    
+        110.4258593224578
+        15.86305603628387
+         111.012237758085
+         11.1198197587999
+        20.63648710268699
+        111.7006670839266
+        8.252704073577062
+        11.12744637429297
+        15.39104579222428
+        111.0661762383256
+ 1.46e+10    
+         111.037397566178
+        16.07854450638836
+        111.5892671699597
+        11.25580544482118
+        20.82949973499704
+        112.2807847021929
+        8.350414718484855
+           11.26340940556
+        15.60485064539154
+        111.6806827405327
+ 1.47e+10    
+        111.6518613826606
+        16.29610178569087
+        112.1673557407171
+        11.39232328345073
+        21.02324605286426
+        112.8619550712158
+        8.448144928699508
+        11.39990473207752
+        15.82073901758209
+        112.2981291553371
+ 1.48e+10    
+         112.269036717677
+         16.5156094142998
+        112.7463441822978
+        11.52931182971041
+        21.21766342869385
+        113.4440161744031
+        8.545841066281573
+         11.5368708694901
+        16.03859156691362
+        112.9183033014559
+ 1.49e+10    
+        112.8887116666075
+        16.73695111390158
+        113.3260778552887
+        11.66671067088931
+        21.41269120524039
+        114.0268107248149
+        8.643449980103144
+        11.67424736076868
+        16.25829114975515
+        113.5409950888466
+ 1.5e+10     
+        113.5106766261486
+        16.96001283496788
+        113.9064068016852
+        11.80446045055249
+        21.60827069247898
+        114.6101862048244
+        8.740919031874697
+        11.81197479995111
+        16.47972286824672
+        114.1659966651176
+ 1.51e+10    
+        114.1347244442002
+        17.18468280097465
+        114.4871857719847
+        11.94250289105092
+        21.80434516266749
+        115.1939948996362
+        8.838196121397715
+        11.94999485440081
+         16.7027741147773
+        114.7931025602366
+ 1.52e+10    
+        114.7606505678414
+        17.41085154970241
+        115.0682742467204
+         12.0807808145641
+        22.00085984367573
+        115.7780939247731
+        8.935229711047935
+         12.0882502856152
+        16.92733461348867
+        115.4221098294544
+ 1.53e+10    
+        115.3882531892807
+         17.6384119716818
+        115.6495364525542
+        12.21923816270307
+        22.19776191065268
+        116.3623452476311
+        9.031968849490116
+        12.22668496861348
+        17.15329645887284
+        116.0528181943578
+ 1.54e+10    
+        116.0173333896614
+        17.86725934584742
+        116.2308413730358
+         12.3578200147046
+        22.39500047610294
+        116.9466157032163
+         9.12836319462618
+        12.36524390993443
+        17.38055415152813
+        116.6850301819378
+ 1.55e+10    
+        116.6476952805965
+        18.09729137246321
+        116.8120627541474
+        12.49647260424532
+        22.59252657844091
+        117.5307770041819
+        9.224363035780211
+        12.50387326427354
+        17.60900463113899
+        117.3185512615734
+ 1.56e+10    
+        117.2791461432974
+        18.32840820337786
+         117.393079104757
+        12.63514333490524
+        22.79029316909204
+        118.1147057452801
+        9.319919315121002
+        12.64252034979019
+        17.83854730674077
+        117.9531899798071
+ 1.57e+10    
+         117.911496565159
+        18.56051246967322
+        117.9737736921045
+        12.77378079430903
+        22.98825509820493
+        118.6982834023593
+        9.414983648323668
+        12.78113366211339
+          18.069084084333
+        118.5887580927885
+ 1.58e+10    
+        118.5445605736432
+        18.79350930675628
+        118.5540345324343
+        12.91233476697437
+        23.18636909904026
+        119.2813963260308
+        9.509508344474119
+        12.91966288707554
+        18.30051939189909
+        119.2250706962524
+ 1.59e+10    
+        119.1781557673146
+         19.0273063769582
+        119.1337543769249
+        13.05075624589428
+        23.38459377109975
+        119.8639357301391
+        9.603446425215127
+        13.05805891220287
+        18.53276020189273
+         119.861946352893
+ 1.6e+10     
+        119.8121034438645
+        19.26181388968844
+        119.7128306930216
+        13.18899744288359
+        23.58288956205636
+        120.4457976751733
+        9.696751643137784
+         13.1962738369902
+        18.76571605124589
+        120.4992072169872
+ 1.61e+10    
+        120.4462287249516
+        19.49694461920095
+        120.2911656413253
+        13.32701179771433
+        23.78121874854602
+        121.0268830467575
+        9.789378499418211
+        13.33426098198954
+        18.99929905895681
+        121.1366791561159
+ 1.62e+10    
+        121.0803606777025
+        19.73261392002116
+        120.8686660481616
+        13.46475398606991
+        23.97954541588081
+        121.6070975293672
+        9.881282260702273
+        13.47197489673827
+        19.23342394131004
+        121.7741918698262
+ 1.63e+10    
+        121.7143324326804
+        19.96873974008626
+        121.4452433739732
+        13.60217992634355
+        24.17783543674024
+        122.1863515754191
+        9.972418975237851
+        13.60937136655528
+        19.46800802478312
+        122.4115790050776
+ 1.64e+10    
+        122.3479812981596
+        20.20524263164475
+        122.0208136776746
+        13.73924678530778
+        24.37605644889763
+        122.7645603698776
+        10.06274548825761
+          13.746407418231
+        19.70297125668982
+        123.0486782682991
+ 1.65e+10    
+        122.9811488705197
+        20.44204575996588
+        122.5952975771074
+        13.87591298268198
+        24.57417783203694
+        123.3416437905471
+        10.15221945661204
+        13.88304132463833
+         19.9382362136138
+        123.6853315339023
+ 1.66e+10    
+        123.6136811405815
+        20.67907490990245
+        123.1686202057481
+        14.01213819462266
+        24.77217068371355
+         123.917526364187
+        10.24079936265505
+        14.01923260829001
+        20.17372810767766
+        124.3213849490653
+ 1.67e+10    
+        124.2454285956981
+        20.91625849035486
+        123.7407111658023
+        14.14788335616381
+          24.970007794512
+        124.4921372186263
+        10.32844452738261
+        14.15494204386778
+        20.40937479069942
+        124.9566890346317
+ 1.68e+10    
+        124.8762463174322
+         21.1535275366787
+        124.3115044778454
+        14.28311066263047
+        25.16766362245273
+         125.065410031028
+        10.41511512282604
+        14.29013165974932
+        20.64510675628173
+        125.5910987819399
+ 1.69e+10    
+        125.5059940746281
+        21.39081571107998
+        124.8809385271416
+        14.41778357005257
+        25.36511426669681
+        125.6372829724716
+        10.50077218370135
+        14.42476473855626
+        20.88085713988033
+        126.2244737454189
+ 1.7e+10     
+        126.1345364117094
+        21.62805930104121
+        125.4489560068053
+        14.55186679460235
+        25.56233744059977
+        126.2076986490137
+        10.58537761831568
+        14.55880581674942
+        21.11656171689763
+        126.8566781307762
+ 1.71e+10    
+        126.7617427320254
+        21.86519721581828
+        126.0155038579452
+        14.68532631107997
+        25.75931244416097
+        126.7766040394035
+        10.66889421873293
+        14.69222068329364
+        21.35215889884494
+        127.4875808786086
+ 1.72e+10    
+        127.3874873760771
+        22.10217098105145
+        126.5805332069429
+        14.81812935047189
+         25.9560201359165
+         127.343950429608
+        10.75128567019997
+        14.82497637741704
+        21.58758972761821
+        128.1170557432732
+ 1.73e+10    
+        128.0116496944597
+        22.33892473152939
+        127.1439993000204
+        14.95024439660518
+        26.15244290432102
+         127.909693344324
+        10.83251655983553
+        14.95704118548781
+        21.82279786793009
+        128.7449813668518
+ 1.74e+10    
+        128.6341141153587
+        22.57540520214649
+        127.7058614352409
+        15.08164118192291
+        26.34856463866403
+        128.4737924756475
+        10.91255238458402
+        15.08838463703116
+        22.05772959793899
+        129.3712413480487
+ 1.75e+10    
+        129.2547702064529
+        22.81156171709418
+           128.2660828921
+        15.21229068240095
+        26.54437069956206
+        129.0362116090599
+         10.9913595584361
+        15.21897749990936
+        22.29233379812016
+        129.9957243058794
+ 1.76e+10    
+         129.873512731076
+          23.047346177324
+        128.8246308588529
+        15.34216511163278
+        26.73984788907236
+        129.5969185469131
+        11.06890541891982
+        15.34879177468805
+        22.52656193841859
+        130.6183239379908
+ 1.77e+10    
+        130.4902416985036
+        23.28271304632296
+        129.3814763577303
+        15.47123791410315
+        26.93498442046753
+        130.1558850295738
+        11.14515823286444
+        15.47780068821015
+        22.76036806372376
+        131.2389390734795
+ 1.78e+10    
+        131.1048624082363
+        23.51761933423937
+          129.93659416819
+        15.59948375767424
+        27.12976988771133
+        130.7130866543997
+         11.2200872014405
+         15.6059786863998
+        22.99370877770934
+         131.857473720078
+ 1.79e+10    
+         131.717285488168
+        23.75202458039906
+        130.4899627483542
+        15.72687852530646
+         27.3241952346762
+        131.2685027927129
+        11.29366246448039
+        15.73330142631799
+        23.22654322507768
+        132.4738371055832
+ 1.8e+10     
+        132.3274269265295
+        23.98589083424957
+        131.0415641547802
+        15.85339930603715
+         27.5182527241397
+        131.8221165049395
+        11.36585510408268
+        15.85974576749193
+        23.45883307224833
+        133.0879437134111
+ 1.81e+10    
+        132.9352080975132
+        24.21918263477249
+        131.5913839607041
+        15.97902438523878
+        27.71193590659725
+        132.3739144540785
+        11.43663714750612
+        15.98528976253896
+        23.69054248653365
+        133.6997133121831
+ 1.82e+10    
+        133.5405557805072
+        24.45186698840509
+        132.1394111729124
+        16.10373323417998
+        27.90523958892737
+         132.923886817664
+        11.50598156935729
+        16.10991264710712
+        23.92163811383915
+        134.3090709792408
+ 1.83e+10    
+        134.1434021728602
+        24.68391334550567
+        132.6856381473714
+        16.22750649891021
+        28.09815980294364
+        133.4720271983813
+        11.57386229307796
+        16.23359482915226
+        24.15208905493127
+        134.9159471180143
+ 1.84e+10    
+        134.7436848961258
+        24.91529357540951
+        133.2300605037639
+        16.35032598849227
+        28.29069377386869
+        134.0183325334976
+        11.64025419173843
+        16.35631787757454
+        24.38186684031278
+        135.5202774691811
+ 1.85e+10    
+        135.3413469957533
+        25.14598194011031
+        133.7726770390676
+        16.47217466260259
+        28.48283988876129
+        134.5628030032598
+        11.70513308814311
+        16.47806451023423
+        24.61094540374668
+        136.1220031155456
+ 1.86e+10    
+         135.936336934189
+        25.37595506661108
+        134.3134896403087
+        16.59303661852299
+        28.67459766492943
+        135.1054419384176
+        11.76847575425608
+        16.59881858136721
+        24.83930105446786
+        136.7210704806092
+ 1.87e+10    
+         136.528608577387
+        25.60519191798422
+        134.8525031966277
+        16.71289707754542
+        28.86596771835927
+        135.6462557270195
+        11.83025990995374
+        16.71856506842237
+        25.06691244812929
+        137.3174313208004
+ 1.88e+10    
+        137.1181211747262
+        25.83367376318448
+        135.3897255107845
+        16.83174237081182
+        29.05695173219043
+        136.1852537206288
+        11.89046422111393
+        16.83729005834121
+        25.29376055651856
+        137.9110427113453
+ 1.89e+10    
+        137.7048393323638
+        26.06138414565534
+        135.9251672102336
+        16.94955992461103
+        29.24755242526552
+        136.7224481401072
+        11.94906829704949
+        16.95498073329936
+        25.51982863609067
+        138.5018670257854
+ 1.9e+10     
+        138.2887329800492
+        26.28830885077343
+        136.4588416578866
+        17.06633824515482
+        29.43777352078038
+         137.257853981099
+        12.00605268729671
+         17.0716253559334
+        25.74510219535913
+         139.089871909152
+ 1.91e+10    
+        138.8697773314645
+        26.51443587217428
+        136.9907648626935
+         17.1820669028556
+        29.62761971506375
+        137.7914889193589
+         12.0613988777681
+        17.18721325407024
+        25.96956896118802
+        139.6750302448321
+ 1.92e+10    
+        139.4479528381463
+        26.73975537700327
+          137.52095539015
+        17.29673651612718
+        29.81709664650935
+        138.3233732160563
+        12.11508928628153
+        17.30173480498318
+        26.19321884402914
+        140.2573201151681
+ 1.93e+10    
+        140.0232451370864
+        26.96425967013817
+        138.0494342728512
+        17.41033873473098
+        30.00621086468572
+        138.8535296231757
+         12.1671072574761
+        17.41518141919335
+        26.41604390214831
+        140.8367247558538
+ 1.94e+10    
+        140.5956449920954
+        27.18794315742765
+        138.5762249212027
+        17.52286622269013
+        30.19496979964702
+        139.3819832891471
+        12.21743705712741
+         17.5275455238379
+        26.63803830488545
+        141.4132325042009
+ 1.95e+10    
+        141.1651482290601
+        27.41080230799218
+        139.1013530343899
+        17.63431264079277
+        30.38338173146614
+        139.9087616648216
+        12.26606386587495
+         17.6388205456262
+        26.85919829499342
+        141.9868367413662
+ 1.96e+10    
+        141.7317556652154
+        27.63283561563567
+        139.6248465117181
+        17.74467262870766
+         30.5714557600127
+        140.4338944099052
+        12.31297377237498
+        17.74900089340398
+        27.07952215010108
+        142.5575358286479
+ 1.97e+10    
+        142.2954730325782
+        27.85404355941374
+        140.1467353644111
+        17.85394178673351
+         30.7592017749937
+        140.9574132999663
+        12.35815376589277
+         17.8580819403469
+        27.29901014334818
+        143.1253330379699
+ 1.98e+10    
+         142.856310895705
+        28.07442856340661
+        140.6670516279775
+         17.9621166572034
+        30.94663042627877
+        141.4793521341198
+        12.40159172834876
+        17.96606000580465
+        27.51766450323671
+        143.6902364766903
+ 1.99e+10    
+         143.414284563945
+        28.29399495574748
+        141.1858292752204
+        18.06919470556909
+        31.13375309452513
+        141.9997466434848
+         12.4432764258338
+        18.07293233681503
+         27.7354893727457
+         144.252259006877
+ 2e+10       
+        143.9694139983789
+         28.5127489269525
+         141.703104129995
+        18.17517430118354
+        31.32058186212156
+        142.5186344005254
+         12.4831974996092
+          18.178697089311
+        27.95249076775946
+        144.8114181592265
+ 2.01e+10    
+        144.5217237136401
+        28.73069848760362
+        142.2189137817801
+        18.28005469780645
+        31.50712948446611
+        143.0360547293465
+        12.52134545660748
+        18.28335330903901
+          28.168676534854
+         145.367736041788
+ 2.02e+10    
+         145.071242674832
+        28.94785342543313
+        142.7332975011575
+        18.38383601385339
+        31.69340936159325
+          143.55204861705
+        12.55771165945096
+        18.38690091221164
+         28.3840563084913
+        145.9212392436871
+ 2.03e+10    
+        145.6180041897673
+        29.16422526186116
+        143.2462961562647
+        18.48651921241045
+        31.87943551016398
+         144.066658626223
+        12.59228831600466
+        18.48934066591374
+        28.59864146766875
+        146.4719587340502
+ 2.04e+10    
+        146.1620457967622
+        29.37982720803502
+        143.7579521302964
+        18.58810608103683
+        32.06522253583282
+        144.5799288086318
+        12.62506846848179
+        18.59067416828352
+        28.81244509207384
+        147.0199297563427
+ 2.05e+10    
+        146.7034091482258
+        29.59467412042195
+        144.2683092401242
+        18.68859921137549
+        32.25078560600386
+        145.0919046202099
+        12.65604598211943
+        18.69090382848885
+        29.02548191779145
+        147.5651917183378
+ 2.06e+10    
+        147.2421398903087
+        29.80878245600465
+        144.7774126560854
+        18.78800197859537
+        32.43614042298562
+        145.6026328373844
+        12.68521553344235
+        18.79003284651923
+        29.23776829261147
+        148.1077880779528
+ 2.07e+10    
+        147.7782875388581
+        30.02217022713084
+        145.2853088230174
+        18.88631852068344
+        32.62130319755783
+        146.1121614748235
+        12.71257259813464
+        18.88806519281401
+         29.4493221309894
+        148.6477662251941
+ 2.08e+10    
+        148.3119053519593
+        30.23485695606803
+         145.792045382579
+        18.98355371761121
+        32.80629062295758
+        146.6205397046506
+        12.73811343853677
+        18.98500558774704
+        29.66016286870298
+        149.1851773604559
+ 2.09e+10    
+        148.8430501993324
+         30.4468636293101
+        146.2976710969146
+        19.07971317039323
+        32.99111984929424
+        147.1278177771855
+        12.76183509078873
+        19.08085948098757
+        29.87031141725823
+        149.7200763694377
+ 2.1e+10     
+        149.3717824288669
+         30.6582126516912
+        146.8022357737079
+        19.17480318006027
+        33.17580845840104
+        147.6340469432542
+        12.78373535163713
+        19.17563303075731
+        30.07979011809062
+        150.2525216949325
+ 2.11e+10    
+        149.8981657305732
+        30.86892780034974
+         147.305790192665
+        19.26883072656614
+        33.36037443913062
+        148.1392793781193
+        12.80381276492653
+        19.26933308300391
+        30.28862269660969
+        150.7825752057647
+ 2.12e+10    
+        150.4222669982462
+        31.07903417859828
+        147.8083860334737
+        19.36180344764919
+        33.54483616310024
+        148.6435681070634
+         12.8220666077955
+        19.36196715050902
+        30.49683421613451
+        151.3103020631457
+ 2.13e+10    
+        150.9441561891234
+        31.28855816974149
+        148.3100758052647
+        19.45372961766714
+        33.72921236089238
+        149.1469669326665
+        12.83849687659495
+        19.45354339195193
+        30.70445103176831
+        151.8357705847236
+ 2.14e+10    
+        151.4639061818319
+        31.49752739089497
+        148.8109127776158
+        19.54461812642545
+        33.91352209871604
+        149.6495303638038
+        12.85310427255081
+        19.54407059094547
+        30.91150074425626
+        152.3590521066067
+ 2.15e+10    
+        151.9815926329114
+        31.70597064684739
+         149.310950913117
+        19.63447845801699
+         34.0977847555317
+        150.1513135463974
+        12.86589018718917
+        19.63355813506466
+        31.11801215387593
+        152.8802208436475
+ 2.16e+10    
+        152.4972938322101
+        31.91391788401672
+        149.8102448015333
+        19.72332066969255
+        34.28202000064407
+        150.6523721959351
+        12.87685668754426
+        19.72201599488536
+        31.32401521440044
+        153.3993537482582
+ 2.17e+10    
+        153.0110905574338
+         32.1214001445415
+        150.3088495955755
+        19.81115537077994
+        34.46624777176522
+        151.1527625317873
+        12.88600650116882
+        19.80945470305072
+        31.52954098718402
+        153.9165303680482
+ 2.18e+10    
+        153.5230659281407
+        32.32844952055412
+        150.8068209483047
+        19.89799370166889
+        34.65048825354957
+         151.652541213327
+        12.89334300096582
+        19.89588533338345
+        31.73462159540921
+        154.4318327025619
+ 2.19e+10    
+        154.0333052594575
+        32.53509910867829
+         151.304214952182
+        19.98384731287867
+         34.8347618566025
+        152.1517652778713
+        12.89887018986118
+        19.98131948006091
+        31.93929017853999
+        154.9453450593918
+ 2.2e+10     
+        154.5418959158052
+        32.74138296479155
+        151.8010880797728
+        20.06872834422706
+        35.01908919696383
+        152.6504920804521
+        12.90259268533638
+        20.06576923686848
+        32.14358084702214
+        155.4571539099468
+ 2.21e+10    
+        155.0489271648905
+        32.94733605909565
+        152.2974971261204
+        20.15264940411304
+         35.2034910760648
+        153.1487792354148
+        12.90451570383934
+        20.14924717654976
+        32.34752863726992
+        155.9673477451446
+ 2.22e+10    
+        155.5544900322479
+        33.15299423153211
+        152.7934991527907
+        20.23562354893267
+        35.38798846116035
+        153.6466845598582
+        12.90464504509264
+        20.23176633026651
+        32.55116946697916
+        156.4760169312959
+ 2.23e+10    
+         156.058677156579
+        33.35839414758204
+        153.2891514335894
+         20.3176642626406
+         35.5726024662334
+        154.1442660189003
+        12.90298707631606
+        20.31334016718615
+        32.75454009080502
+        156.9832535664426
+ 2.24e+10    
+        156.5615826461466
+        33.56357325448599
+        153.7845114019583
+        20.39878543647245
+        35.75735433337216
+        154.6415816727823
+        12.89954871638231
+        20.39398257420917
+        32.95767805643742
+        157.4891513374035
+ 2.25e+10    
+        157.0633019364641
+        33.76856973791869
+        154.2796366000415
+        20.47900134884175
+        35.94226541461664
+        155.1386896257851
+        12.89433741992217
+        20.47370783585289
+        33.16062166111452
+        157.9938053777791
+ 2.26e+10    
+        157.5639316495256
+        33.97342247915402
+        154.7745846294199
+        20.55832664542521
+        36.12735715427281
+        155.6356479769671
+         12.8873611613965
+        20.55253061430253
+         33.3634099086027
+         158.497312127155
+ 2.27e+10    
+        158.0635694547844
+        34.17817101274863
+        155.2694131035124
+        20.63677631944826
+        36.31265107169219
+        156.1325147726967
+        12.87862841915138
+        20.63046592964607
+        33.56608246667867
+        158.9997691917362
+ 2.28e+10    
+        158.5623139321144
+        34.38285548477725
+        155.7641796016214
+        20.71436569218228
+         36.4981687445121
+        156.6293479609727
+        12.86814815947107
+        20.70752914030146
+        33.76867962514127
+        159.5012752066327
+ 2.29e+10    
+        159.0602644369538
+        34.58751661164668
+        156.2589416246262
+        20.79111039366705
+        36.68393179235485
+        157.1262053475157
+        12.85592982064649
+        20.78373592365146
+        33.97124225438611
+        160.0019297000284
+ 2.3e+10     
+        159.5575209678145
+        34.79219563951634
+        156.7537565523016
+        20.86702634366666
+        36.86996186098079
+        157.6231445536075
+        12.84198329707133
+        20.85910225689536
+        34.17381176456477
+        160.5018329594092
+ 2.31e+10    
+        160.0541840363661
+        34.99693430434955
+        157.2486816022502
+        20.94212973287012
+        37.05628060689121
+        158.1202229756616
+        12.82631892338136
+        20.93364439812888
+        34.37643006535953
+        161.0010859000763
+ 2.32e+10    
+        160.5503545402422
+        35.20177479261829
+        157.7437737904301
+         21.0164370043466
+        37.24290968237613
+        158.6174977465014
+        12.80894745865088
+        21.00737886766259
+        34.57913952639504
+        161.4997899361078
+ 2.33e+10    
+        161.0461336387474
+        35.40675970268623
+        158.2390898932612
+        21.08996483526275
+        37.42987072100328
+        159.1150256983219
+        12.78988007065808
+        21.08032242958802
+        34.78198293830991
+         161.998046853952
+ 2.34e+10    
+        161.5416226316066
+        35.61193200688503
+          158.73468641129
+        21.16273011887132
+        37.61718532354193
+        159.6128633273055
+        12.76912832023259
+        21.15249207360024
+        34.98500347450818
+        162.4959586888149
+ 2.35e+10    
+        162.0369228408978
+        35.81733501430632
+        159.2306195343872
+        21.23474994677825
+         37.8048750443162
+        160.1110667598727
+        12.74670414569688
+        21.22390499708505
+        35.18824465361161
+        162.9936276039899
+ 2.36e+10    
+         162.532135496294
+        36.02301233432433
+        159.7269451084664
+        21.30604159149509
+        37.99296137798333
+        160.6096917205322
+        12.72261984741264
+        21.29457858747956
+        35.39175030262935
+        163.4911557732737
+ 2.37e+10    
+        163.0273616237242
+        36.22900784086234
+         160.223718603684
+        21.37662248928232
+        38.18146574672928
+        161.1087935013004
+        12.69688807244193
+        21.36453040491077
+        35.59556452085877
+        163.9886452665974
+ 2.38e+10    
+        163.5227019375646
+        36.43536563741879
+        160.7209950841097
+        21.44651022329129
+        38.37040948787768
+        161.6084269326689
+        12.66952179933466
+        21.43377816512152
+        35.79973164453576
+        164.4861979389841
+ 2.39e+10    
+        164.0182567364423
+        36.64213002286137
+        161.2188291788337
+        21.51572250700663
+         38.5598138419042
+        162.1086463560738
+        12.64053432304978
+        21.50233972268693
+        36.00429621224301
+        164.9839153229501
+ 2.4e+10     
+        164.5141258027332
+        36.84934545800216
+        161.7172750544876
+        21.58427716799653
+        38.74969994085039
+        162.6095055978478
+        12.60993924002014
+        21.57023305452862
+        36.20930293108869
+        165.4818985244293
+ 2.41e+10    
+        165.0104083058239
+         37.0570565329584
+        162.2163863891475
+        21.65219213197275
+        38.94008879713139
+        163.1110579446132
+        12.57775043336856
+        21.63747624372983
+        36.41479664366547
+          165.98024812232
+ 2.42e+10    
+        165.5072027091911
+        37.26530793530865
+        162.7162163475924
+          21.719485407165
+        39.13100129272929
+         163.613356120086
+        12.54398205828215
+        21.70408746365633
+        36.62082229579633
+        166.4790640717096
+ 2.43e+10    
+        166.0046066813407
+        37.47414441904552
+        163.2168175578925
+         21.7861750690106
+        39.32245816876713
+        164.1164522632555
+        12.50864852755271
+        21.77008496238648
+        36.82742490507402
+        166.9784456108528
+ 2.44e+10    
+        166.5027170106486
+        37.68361077433427
+        163.7182420892909
+        21.85227924516404
+        39.51448001545493
+        164.6203979079044
+         12.4717644972883
+        21.83548704745336
+        37.03464953019895
+        167.4784911719389
+ 2.45e+10    
+        167.0016295241204
+         37.8937517980718
+        164.2205414313536
+        21.91781610082537
+        39.70708726240191
+        165.1252439634319
+        12.43334485280198
+        21.90031207090108
+        37.24254124111798
+           167.9792982957
+ 2.46e+10    
+        167.5014390100878
+        38.10461226525455
+        164.7237664743553
+        21.98280382439138
+        39.90030016928871
+        165.6310406969531
+        12.39340469468336
+        21.96457841465762
+        37.45114508996745
+        168.4809635498784
+ 2.47e+10    
+        168.0022391448362
+        38.31623690114702
+        165.2279674908712
+        22.04726061342697
+        40.09413881688971
+        166.1378377166244
+        12.35195932505609
+        22.02830447622571
+        37.66050608281858
+        168.9835824515779
+ 2.48e+10    
+         168.504122423177
+         38.5286703542574
+        165.7331941185417
+        22.11120466096046
+        40.28862309844167
+        166.6456839561735
+        12.30902423402703
+        22.09150865469145
+        37.87066915222752
+        169.4872493935056
+ 2.49e+10    
+        169.0071800929264
+        38.74195717010808
+        166.2394953439818
+        22.17465414209934
+        40.48377271134975
+        167.1546276605905
+        12.26461508632861
+        22.15420933705317
+        38.08167913058526
+        169.9920575741031
+ 2.5e+10     
+        169.5115020932887
+        38.95614176580468
+        166.7469194877993
+        22.23762720096793
+        40.67960714922415
+        167.6647163729438
+        12.21874770815889
+        22.21642488486881
+        38.29358072426511
+        170.4980989315578
+ 2.51e+10    
+        170.0171769970933
+        39.17126840539292
+        167.2555141906938
+        22.30014193796494
+        40.87614569423985
+        168.1759969222911
+        12.17143807422043
+        22.27817362122171
+         38.5064184885649
+        171.0054640816773
+ 2.52e+10    
+        170.5242919568651
+        39.38738117599979
+        167.7653264006069
+        22.36221639733946
+        41.07340740981437
+         168.688515412642
+        12.12270229496132
+        22.33947381800504
+        38.72023680343472
+        171.5142422595972
+ 2.53e+10    
+        171.0329326546683
+        39.60452396474996
+        168.2764023608835
+        22.42386855508373
+        41.27141113359232
+        169.2023172129425
+        12.07255660401837
+        22.40034368352202
+        38.93507984998828
+        172.0245212652902
+ 2.54e+10    
+        171.5431832556714
+        39.82274043645032
+        168.7887875994258
+        22.48511630714074
+        41.47017547073551
+        169.7174469480487
+        12.02101734586451
+         22.4608013504018
+        39.15099158778727
+         172.536387412835
+ 2.55e+10    
+        172.0551263653852
+        40.04207401203269
+        169.3025269187936
+        22.54597745792325
+        41.66971878750537
+        170.2339484906426
+        11.96810096366115
+        22.52086486382824
+        39.36801573289062
+        173.0499254833934
+ 2.56e+10    
+        172.5688429904917
+        40.26256784774463
+        169.8176643872339
+        22.60646970914228
+        41.87005920513585
+        170.7518649540745
+        11.91382398731499
+        22.58055217007932
+        39.58619573666163
+        173.5652186818427
+ 2.57e+10    
+        173.0844125032042
+        40.48426481507833
+        170.3342433306024
+        22.66661064894177
+        42.07121459398662
+        171.2712386860788
+        11.85820302173978
+        22.63988110537495
+        39.80557476531963
+        174.0823485970002
+ 2.58e+10    
+         173.601912609081
+        40.70720748142634
+        170.8523063251433
+        22.72641774133614
+        42.27320256797156
+        171.7921112633458
+        11.80125473532286
+        22.69886938503045
+        40.02619568022936
+        174.6013951653758
+ 2.59e+10    
+         174.121419318205
+        40.93143809145047
+        171.3718951911051
+        22.78590831594637
+        42.47604047925458
+        172.3145234869041
+        11.74299584859486
+        22.75753459291177
+          40.248101018913
+         175.122436638376
+ 2.6e+10     
+        174.6430069196562
+        41.15699854915334
+        171.8930509871559
+        22.84509955803212
+        42.67974541320662
+        172.8385153782889
+        11.68344312310239
+        22.81589417119001
+        40.47133297677531
+        175.6455495528835
+ 2.61e+10    
+        175.1667479591738
+        41.38393040063886
+        172.4158140055734
+        22.90400849881475
+         42.8843341836175
+        173.3641261764639
+        11.62261335048209
+        22.87396541039113
+        40.69593338952889
+        176.1708087051346
+ 2.62e+10    
+        175.6927132199328
+        41.61227481754747
+        172.9402237681775
+        22.96265200608761
+        43.08982332815553
+        173.8913943354595
+        11.56052334173424
+        22.93176543973721
+        40.92194371630544
+        176.6982871278049
+ 2.63e+10    
+        176.2209717063259
+        41.84207258115329
+        173.4663190229755
+        23.02104677510964
+          43.296229104068
+        174.4203575227027
+        11.49718991669465
+          22.989311217775
+        41.14940502344108
+        177.2280560702143
+ 2.64e+10    
+        176.7515906306602
+        42.07336406710905
+        173.9941377415015
+         23.0792093197764
+        43.50356748411784
+        174.9510526180072
+        11.43262989370218
+        23.04661952328812
+        41.37835796892068
+        177.7601849815648
+ 2.65e+10    
+         177.284635402673
+        42.30618923082248
+        174.5237171168068
+        23.13715596406577
+        43.71185415274821
+        175.4835157131921
+         11.3668600794605
+        23.10370694648825
+        41.60884278746886
+         178.294741497111
+ 2.66e+10    
+         177.820169621759
+        42.54058759345331
+        175.0550935620892
+        23.19490283375189
+        43.92110450246972
+        176.0177821122999
+        11.29989725909082
+         23.1605898804807
+        41.84089927626945
+        178.8317914271669
+ 2.67e+10    
+        178.3582550718084
+        42.77659822851118
+        175.5883027099225
+        23.25246584838474
+        44.13133363046585
+        176.5538863323952
+        11.23175818637382
+        23.21728451300017
+        42.07456678130423
+        179.3713987488557
+ 2.68e+10    
+        178.8989517185595
+        43.01425974904315
+        176.1233794120737
+         23.3098607135269
+        44.34255633540614
+        177.0918621048967
+        11.16245957417755
+        23.27380681841224
+        42.30988418429082
+        179.9136256004972
+ 2.69e+10    
+        179.4423177093542
+        43.25361029539503
+        176.6603577398637
+        23.36710291324747
+        44.55478711446676
+        177.6317423774407
+        11.09201808506917
+        23.33017254997483
+        42.54688989020805
+        180.4585322785334
+ 2.7e+10     
+         179.988409375195
+        43.49468752353035
+        177.1992709850677
+        23.42420770286355
+        44.76804016054896
+        178.1735593162275
+        11.02045032210676
+        23.38639723235628
+        42.78562181539291
+          181.00617723689
+ 2.71e+10    
+         180.537281235002
+        43.73752859389181
+         177.740151661316
+        23.48119010192705
+        44.98232935969097
+        178.7173443088426
+         10.9477728198091
+        23.44249615440363
+        43.02611737619275
+        181.5566170886735
+ 2.72e+10    
+        181.0889860019633
+        43.98217016079209
+        178.2830315059753
+        23.53806488745113
+        45.19766828866805
+        179.2631279675142
+        10.87400203529995
+        23.49848436215807
+        43.26841347815962
+        182.1099066100957
+ 2.73e+10    
+        181.6435745918793
+        44.22864836231647
+        178.8279414824904
+        23.59484658737102
+        45.41407021277434
+        179.8109401327951
+        10.79915433962367
+        23.55437665211033
+        43.51254650576979
+          182.66609874653
+ 2.74e+10    
+        182.2010961333924
+        44.47699881072354
+        179.3749117831605
+        23.65154947423454
+        45.63154808378319
+        180.3608098776365
+        10.72324600922947
+        23.61018756469332
+        43.75855231265477
+        183.2252446205906
+ 2.75e+10    
+        182.7615979800098
+        44.72725658333038
+        179.9239718323312
+        23.70818755911694
+        45.85011453807831
+        180.9127655118351
+        10.64629321762079
+        23.66593137800592
+         44.0064662123275
+        183.7873935421392
+ 2.76e+10    
+        183.3251257238085
+        44.97945621386385
+         180.475150289977
+        23.76477458575586
+        46.06978189495256
+        181.4668345868355
+        10.56831202716633
+        23.72162210176247
+        44.25632296939069
+        184.3525930201109
+ 2.77e+10    
+        183.8917232107394
+        45.23363168426812
+        181.0284750556553
+        23.82132402490057
+        46.29056215506831
+        182.0230439008572
+        10.48931838107084
+        23.77727347146492
+        44.50815679120987
+        184.9208887760686
+ 2.78e+10    
+        184.4614325574134
+        45.48981641695062
+        181.5839732728135
+        23.87784906887154
+        46.51246699907576
+        182.5814195043351
+        10.40932809550092
+        23.83289894279073
+        44.76200132004013
+         185.492324759379
+ 2.79e+10    
+        185.0342941692906
+        45.74804326745393
+        182.1416713334291
+        23.93436262632444
+         46.7355077863826
+        183.1419867056489
+        10.32835685186355
+        23.88851168619274
+        45.01788962558838
+        186.0669431639185
+ 2.8e+10     
+         185.610346760176
+        46.00834451753921
+        182.7015948829594
+        23.99087731721503
+         46.9596955540725
+        183.7047700771219
+        10.24642018923435
+        23.94412458170637
+        45.27585419799964
+        186.6447844462106
+ 2.81e+10    
+        186.1896273729274
+        46.27075186866892
+          183.26376882559
+        24.04740546795993
+        47.18504101596744
+        184.2697934612785
+        10.16353349693248
+        23.99975021395896
+        45.53592694125477
+        187.2258873449077
+ 2.82e+10    
+        186.7721714012812
+        46.53529643587213
+        183.8282173297582
+        24.10395910678765
+        47.41155456182734
+        184.8370799773279
+        10.07971200723807
+        24.05540086737644
+        45.79813916695934
+        187.8102889015127
+ 2.83e+10    
+        187.3580126127276
+        46.80200874198432
+        184.3949638339383
+         24.1605499592767
+        47.63924625668682
+        185.4066520278735
+        9.994970788251383
+        24.11108852158387
+        46.06252158852014
+        188.3980244822671
+ 2.84e+10    
+        187.9471831723317
+        47.07091871224519
+        184.9640310526651
+        24.21718944407577
+        47.86812584032025
+        185.9785313058192
+        9.909324736888387
+        24.16682484699286
+        46.32910431568709
+        188.9891278011042
+ 2.85e+10    
+        188.5397136674276
+        47.34205566924194
+        185.5354409827957
+        24.27388866880189
+        48.09820272683588
+        186.5527388014644
+        9.822788572011707
+        24.22262120057521
+        46.59791684945366
+         189.583630943592
+ 2.86e+10    
+        189.1356331331058
+        47.61544832819052
+        186.1092149099701
+        24.33065842611144
+        48.32948600439059
+        187.1292948097678
+        9.735376827693617
+         24.2784886218148
+        46.86898807730177
+        190.1815643917805
+ 2.87e+10    
+        189.7349690784204
+        47.89112479253668
+        186.6853734152788
+        24.38750918994153
+        48.56198443502544
+        187.7082189377707
+        9.647103846607717
+        24.33443782883488
+        47.14234626877691
+        190.7829570498687
+ 2.88e+10    
+        190.3377475132325
+        48.16911254987075
+        187.2639363821105
+        24.44445111191593
+        48.79570645461481
+        188.2895301121584
+        9.557983773548186
+        24.39047921469778
+        47.41801907138597
+        191.3878362706207
+ 2.89e+10    
+        190.9439929756256
+        48.44943846814107
+        187.8449230031663
+        24.50149401791273
+        49.03066017292815
+        188.8732465869539
+        9.468030549072193
+        24.44662284387031
+        47.69603350680076
+         191.996227882451
+ 2.9e+10     
+        191.5537285598284
+        48.73212879215958
+        188.4283517876327
+        24.55864740478973
+        49.26685337379992
+        189.4593859513291
+        9.377257903264921
+         24.5028784488538
+        47.97641596736266
+        192.6081562171094
+ 2.91e+10    
+        192.1669759445672
+        49.01720914038474
+        189.0142405684975
+         24.6159204372631
+        49.50429351540362
+        190.0479651375135
+        9.285679349623623
+        24.55925542697245
+        48.25919221287114
+        193.2236441378946
+ 2.92e+10    
+        192.7837554217938
+         49.3047045019749
+        189.6026065099948
+        24.67332194493694
+        49.74298773062808
+        190.6390004288074
+        9.193308179058963
+        24.61576283731776
+        48.54438736765073
+        193.8427130683261
+ 2.93e+10    
+        193.4040859257276
+         49.5946392341017
+        190.1934661151728
+        24.73086041947878
+        49.98294282755145
+        191.2325074676642
+        9.100157454011008
+         24.6724093978445
+        48.83202591788348
+        194.4653830212189
+ 2.94e+10    
+        194.0279850621462
+        49.88703705951247
+        190.7868352335623
+        24.78854401193913
+         50.2241652900104
+        191.8285012638515
+        9.006240002679061
+        24.72920348261563
+        49.12213170919764
+        195.0916726280877
+ 2.95e+10    
+        194.6554691378866
+        50.18192106433641
+        191.3827290689536
+        24.84638053021049
+        50.46666127826246
+         192.426996202674
+        8.911568413361659
+        24.78615311919092
+        49.41472794450526
+        195.7215991688311
+ 2.96e+10    
+        195.2865531904792
+        50.47931369612061
+        191.9811621872485
+        24.90437743662264
+         50.7104366297356
+        193.0280060532403
+        8.816155028906175
+        24.84326598615852
+        49.70983718207609
+        196.3551786016329
+ 2.97e+10    
+        195.9212510178874
+        50.77923676209372
+         192.582148524399
+         24.9625418456729
+        50.95549685986635
+        193.6315439767801
+        8.720011941265977
+        24.90054941080338
+        50.00748133384253
+         196.992425593031
+ 2.98e+10    
+        196.5595752082951
+         51.0817114276435
+        193.1857013944055
+        25.02088052188575
+         51.2018471630206
+         194.237622534992
+        8.623150986163131
+        24.95801036691186
+        50.30768166392454
+        197.6333535480995
+ 2.99e+10    
+        197.2015371698964
+        51.38675821500453
+        193.7918334973839
+        25.07939987780076
+        51.44949241349543
+        194.8462536984157
+        8.525583737855232
+        25.01565547270756
+        50.61045878736893
+         198.277974640698
+ 3e+10       
+        197.8471471606511
+        51.69439700214757
+        194.4005569276701
+        25.13810597208578
+        51.69843716659969
+        195.4574488548236
+        8.427321504005686
+        25.07349098891669
+        50.91583266909316
+        198.9262998437376
+ 3.01e+10    
+        198.4964143179542
+        52.00464702186237
+        195.0118831819781
+         25.1970045077717
+         51.9486856598105
+        196.0712188176244
+        8.328375320654544
+        25.13152281695986
+        51.22382262302832
+        199.5783389594284
+ 3.02e+10    
+        199.1493466882021
+        52.31752686102996
+        195.6258231675872
+        25.25610083060762
+        52.20024181400331
+        196.6875738342683
+        8.228755947290047
+        25.18975649726671
+        51.53444731145231
+        200.2341006494551
+ 3.03e+10    
+        199.8059512561965
+        52.63305446007492
+        196.2423872105552
+        25.31539992753301
+         52.4531092347537
+        197.3065235946474
+        8.128473862019154
+         25.2481972077122
+        51.84772474450758
+        200.8935924650542
+ 3.04e+10    
+        200.4662339743697
+        52.95124711259385
+        196.8615850639558
+        25.37490642526439
+        52.70729121370702
+        197.9280772394933
+        8.027539256835601
+         25.3068497621707
+        52.16367227989743
+        201.5568208769467
+ 3.05e+10    
+        201.1301997917973
+        53.27212146515293
+        197.4834259161256
+        25.43462458899531
+        52.96279073001664
+        198.5522433687547
+         7.92596203298552
+        25.36571860918632
+        52.48230662275374
+        202.2237913050994
+ 3.06e+10    
+          201.79785268296
+        53.59569351724974
+        198.1079183989187
+        25.49455832120567
+        53.21961045184506
+        199.1790300499574
+        7.823751796428342
+        25.42480783075618
+        52.80364382567093
+        202.8945081482774
+ 3.07e+10    
+        202.4691956762421
+        53.92197862143399
+        198.7350705959661
+        25.55471116058028
+        53.47775273792955
+        199.8084448265372
+        7.720917853393573
+         25.4841211412261
+        53.12769928890064
+        203.5689748133596
+ 3.08e+10    
+        203.1442308821326
+        54.25099148358105
+         199.364890050928
+        25.61508628103258
+        53.73721963920691
+        200.4404947261443
+        7.617469206031686
+        25.54366188629421
+        53.45448776070011
+        204.2471937443897
+ 3.09e+10    
+         203.822959521109
+         54.5827461633164
+        199.9973837757358
+        25.67568649083375
+        53.99801290049876
+        201.0751862689155
+         7.51341454815908
+         25.6034330421221
+        53.78402333783421
+        204.9291664513433
+ 3.1e+10     
+        204.5053819511816
+        54.91725607458272
+        200.6325582588211
+        25.73651423184316
+        54.26013396225218
+        201.7125254757034
+        7.408762261096147
+         25.6634372145513
+        54.11631946621964
+        205.6148935385698
+ 3.11e+10    
+        205.1914976950813
+        55.25453398634828
+        201.2704194733255
+        25.79757157883995
+        54.52358396233639
+        202.3525178762656
+        7.303520409598278
+        25.72367663842212
+        54.45138894171158
+        206.3043747329107
+ 3.12e+10    
+        205.8813054670723
+        55.59459202345021
+        201.9109728852846
+        25.85886023895327
+        54.78836373789358
+        202.9951685174095
+         7.19769673787907
+        25.78415317699438
+        54.78924391102738
+        206.9976089114504
+ 3.13e+10    
+        206.5748031993738
+        55.93744166757373
+         202.554223461791
+        25.92038155119002
+        55.05447382724029
+        203.6404819710862
+        7.091298665725985
+        25.84486832146764
+        55.12989587280284
+        207.6945941289057
+ 3.14e+10    
+        207.2719880681776
+        56.28309375835538
+        203.2001756791142
+        25.98213648605801
+        55.32191447182005
+        204.2884623424321
+        6.984333284707219
+        25.90582319059865
+        55.47335567877674
+        208.3953276446129
+ 3.15e+10    
+        207.9728565192477
+         56.6315584946156
+        203.8488335307997
+         26.0441256452833
+        55.59068561820472
+        204.9391132777578
+        6.876807354470632
+        25.96701853041576
+        55.81963353510229
+        209.0998059491167
+ 3.16e+10    
+        208.6774042930875
+        56.98284543571083
+        204.5002005357118
+        26.10634926162051
+        55.86078692014195
+        205.5924379724757
+        6.768727299133873
+        26.02845471402764
+        56.16873900377992
+        209.8080247903402
+ 3.17e+10    
+         209.385626449678
+        57.33696350300804
+        205.1542797460562
+        26.16880719875423
+        56.13221774065008
+        206.2484391789716
+        6.660099203765817
+        26.09013174152491
+        56.52068100420759
+        210.5199791993164
+ 3.18e+10    
+        210.0975173927608
+        57.69392098147236
+        205.8110737553381
+        26.23149895129077
+        56.40497715415616
+        206.9071192144142
+        6.550928810959572
+        26.15204923997441
+        56.87546781485055
+        211.2356635154897
+ 3.19e+10    
+        210.8130708936655
+         58.0537255213704
+        206.4705847062878
+        26.29442364483833
+        56.67906394867766
+        207.5684799684973
+        6.441221517496619
+        26.21420646350301
+        57.23310707502008
+        211.9550714115562
+ 3.2e+10     
+        211.5322801146872
+        58.41638414008447
+        207.1328142987259
+        26.35758003617529
+        56.95447662804566
+        208.2325229111195
+          6.3309823711025
+        26.27660229347094
+        57.59360578676628
+        212.6781959178532
+ 3.21e+10    
+        212.2551376319856
+        58.78190322403481
+        207.7977637973844
+        26.42096651350463
+        57.23121341416868
+         208.899249099997
+         6.22021606729411
+        26.33923523873302
+         57.9569703168762
+        213.4050294462786
+ 3.22e+10    
+        212.9816354580268
+        59.15028853071148
+         208.465434039671
+         26.4845810967937
+        57.50927224933571
+        209.5686591882074
+        6.108926946318755
+        26.40210343598667
+        58.32320639897974
+        214.1355638137405
+ 3.23e+10    
+        213.7117650635437
+        59.52154519080656
+        209.1358254433751
+        26.54842143819846
+        57.78865079855695
+        210.2407534316618
+        5.997118990185371
+        26.46520465020541
+        58.69231913575793
+        214.8697902651368
+ 3.24e+10    
+        214.4455173990289
+        59.89567771045232
+        209.8089380143196
+         26.6124848225715
+        58.06934645194302
+        210.9155316965115
+        5.884795819787815
+        26.52853627515707
+        59.06431300125392
+        215.6076994958493
+ 3.25e+10    
+        215.1828829157484
+        60.27268997355941
+        210.4847713539528
+        26.67676816805118
+        58.35135632711754
+        211.5929934664767
+        5.771960692120912
+        26.59209533400512
+        59.43919184328207
+        216.3492816737596
+ 3.26e+10    
+        215.9238515862853
+        60.65258524425429
+        211.1633246668788
+        26.74126802673382
+        58.63467727166726
+        212.2731378501085
+        5.658616497589543
+        26.65587847999305
+        59.81695888593649
+        217.0945264607857
+ 3.27e+10    
+        216.6684129246013
+        61.03536616941363
+        211.8445967683265
+        26.80598058542522
+        58.91930586562389
+        212.9559635879748
+          5.5447657574109
+        26.71988199720973
+        60.19761673219539
+         217.843423033933
+ 3.28e+10    
+        217.4165560056326
+        61.42103478129631
+        212.5285860915546
+        26.87090166647297
+        59.20523842398008
+        213.6414690597764
+        5.430410621110926
+        26.78410180143599
+         60.5811673666198
+        218.5959601058625
+ 3.29e+10    
+        218.1682694844107
+        61.80959250026891
+        213.2152906951964
+         26.9360267286766
+        59.49247099923645
+        214.3296522913839
+        5.315552864114354
+        26.84853344107045
+        60.96761215814611
+        219.3521259449775
+ 3.3e+10     
+        218.9235416147143
+        62.20104013762505
+        213.9047082705322
+        27.00135086827687
+        59.78099938397975
+        215.0205109618067
+        5.200193885430227
+         26.9131720981348
+        61.35695186297093
+         220.111908395034
+ 3.31e+10    
+         219.682360267259
+        62.59537789849811
+         214.596836148708
+         27.0668688200222
+        60.07081911349158
+        215.7140424100839
+        5.084334705432273
+        26.97801258935718
+        61.74918662752643
+        220.8752948942694
+ 3.32e+10    
+        220.4447129474216
+        62.99260538486276
+        215.2916713078744
+        27.13257495831147
+        60.36192546838614
+        216.4102436421039
+        4.967975963735032
+        27.04304936733256
+        62.14431599154437
+        221.6422724940584
+ 3.33e+10    
+        221.2105868125089
+        63.39272159862919
+        215.9892103802688
+        27.19846329841361
+        60.65431347727493
+        217.1091113373483
+        4.851117917166476
+        27.10827652176008
+        62.54233889121086
+        222.4128278770996
+ 3.34e+10    
+        221.9799686885765
+        63.79572494482549
+        216.6894496592303
+        27.26452749776191
+        60.94797791946188
+        217.8106418555625
+        4.733760437837763
+        27.17368778075702
+        62.94325366240752
+        223.1869473751348
+ 3.35e+10    
+         222.752845086796
+        64.20161323486681
+        217.3923851061382
+        27.33076085732322
+        61.24291332766209
+        218.5148312433533
+        4.615903011309815
+        27.23927651224638
+        63.34705804403819
+        223.9646169862017
+ 3.36e+10    
+        223.5292022193831
+        64.61038368991417
+        218.0980123572947
+        27.39715632304172
+        61.53911399074889
+        219.2216752407126
+        4.497544734859034
+        27.30503572542094
+        63.75374918144364
+        224.7458223914394
+ 3.37e+10    
+        224.3090260150904
+        65.02203294431868
+        218.8063267307322
+        27.46370648735571
+        61.83657395652521
+        219.9311692874683
+         4.37868431584109
+        27.37095807228049
+        64.16332362990052
+        225.5305489714337
+ 3.38e+10    
+        225.0923021342705
+        65.43655704915125
+        219.5173232329547
+        27.53040359078779
+        62.13528703451924
+        220.6433085296629
+        4.259320070154239
+         27.4370358492421
+        64.57577735820311
+        226.3187818221206
+ 3.39e+10    
+        225.8790159835122
+        65.85395147581778
+        220.2309965656153
+        27.59723952360698
+          62.435246798805
+        221.3580878258608
+        4.139449920803045
+        27.50326099882398
+        64.99110575233121
+        227.1105057702517
+ 3.4e+10     
+        226.6691527298714
+        66.27421111975929
+        220.9473411321206
+        27.66420582756335
+         62.7364465908451
+        222.0755017533841
+        4.019071396562547
+        27.56962511140113
+        65.40930361919924
+         227.905705388423
+ 3.41e+10    
+        227.4626973146772
+        66.69733030423383
+        221.6663510441716
+         27.7312936976934
+        63.03887952235664
+        222.7955446144771
+        3.898181630743904
+        27.63611942703288
+        65.83036519048713
+        228.7043650096814
+ 3.42e+10    
+         228.259634466953
+        67.12330278418358
+        222.3880201282338
+        27.79849398419656
+        63.34253847819878
+        223.5182104423992
+        3.776777360062225
+        27.70273483736108
+        66.25428412655491
+        229.5064687417102
+ 3.43e+10    
+        229.0599487164303
+        67.55212175018417
+        223.1123419319487
+        27.86579719438225
+        63.64741611928185
+        224.2434930074545
+        3.654854923607189
+        27.76946188757983
+        66.68105352043654
+        230.3120004806049
+ 3.44e+10    
+        229.8636244061837
+        67.98377983247447
+        223.8393097304692
+        27.93319349468614
+        63.95350488549717
+        224.9713858229458
+        3.532410261917029
+        27.83629077847471
+        67.11066590191624
+         231.120943924244
+ 3.45e+10    
+        230.6706457048847
+        68.41826910506953
+        224.5689165327331
+        28.00067271275643
+        64.26079699866668
+        225.7018821510638
+         3.40943891615677
+        27.90321136853135
+        67.54311324168191
+        231.9332825852604
+ 3.46e+10    
+         231.480996618681
+        68.85558108995298
+         225.301155087674
+        28.06822433960876
+        64.56928446551302
+        226.4349750087117
+        3.285936027401329
+        27.97021317611384
+        67.97838695556214
+        232.7489998036293
+ 3.47e+10    
+        232.2946610027177
+        69.29570676135134
+        226.0360178903628
+        28.13583753184923
+        64.87895908064722
+        227.1706571732587
+        3.161896336024016
+        28.03728538171118
+        68.41647790883916
+        233.5680787588711
+ 3.48e+10    
+        233.1116225723044
+        69.73863655008707
+        226.7734971880872
+        28.20350111396616
+        65.18981242957682
+        227.9089211882351
+        3.037314181191803
+        28.10441683025266
+        68.85737642064316
+        234.3905024818891
+ 3.49e+10    
+        233.9318649137276
+        70.18436034801175
+        227.5135849863671
+        28.27120358068845
+        65.50183589173059
+        228.6497593689543
+        2.912183500466542
+        28.17159603348979
+        69.30107226842192
+        235.2162538664269
+ 3.5e+10     
+        234.7553714947308
+        70.63286751251755
+        228.2562730549057
+        28.33893309941167
+        65.81502064350062
+        229.3931638080804
+         2.78649782951468
+        28.23881117244629
+        69.74755469249071
+        236.0453156801865
+ 3.51e+10    
+        235.5821256746613
+        71.08414687112807
+        229.0015529334795
+        28.40667751269034
+         66.1293576613029
+        230.1391263811274
+        2.660250301925096
+        28.30605009993501
+        70.19681240065978
+        236.8776705755896
+ 3.52e+10    
+        236.4121107142961
+         71.5381867261668
+        229.7494159377673
+        28.47442434079696
+        66.44483772465334
+        230.8876387519023
+        2.533433649135358
+        28.37330034314044
+        70.64883357293742
+        237.7133011001987
+ 3.53e+10    
+        237.2453097853504
+        71.99497485950289
+         230.499853165114
+        28.54216078434599
+        66.76145141925961
+        231.6386923778808
+        2.406040200468308
+        28.44054910626787
+        71.10360586631037
+        238.5521897068086
+ 3.54e+10    
+        238.0817059796778
+        72.45449853737442
+        231.2528555002379
+        28.60987372698358
+        67.07918914012951
+         232.392278515529
+         2.27806188327836
+        28.50778327325738
+        71.56111641960069
+        239.3943187632131
+ 3.55e+10    
+        238.9212823181813
+        72.91674451528912
+        232.0084136208774
+        28.67754973814229
+         67.3980410946937
+        233.1483882255664
+        2.149490223209143
+        28.57498941056324
+        72.02135185839899
+        240.2396705616568
+ 3.56e+10    
+        239.7640217594194
+        73.38169904299889
+        232.7665180033788
+        28.74517507585988
+        67.71799730594446
+        233.9070123781706
+         2.02031634456231
+         28.6421537699978
+        72.48429830007157
+        241.0882273279791
+ 3.57e+10    
+        240.6099072079444
+        73.84934786955371
+        233.5271589282268
+         28.8127356896623
+        68.03904761558645
+        234.6681416581213
+        1.890530970778909
+        28.70926229163909
+        72.94994135884413
+        241.9399712304605
+ 3.58e+10    
+        241.4589215223529
+        74.31967624842753
+         234.290326485513
+         28.8802172235103
+        68.36118168720461
+        235.4317665699002
+        1.760124425033148
+         28.7763006068031
+        73.41826615095961
+        242.7948843883761
+ 3.59e+10    
+         242.311047523078
+        74.79266894272098
+         235.056010580357
+        28.94760501880862
+        68.68438900944203
+        236.1978774427238
+        1.629086630939897
+        28.84325404107808
+        73.88925729991024
+        243.6529488802678
+ 3.6e+10     
+        243.1662679999167
+        75.26831023043667
+        235.8242009382626
+        29.01488411747864
+        69.00865889919375
+        236.9664644355297
+        1.497407113375966
+         28.9101076174224
+        74.36289894174257
+        244.5141467519391
+ 3.61e+10    
+        244.0245657193129
+        75.74658390983198
+        236.5948871104263
+        29.08203926509281
+        69.33398050481189
+        237.7375175419131
+        1.365074999416032
+        28.97684605932457
+        74.83917473043809
+        245.3784600241868
+ 3.62e+10    
+        244.8859234313844
+        76.22747330483944
+        237.3680584789856
+        29.14905491407056
+        69.66034280932314
+        238.5110265950047
+        1.232079019383531
+        29.04345379402529
+        75.31806784336371
+        246.2458707002697
+ 3.63e+10    
+        245.7503238767235
+        76.71096127056539
+        238.1437042622208
+        29.21591522693617
+        69.98773463365902
+        239.2869812723043
+        1.098407508017299
+         29.1099149558007
+        75.79956098679729
+        247.1163607731256
+ 3.64e+10    
+        246.6177497929641
+        77.19703019885746
+        238.9218135197004
+        29.28260407963708
+        70.31614463989663
+        240.0653711004628
+       0.9640484057543324
+        29.17621338930668
+        76.28363640152261
+        247.9899122323465
+ 3.65e+10    
+        247.4881839211273
+        77.68566202394602
+        239.7023751573752
+        29.34910506492258
+        70.64556133451117
+        240.8461854600167
+       0.8289892601294016
+         29.2423326529843
+        76.77027586849952
+        248.8665070709181
+ 3.66e+10    
+        248.3616090117484
+        78.17683822815465
+        240.4853779326223
+        29.41540149578286
+         70.9759730716394
+        241.6294135900754
+       0.6932172272913784
+        29.30825602252418
+        77.25946071459998
+        249.7461272917246
+ 3.67e+10    
+        249.2380078308007
+        78.67053984768333
+        241.2708104592431
+        29.48147640894709
+        71.30736805635372
+        242.4150445929613
+       0.5567190736377787
+        29.37396649439157
+        77.75117181841867
+        250.6287549138366
+ 3.68e+10    
+        250.1173631654144
+         79.1667474784598
+        242.0586612124061
+        29.54731256844046
+        71.63973434794548
+        243.2030674388056
+        0.419481177566885
+         29.4394467894104
+        78.24538961615251
+        251.5143719785839
+ 3.69e+10    
+        250.9996578294005
+        79.66544128206218
+         242.848918533546
+        29.61289246920023
+        71.97305986321908
+         243.993470970101
+       0.2814895313485684
+        29.50467935640516
+        78.74209410754705
+        252.4029605554155
+ 3.7e+10     
+        251.8848746685894
+        80.16660099170836
+        243.6415706352159
+        29.67819834074952
+        72.30733237979534
+        244.7862439062084
+       0.1427297431142236
+        29.56964637590215
+        79.24126486191494
+        253.2945027475643
+ 3.71e+10    
+        252.7729965659834
+         80.6702059183157
+        244.4366056058909
+        29.74321215092838
+        72.64253953942359
+        245.5813748478234
+     0.003187038965702271
+         29.6343297638878
+        79.74288102422125
+        254.1889806975168
+ 3.72e+10    
+         253.664006446736
+        81.17623495662616
+        245.2340114147272
+         29.8079156096825
+        72.97866885130276
+        246.3788522813998
+      -0.1371537347959082
+        29.69871117562425
+        80.24692132123504
+        255.0863765922886
+ 3.73e+10    
+        254.5578872829647
+         81.6846665913999
+        246.0337759162784
+         29.8722901729079
+        73.31570769541131
+        247.1786645835348
+      -0.2783081093215802
+        29.76277200952182
+        80.75336406774952
+        255.9866726685289
+ 3.74e+10    
+        255.4546220983909
+        82.19547890367436
+        246.8358868551669
+        29.93631704635222
+        73.65364332584463
+        247.9808000253126
+      -0.4202919907450156
+        29.82649341106786
+        81.26218717286832
+        256.8898512174397
+ 3.75e+10    
+        256.3541939728349
+        82.70864957708868
+        247.6403318707097
+        29.99997718957069
+         73.9924628741604
+        248.7852467766082
+      -0.5631216575928901
+        29.88985627681084
+        81.77336814635647
+         257.795894589538
+ 3.76e+10    
+        257.2565860465498
+        83.22415590427238
+        248.4470985015065
+        30.06325131993827
+        74.33215335273232
+        249.5919929103591
+      -0.7068137580745173
+        29.95284125839998
+        82.28688410505667
+        258.7047851992403
+ 3.77e+10    
+        258.1617815244118
+        83.74197479330059
+        249.2561741899825
+        30.12611991671533
+        74.67270165810989
+        250.4010264067919
+      -0.8513853072492719
+        30.01542876667962
+        82.80271177936999
+        259.6165055293044
+ 3.78e+10    
+          259.06976367997
+        84.26208277420815
+        250.0675462868972
+        30.18856322516737
+        75.01409457438538
+        251.2123351576187
+      -0.9968536840738276
+        30.07759897583774
+        83.32082751980016
+        260.5310381351134
+ 3.79e+10    
+        259.9805158593617
+        84.78445600557086
+        250.8812020558036
+        30.25056126073877
+        75.35631877656789
+        252.0259069701977
+       -1.143236628326821
+         30.1393318276077
+        83.84120730356004
+        261.4483656488133
+ 3.8e+10     
+        260.8940214850978
+        85.30907028114412
+        251.6971286774755
+        30.31209381327848
+         75.6993608339629
+         252.841729571654
+       -1.290552237412308
+        30.20060703552366
+        84.36382674124066
+        262.3684707833159
+ 3.81e+10    
+        261.8102640597182
+        85.83590103656609
+        252.5153132542966
+        30.37314045131887
+        76.04320721355857
+        253.6597906129757
+       -1.438818963040876
+        30.26140408922815
+        84.88866108354071
+        263.2913363361609
+ 3.82e+10    
+        262.7292271693336
+        86.36492335611875
+        253.3357428146075
+        30.43368052640547
+        76.38784428341654
+        254.4800776730666
+       -1.588055607788925
+        30.32170225883133
+         85.4156852280575
+        264.2169451932511
+ 3.83e+10    
+        263.6508944870468
+        86.89611197954791
+        254.1584043170206
+        30.49369317747879
+        76.73325831607022
+        255.3025782627774
+       -1.738281321535506
+        30.38148059932276
+        85.94487372613719
+        265.1452803324698
+ 3.84e+10    
+        264.5752497762693
+        87.42944130894402
+        254.9832846546965
+        30.55315733530562
+        77.07943549192478
+        256.1272798288962
+       -1.889515597777094
+        30.44071795503243
+        86.47620078978245
+        266.0763248271642
+ 3.85e+10    
+        265.5022768939213
+        87.96488541567732
+        255.8103706595854
+        30.61205172696113
+        77.42636190266546
+        256.9541697581149
+       -2.041778269819942
+         30.4993929641434
+        87.00964029862078
+        267.0100618495309
+ 3.86e+10    
+        266.4319597935385
+        88.50241804739123
+        256.6396491066334
+        30.67035488036021
+        77.77402355466795
+        257.7832353809598
+       -2.195089506850101
+         30.5574840632532
+        87.54516580692652
+         267.946474673876
+ 3.87e+10    
+        267.3642825282823
+        89.04201263505172
+         257.471106717958
+        30.72804512883713
+        78.12240637241347
+        258.6144639756992
+       -2.349469809880933
+        30.61496949198494
+        88.08275055070231
+        268.8855466797841
+ 3.88e+10    
+        268.2992292538447
+        89.58364230005039
+        258.3047301669836
+        30.78510061577412
+        78.47149620190901
+        259.4478427722192
+       -2.504940007578743
+         30.6718272976462
+        88.62236745481326
+        269.8272613551741
+ 3.89e+10    
+        269.2367842312797
+        90.12727986136245
+        259.1405060825533
+        30.84149929927662
+        78.82127881410858
+        260.2833589558673
+       -2.661521251965587
+        30.72803533993646
+        89.16398914017665
+        270.7716022992678
+ 3.9e+10     
+        270.1769318297352
+        90.67289784275562
+        259.9784210529987
+        30.89721895689615
+        79.17173990834013
+        261.1209996712769
+       -2.819235014000419
+        30.78357129570112
+        89.70758793100504
+        271.7185532254561
+ 3.91e+10    
+        271.1196565291111
+        91.22046848005334
+        260.8184616301888
+        30.95223719039924
+        79.52286511573499
+        261.9607520261615
+       -2.978103079037688
+        30.83841266373269
+        90.25313586210186
+        272.6680979640882
+ 3.92e+10    
+        272.0649429226376
+        91.76996372844772
+         261.660614333537
+        31.00653143058184
+        79.87464000265794
+        262.8026030950769
+       -3.138147542164607
+        30.89253676961741
+        90.80060468620746
+        273.6202204651652
+ 3.93e+10    
+        273.0127757193749
+        92.32135526986113
+        262.5048656539886
+        31.06007894212894
+        80.22705007414335
+        263.6465399231694
+       -3.299390803416237
+        30.94592077062766
+        91.34996588139691
+        274.5749048009588
+ 3.94e+10    
+         273.963139746647
+        92.87461452035872
+        263.3512020579691
+         31.1128568285184
+         80.5800807773298
+        264.4925495298875
+       -3.461855562869277
+        30.99854166065854
+        91.90119065852656
+        275.5321351685519
+ 3.95e+10    
+        274.9160199524019
+        93.42971263760799
+        264.1996099913123
+         31.1648420369685
+        80.93371750489922
+        265.3406189126781
+       -3.625564815614458
+        31.05037627520896
+        92.45424996872951
+        276.4918958923012
+ 3.96e+10    
+        275.8714014075124
+        93.98662052838476
+         265.050075883152
+        31.21601136342849
+        81.28794559851623
+        266.1907350506529
+       -3.790541846608002
+        31.10140129640559
+        93.00911451095772
+        277.4541714262367
+ 3.97e+10    
+        276.8292693080115
+        94.54530885612488
+        265.9025861497897
+        31.26634145761132
+        81.64275035226846
+        267.0428849082334
+         -3.9568102254023
+        31.15159325806999
+         93.5657547395718
+        278.4189463563867
+ 3.98e+10    
+        277.7896089772681
+        95.10574804852085
+         266.757127198535
+        31.31580882806838
+        81.99811701610982
+         267.897055438774
+       -4.124393800756342
+        31.20092855082707
+        94.12414087197436
+        279.3862054030428
+ 3.99e+10    
+        278.7524058681083
+        95.66790830516223
+        267.6136854315187
+        31.36438984730465
+        82.35403079930191
+        268.7532335881592
+       -4.293316695125861
+         31.2493834272555
+        94.68424289628908
+        280.3559334229629
+ 4e+10       
+        279.7176455648845
+        96.23175960521799
+        268.4722472494768
+        31.41206075693428
+        82.71047687385739
+        269.6114062983857
+       -4.463603299033992
+        31.29693400707836
+        95.24603057908251
+        281.3281154115156
+ 4.01e+10    
+        280.6853137854935
+        96.79727171516086
+        269.3327990555111
+        31.45879767287617
+        83.06744037798359
+        270.4715605111139
+       -4.635278265322779
+        31.34355628239339
+        95.80947347312784
+        282.3027365047694
+ 4.02e+10    
+        281.6553963833408
+        97.36441419653106
+         270.195327258826
+        31.50457659058735
+         83.4249064195248
+        271.3336831712036
+       -4.808366503285886
+        31.38922612294318
+        96.37454092520824
+        283.2797819815297
+ 4.03e+10    
+        282.6278793492653
+        97.93315641373938
+        271.0598182784329
+         31.5493733903355
+        83.78286007940557
+         272.197761230232
+       -4.982893172682729
+        31.43391928142318
+        96.94120208396342
+         284.259237265327
+ 4.04e+10    
+        283.6027488134224
+        98.50346754190888
+        271.9262585468386
+         31.5931638425078
+        84.14128641507226
+        273.0637816499806
+       -5.158883677635387
+         31.4776113988273
+        97.50942590777039
+        285.2410879263538
+ 4.05e+10    
+        284.5799910471187
+        99.07531657475303
+        272.7946345137042
+        31.63592361295747
+        84.50017046393388
+        273.9317314059149
+       -5.336363660407754
+         31.5202780098315
+        98.07918117266583
+        286.2253196833639
+ 4.06e+10    
+        285.5595924646113
+        99.64867233248886
+        273.6649326494804
+        31.67762826838504
+        84.85949724680162
+        274.8015974906365
+       -5.515358995068477
+        31.56189454821229
+        98.65043648030209
+        287.2119184055175
+ 4.07e+10    
+        286.5415396248732
+         100.223503469786
+        274.5371394490231
+        31.71825328175563
+        85.21925177132765
+        275.6733669173153
+       -5.695895781037778
+        31.60243635230162
+        99.22316026593901
+        288.2008701142011
+ 4.08e+10    
+        287.5258192333187
+        100.7997784837464
+         275.411241435176
+        31.75777403775012
+        85.57941903544018
+        276.5470267231128
+        -5.87800033651858
+        31.64187867047614
+        99.79732080647052
+        289.1921609847916
+ 4.09e+10    
+        288.5124181434983
+          101.37746572192
+        276.2872251623464
+         31.7961658382498
+        85.93998403077855
+        277.4225639725703
+       -6.061699191813548
+        31.68019666668073
+        100.3728862284828
+        290.1857773484019
+ 4.1e+10     
+        289.5013233587636
+        101.9565333903484
+         277.165077220044
+        31.83340390785435
+        86.30093174612468
+        278.2999657609947
+       -6.247019082527514
+        31.71736542598488
+        100.9498245163457
+        291.1817056935792
+ 4.11e+10    
+        290.4925220338994
+        102.5369495616371
+        278.0447842363994
+        31.86946339943088
+        86.66224717083145
+        279.1792192178162
+       -6.433986942657428
+        31.75335996017147
+        101.5281035203313
+        292.1799326679761
+ 4.12e+10    
+        291.4860014767308
+        103.1186821830618
+        278.9263328816751
+         31.9043193996954
+        87.02391529824992
+        280.0603115099325
+       -6.622629897569087
+        31.78815521335759
+        102.1076909647662
+        293.1804450799909
+ 4.13e+10    
+        292.4817491497039
+        103.7016990846948
+        279.8097098717309
+        31.93794693482376
+        87.38592112915117
+        280.9432298450349
+       -6.812975256862811
+        31.82172606764588
+         102.688554456208
+          294.18322990038
+ 4.14e+10    
+        293.4797526714408
+        104.2859679875632
+        280.6949019714926
+        31.97032097609256
+        87.74824967514616
+        281.8279614749151
+       -7.005050507128145
+        31.85404734880571
+        103.2706614916492
+        295.1882742638395
+ 4.15e+10    
+        294.4799998182721
+        104.8714565118284
+        281.5818959983814
+        32.00141644554914
+        88.11088596210128
+        282.7144936987606
+       -7.198883304588668
+        31.88509383198441
+        103.8539794667489
+        296.1955654705677
+ 4.16e+10    
+        295.4824785257464
+        105.4581321849908
+        282.4706788257321
+         32.0312082217089
+        88.47381503354936
+         283.602813866422
+       -7.394501467637919
+        31.91484024744578
+        104.4384756840842
+        297.2050909877946
+ 4.17e+10    
+        296.4871768901225
+        106.0459624501162
+        283.3612373861884
+         32.0596711452805
+        88.83702195409698
+         284.492909381678
+       -7.591932969267089
+        31.94326128633711
+        105.0241173614302
+        298.2168384512979
+ 4.18e+10    
+        297.4940831698379
+        106.6349146740839
+        284.2535586750782
+        32.08678002491717
+        89.20049181282729
+        285.3847677054756
+       -7.791205929386247
+         31.9703316064826
+        105.6108716400561
+         299.230795666892
+ 4.19e+10    
+        298.5031857869625
+        107.2249561558534
+        285.1476297537649
+        32.11250964299333
+        89.56420972669697
+        286.2783763591513
+       -7.992348607038694
+        31.99602583820261
+        106.1987055930456
+        300.2469506118981
+ 4.2e+10     
+        299.5144733286336
+        107.8160541347509
+        286.0434377529903
+        32.13683476140606
+        89.92816084392891
+        287.1737229276444
+       -8.195389392511256
+        32.02031859015845
+        106.7875862336345
+        301.2652914365962
+ 4.21e+10    
+        300.5279345484777
+        108.4081757987729
+        286.9409698761834
+        32.15973012740085
+        90.29233034739927
+        288.0707950626897
+       -8.400356799340134
+        32.04318445522082
+        107.3774805235671
+        302.2858064656588
+ 4.22e+10    
+        301.5435583680118
+        109.0012882929045
+        287.8402134027583
+        32.18117047941906
+        90.65670345801804
+        288.9695804859916
+       -8.607279456214268
+         32.0645980163624
+        107.9683553814685
+        303.3084841995719
+ 4.23e+10    
+         302.561333878039
+        109.5953587274545
+        288.7411556913949
+        32.20113055296939
+         91.0212654381049
+        289.8700669923919
+       -8.816186098777104
+        32.08453385257215
+        108.5601776912326
+        304.3333133160303
+ 4.24e+10    
+        303.5812503400218
+        110.1903541864017
+        289.6437841832906
+        32.21958508651881
+        91.38600159475733
+        290.7722424530109
+       -9.027105561327861
+        32.10296654479198
+        109.1529143104241
+        305.3602826713341
+ 4.25e+10    
+        304.6032971874527
+        110.7862417357561
+        290.5480864054064
+        32.23650882740506
+        91.75089728321346
+         291.676094818379
+       -9.240066768424006
+         32.1198706818741
+        109.7465320786924
+        306.3893813017543
+ 4.26e+10    
+        305.6274640272027
+        111.3829884319291
+        291.4540499736837
+        32.25187653776828
+        92.11593791020724
+        292.5816121215548
+       -9.455098726385268
+        32.13522086655789
+        110.3409978261987
+        307.4205984249012
+ 4.27e+10    
+        306.6537406408721
+        111.9805613301122
+         292.361662596245
+        32.26566300050125
+        92.48110893731638
+        293.4887824812251
+       -9.672230514701649
+        32.14899172146673
+        110.9362783820519
+        308.4539234410706
+ 4.28e+10    
+        307.6821169861172
+        112.5789274926686
+        293.2709120765817
+        32.27784302521729
+        92.84639588430382
+        294.3975941047838
+       -9.891491277345917
+        32.16115789512182
+         111.532340582752
+        309.4893459345812
+ 4.29e+10    
+          308.71258319798
+        113.1780539975263
+        294.1817863167155
+        32.28839145423592
+        93.21178433245099
+        295.3080352914124
+       -10.11291021399212
+        32.17169406797436
+        112.1291512806444
+        310.5268556751047
+ 4.3e+10     
+        309.7451295902006
+        113.7779079465808
+        295.0942733203474
+        32.29728316858291
+        93.57725992788193
+        296.2200944351254
+       -10.33651657114205
+        32.18057495845372
+        112.7266773523778
+        311.5664426189853
+ 4.31e+10    
+         310.779746656525
+        114.3784564741019
+        296.0083611959864
+        32.30449309400701
+        93.94280838488173
+        297.1337600278156
+       -10.56233963315992
+        32.18777532903101
+        113.3248857073681
+        312.6080969105445
+ 4.32e+10    
+         311.816425072006
+         114.979666755141
+        296.9240381600594
+        32.30999620700992
+        94.30841548920448
+        298.0490206622783
+       -10.79040871321836
+        32.19326999229752
+        113.9237432962657
+        313.6518088833889
+ 4.33e+10    
+        312.8551556942972
+        115.5815060139447
+        297.8412925400041
+        32.31376754088995
+        94.67406710137247
+        298.9658650352184
+       -11.02075314415568
+        32.19703381705645
+        114.5232171194243
+        314.6975690616949
+ 4.34e+10    
+        313.8959295649339
+         116.183941532365
+        298.7601127773466
+        32.31578219179771
+        95.03974915996832
+        299.8842819502501
+       -11.25340226924702
+        32.19904173442822
+        115.1232742353728
+        315.7453681614997
+ 4.35e+10    
+        314.9387379106157
+        116.7869406582716
+        299.6804874307547
+        32.31601532480389
+        95.40544768491463
+        300.8042603208737
+       -11.48838543289034
+        32.19926874396618
+        115.7238817692837
+        316.7951970919776
+ 4.36e+10    
+        315.9835721444832
+        117.3904708139619
+        300.6024051790825
+        32.31444217997684
+        95.77114878074757
+        301.7257891734428
+       -11.72573197120905
+        32.19768991978539
+        116.3250069214448
+        317.8470469567111
+ 4.37e+10    
+        317.0304238673768
+        117.9944995045655
+        301.5258548243858
+        32.31103807847018
+        96.13683863987738
+        302.6488576501135
+       -11.96547120257309
+        32.19428041669941
+        116.9266169757221
+        318.9009090549578
+ 4.38e+10    
+        318.0792848691078
+        118.5989943264484
+        302.4508252949336
+        32.30577842861914
+        96.50250354584131
+        303.5734550117804
+       -12.20763241804012
+        32.18901547636722
+        117.5286793080233
+        319.9567748829085
+ 4.39e+10    
+        319.1301471297105
+        119.2039229756079
+         303.377305648188
+        32.29863873204455
+        96.86812987654473
+        304.4995706409993
+       -12.45224487171809
+        32.18187043344822
+        118.1311613947545
+        321.0146361349408
+ 4.4e+10     
+        320.1830028206982
+        119.8092532560622
+        304.3052850737774
+        32.28959458976337
+        97.23370410749146
+        305.4271940448895
+       -12.69933777105137
+         32.1728207217641
+        118.7340308212679
+        322.0744847048693
+ 4.41e+10    
+        321.2378443063054
+        120.4149530882318
+        305.2347528964477
+        32.27862170830589
+        97.59921281500469
+        306.3563148580277
+       -12.94894026703236
+        32.16184188046734
+        119.3372552903051
+        323.1363126871851
+ 4.42e+10    
+        322.2946641447348
+        121.0209905173113
+         306.165698578994
+        32.26569590583699
+         97.9646426794348
+        307.2869228453199
+       -13.20108144433967
+         32.1489095602149
+         119.940802630429
+        324.2001123782994
+ 4.43e+10    
+        323.3534550893962
+        121.6273337216303
+        307.0981117251798
+        32.25079311828198
+        98.32998048835704
+         308.219007904867
+       -13.45579031140562
+        32.13399952934618
+        120.5446408044452
+         325.265876277773
+ 4.44e+10    
+        324.4142100901368
+        122.2339510210009
+        308.0319820826326
+        32.23388940545516
+        98.69521313975712
+        309.1525600708082
+       -13.71309579041431
+        32.11708768006472
+        121.1487379178124
+        326.3335970895475
+ 4.45e+10    
+         325.476922294476
+        122.8408108850565
+        308.9672995457296
+        32.21496095719088
+        99.06032764520445
+        310.0875695161491
+        -13.9730267072322
+        32.09815003462212
+        121.7530622270387
+        327.4032677231691
+ 4.46e+10    
+        326.5415850488264
+        123.4478819415705
+        309.9040541584565
+        32.19398409947547
+        99.42531113301405
+        311.0240265555816
+       -14.23561178127374
+        32.07716275150354
+        122.3575821480647
+         328.474881295009
+ 4.47e+10    
+        327.6081918997196
+        124.0551329847627
+        310.8422361172569
+        32.17093530057912
+         99.7901508513948
+        311.9619216482797
+       -14.50087961530307
+        32.05410213161367
+        122.9622662646293
+        329.5484311294787
+ 4.48e+10    
+        328.6767365950217
+        124.6625329835879
+          311.78183577386
+        32.14579117718765
+        100.1548341715857
+        312.9012454006866
+       -14.76885868517493
+        32.02894462446251
+        123.5670833366206
+        330.6239107602419
+ 4.49e+10    
+        329.7472130851449
+        125.2700510900077
+        312.7228436380914
+        32.11852850053207
+        100.5193485909793
+        313.8419885692852
+       -15.03957732951518
+         32.0016668343499
+        124.1720023084073
+        331.7013139314222
+ 4.5e+10     
+        330.8196155242612
+        125.8776566472398
+        313.6652503806692
+        32.08912420251558
+        100.8836817362308
+         314.784142063346
+       -15.31306373934543
+        31.97224552654707
+        124.7769923171517
+         332.780634598806
+ 4.51e+10    
+        331.8939382715015
+         126.485319197989
+        314.6090468359724
+        32.05755538183698
+        101.2478213663552
+        315.7276969476722
+       -15.58934594765123
+        31.94065763347583
+        125.3820227011002
+         333.861866931041
+ 4.52e+10    
+        332.9701758921631
+        127.0930084926575
+        315.5542240048071
+        32.02379931010935
+        101.6117553758087
+         316.672644445318
+       -15.86845181889779
+        31.90688026088234
+        125.9870630078549
+        334.9450053108309
+ 4.53e+10    
+        334.0483231588993
+        127.7006944975295
+        316.5007730571412
+        31.98783343797336
+        101.9754717975583
+        317.6189759402965
+        -16.1504090384949
+        31.87089069400692
+         126.592083002619
+        336.0300443361231
+ 4.54e+10    
+        335.1283750529155
+        128.3083474029324
+        317.4486853348291
+        31.94963540120375
+        102.3389588061347
+        318.5666829802691
+       -16.43524510221249
+        31.83266640374658
+        127.1970526764214
+        337.1169788212986
+ 4.55e+10    
+        336.2103267651535
+        128.9159376313743
+        318.3979523543142
+        31.90918302680828
+        102.7022047206729
+        319.5157572792221
+        -16.7229873055507
+        31.79218505281083
+        127.8019422543119
+        338.2058037983472
+ 4.56e+10    
+        337.2941736974767
+        129.5234358456532
+        319.3485658093179
+        31.86645433911891
+        103.0651980079369
+        320.4661907201262
+       -17.01366273306448
+        31.74942450186946
+        128.4067222035335
+        339.2965145180494
+ 4.57e+10    
+        338.3799114638455
+        130.1308129569391
+         320.300517573504
+        31.82142756587233
+        103.4279272853289
+        321.4179753575754
+       -17.30729824764737
+        31.70436281569057
+         129.011363241664
+        340.3891064511437
+ 4.58e+10    
+        339.4675358914885
+        130.7380401328272
+        321.2537997031334
+        31.77408114428091
+        103.7903813238842
+        322.3711034204167
+       -17.60392047977491
+        31.65697826926929
+        129.6158363447304
+        341.4835752894908
+ 4.59e+10    
+         340.557043022073
+        131.3450888053619
+        322.2084044396933
+         31.7243937270921
+        104.1525490512505
+        323.3255673143571
+       -17.90355581671093
+        31.60724935394446
+        130.2201127552918
+        342.5799169472414
+ 4.6e+10     
+         341.648429112864
+        131.9519306790275
+        323.1643242125124
+        31.67234418863502
+        104.5144195546499
+        324.2813596245588
+       -18.20623039167879
+        31.55515478350399
+        130.8241639904913
+        343.6781275619839
+ 4.61e+10    
+        342.7416906378807
+        132.5585377387085
+        324.1215516413538
+        31.61791163085406
+        104.8759820838279
+        325.2384731182156
+       -18.51197007300048
+        31.50067350027673
+        131.4279618500768
+        344.7782034958989
+ 4.62e+10    
+         343.836824289044
+        133.1648822576176
+        325.0800795389979
+        31.56107538932851
+        105.2372260539825
+        326.1969007471118
+       -18.82080045320452
+        31.44378468121048
+        132.0314784243855
+        345.8801413369014
+ 4.63e+10    
+        344.9338269773267
+        133.7709368051844
+        326.0399009137952
+        31.50181503927573
+        105.5981410486803
+        327.1566356501642
+       -19.13274683810744
+        31.38446774393482
+         132.634686102296
+        346.9839378997811
+ 4.64e+10    
+        346.0326958338836
+        134.3766742549145
+        327.0010089722072
+        31.44011040153921
+        105.9587168227528
+        328.1176711559514
+       -19.44783423586906
+        31.32270235280765
+        133.2375575791428
+        348.0895902273305
+ 4.65e+10    
+        347.1334282111841
+        134.9820677922073
+        327.9633971213327
+        31.37594154855853
+        106.3189433051781
+         329.080000785219
+       -19.76608734602542
+        31.25846842494537
+        133.8400658645944
+        349.1970955914715
+ 4.66e+10    
+        348.2360216841405
+        135.5870909221391
+         328.927058971404
+         31.3092888103219
+        106.6788106019442
+        330.0436182533717
+       -20.08753054850114
+        31.19174613623458
+        134.4421842904932
+        350.3064514943747
+ 4.67e+10    
+        349.3404740512187
+        136.1917174772042
+        329.8919883382763
+        31.24013278029825
+        107.0383089988948
+        331.0085174729486
+       -20.41218789260454
+        31.12251592732464
+        135.0438865186566
+        351.4176556695672
+ 4.68e+10    
+        350.4467833355503
+        136.7959216250192
+        330.8581792458882
+        31.16845432135063
+        107.3974289645588
+        331.9746925560768
+       -20.74008308600701
+        31.05075850960122
+        135.6451465486371
+        352.5307060830442
+ 4.69e+10    
+        351.5549477860334
+        137.3996778759845
+        331.8256259287101
+        31.09423457162712
+        107.7561611529596
+        332.9421378169144
+       -21.07123948371054
+        30.97645487113748
+        136.2459387254409
+        353.6456009343558
+ 4.7e+10     
+        352.6649658784252
+        138.0029610909032
+        332.7943228341715
+        31.01745495043049
+        108.1144964064088
+        333.9108477740667
+        -21.4056800770043
+        30.89958628262444
+         136.846237747204
+        354.7623386577012
+ 4.71e+10    
+         353.776836316428
+        138.6057464885596
+        333.7642646250656
+        30.93809716406427
+        108.4724257582794
+        334.8808171529915
+       -21.74342748241504
+        30.82013430327813
+        137.4460186728263
+        355.8809179230063
+ 4.72e+10    
+        354.8905580327638
+        139.2080096532502
+        334.7354461819406
+        30.85614321165485
+        108.8299404357625
+        335.8520408883827
+       -22.08450393065184
+        30.73808078672273
+        138.0452569295584
+         357.001337636998
+ 4.73e+10    
+        356.0061301902433
+        139.8097265422722
+        335.7078626054669
+        30.77157539094859
+        109.1870318626032
+        336.8245141265388
+       -22.42893125554936
+        30.65340788684892
+        138.6439283205453
+        358.1235969442639
+ 4.74e+10    
+        357.1235521828226
+        140.4108734933642
+        336.6815092187858
+        30.68437630408324
+        109.5436916618193
+        337.7982322277076
+       -22.77673088301148
+        30.56609806364648
+        139.2420090323216
+        359.2476952283071
+ 4.75e+10    
+        358.2428236366516
+        141.0114272321019
+        337.6563815698424
+        30.59452886333153
+        109.8999116583994
+        338.7731907684187
+       -23.12792381995845
+        30.47613408901027
+         139.839475642261
+        360.3736321125917
+ 4.76e+10    
+        359.3639444111143
+        141.6113648792427
+        338.6324754336886
+        30.50201629681759
+        110.2556838819826
+        339.7493855437918
+        -23.4825306432805
+        30.38349905251773
+        140.4363051259749
+        361.5014074615756
+ 4.77e+10    
+        360.4869145998513
+        142.2106639580233
+        339.6097868147801
+        30.40682215420419
+        110.6110005695181
+        340.7268125698309
+       -23.84057148879926
+        30.28817636717853
+        141.0324748646628
+        362.6310213817331
+ 4.78e+10    
+        361.6117345317838
+         142.809302401409
+        340.5883119492444
+        30.30893031235047
+        110.9658541679053
+        341.7054680856976
+       -24.20206604024202
+        30.19014977515413
+        141.6279626524133
+        363.7624742225732
+ 4.79e+10    
+        362.7384047721149
+        143.4072585592863
+        341.5680473071276
+        30.20832498093797
+        111.3202373366128
+        342.6853485559611
+       -24.56703351822929
+        30.08940335344649
+        142.2227467034501
+         364.895766577638
+ 4.8e+10     
+          363.86692612333
+        144.0045112056116
+        342.5489895946285
+        30.10499070806613
+        111.6741429502792
+        343.6664506728368
+       -24.93549266928034
+        29.98592151955543
+        142.8168056593287
+        366.0308992854963
+ 4.81e+10    
+        364.9972996261739
+        144.6010395454999
+        343.5311357563042
+        29.99891238581407
+        112.0275641012914
+        344.6487713584005
+       -25.30746175483835
+         29.8796890371034
+        143.4101185960782
+        367.1678734307229
+ 4.82e+10    
+         366.129526560626
+        145.1968232222638
+        344.5144829772614
+        29.89007525576925
+        112.3804941023435
+        345.6323077667848
+       -25.68295854031816
+        29.77069102142641
+          144.00266503129
+        368.3066903448684
+ 4.83e+10    
+        367.2636084468584
+        145.7918423243982
+        345.4990286853266
+         29.7784649145215
+        112.7329264889745
+        346.6170572863522
+       -26.06200028417972
+        29.65891294513154
+        144.5944249311495
+        369.4473516074156
+ 4.84e+10    
+        368.3995470461838
+        146.3860773925067
+        346.4847705531892
+        29.66406731912144
+        113.0848550220853
+        347.6030175418557
+       -26.44460372703063
+        29.54434064361674
+        145.1853787174127
+        370.5898590467188
+ 4.85e+10    
+        369.5373443619857
+        146.9795094261748
+        347.4717065005317
+        29.54686879250221
+        113.4362736904329
+        348.5901863965714
+       -26.83078508075872
+        29.42696032055736
+        145.7755072743269
+        371.7342147409422
+ 4.86e+10    
+        370.6770026406419
+        147.5721198907849
+        348.4598346961383
+        29.42685602886454
+        113.7871767131065
+        349.5785619544171
+       -27.22056001770029
+         29.3067585533525
+        146.3647919554904
+        372.8804210189676
+ 4.87e+10    
+        371.8185243724255
+        148.1638907242717
+        349.4491535599752
+        29.30401609902267
+        114.1375585419785
+         350.568142562048
+       -27.61394365984391
+        29.18372229853519
+        146.9532145906571
+        374.0284804613065
+ 4.88e+10    
+        372.9619122924045
+        148.7548043438218
+        350.4396617652594
+        29.17833645571183
+         114.487413864136
+        351.5589268109314
+       -28.01095056807524
+        29.05783889714238
+        147.5407574924798
+        375.1783959009857
+ 4.89e+10    
+        374.1071693813126
+        149.3448436525115
+        351.4313582404985
+        29.04980493885459
+        114.8367376042892
+        352.5509135394019
+       -28.41159473146447
+        28.92909608004455
+        148.1274034631925
+        376.3301704244242
+ 4.9e+10     
+        375.2542988664148
+        149.9339920458858
+        352.4242421715162
+        28.91840978078739
+        115.1855249271583
+           353.5441018347
+       -28.81588955659878
+        28.79748197323579
+        148.7131358012334
+        377.4838073722925
+ 4.91e+10    
+        376.4033042223549
+        150.5222334184739
+        353.4183130034509
+         28.7841396114442
+         115.533771239838
+        354.5384910349773
+       -29.22384785696427
+        28.66298510308027
+        149.2979383078042
+        378.6393103403609
+ 4.92e+10    
+        377.5541891719885
+        151.1095521702463
+        354.4135704427336
+        28.64698346349765
+        115.8814721941387
+        355.5340807312993
+         -29.635481842379
+        28.52559440151661
+        149.8817952933666
+        379.7966831803259
+ 4.93e+10    
+         378.706957687198
+        151.6959332130058
+        355.4100144590476
+        28.50693077745641
+        116.2286236889069
+        356.5308707696096
+       -30.05080310848051
+        28.38529921121897
+        150.4646915840783
+          380.95593000063
+ 4.94e+10    
+        379.8616139896932
+        152.2813619767179
+        356.4076452872673
+        28.36397140671802
+        116.5752218723212
+        357.5288612526871
+       -30.46982262627078
+        28.24208929071274
+        151.0466125281612
+        382.1170551672581
+ 4.95e+10    
+        381.0181625517955
+        152.8658244157742
+        357.4064634293638
+        28.21809562257599
+        116.9212631441655
+        358.5280525420696
+       -30.89255073172104
+        28.09595481944491
+        151.6275440022051
+        383.2800633045157
+ 4.96e+10    
+        382.1766080972048
+         153.449307015195
+        358.4064696563058
+        28.06929411918084
+        117.2667441580797
+        359.5284452599666
+       -31.31899711544062
+        27.94688640280829
+        152.2074724174086
+        384.4449592958012
+ 4.97e+10    
+        383.3369556017475
+        154.0317967967614
+        359.4076650099263
+        27.91755801845326
+        117.6116618237866
+        360.5300402911425
+       -31.74917081241112
+        27.79487507711826
+        152.7863847257493
+        385.6117482843495
+ 4.98e+10    
+        384.4992102941118
+        154.6132813250865
+        360.4100508047696
+        27.76287887495016
+        117.9560133092958
+        361.5328387847857
+       -32.18308019178993
+         27.6399123145414
+        153.3642684260923
+        386.7804356739662
+ 4.99e+10    
+          385.66337765656
+        155.1937487136152
+        361.4136286299212
+        27.60524868068086
+         118.299796043084
+        362.5368421563488
+       -32.62073294678563
+        27.48199002797502
+        153.9411115702243
+         387.951027129736
+ 5e+10       
+         386.829463425625
+         155.773187630559
+        362.4184003508097
+        27.44465986987363
+        118.6430077162504
+        363.5420520893701
+       -33.06213608460848
+        27.32110057587663
+        154.5169027688253
+        389.1235285787229
+ 5.01e+10    
+        387.9974735927873
+        156.3515873047633
+         363.424368110987
+        27.28110532369184
+        118.9856462846502
+        364.5484705372739
+       -33.50729591649828
+        27.15723676704332
+        155.0916311973679
+        390.2979462106445
+ 5.02e+10    
+        389.1674144051362
+        156.9289375315034
+        364.4315343338913
+         27.1145783748986
+        119.3277099710023
+        365.5560997251497
+       -33.95621804783326
+        26.99039186533877
+        155.6652866019483
+        391.4742864785308
+ 5.03e+10    
+        390.3392923660074
+        157.5052286782128
+        365.4399017245777
+        26.94507281246877
+        119.6691972669739
+        366.5649421515042
+        -34.4089073683227
+        26.82055959436799
+        156.2378593050452
+        392.6525560993601
+ 5.04e+10    
+        391.5131142356042
+        158.0804516901427
+        366.4494732714402
+        26.77258288614784
+        120.0101069352405
+        367.5750005899967
+       -34.86536804228523
+        26.64773414209976
+        156.8093402112112
+         393.832762054683
+ 5.05e+10    
+        392.6888870315989
+        158.6545980959478
+        367.4602522478953
+        26.59710331095732
+        120.3504380115202
+        368.5862780911472
+       -35.32560349901768
+        26.47191016543307
+        157.3797208126887
+        395.0149115912191
+ 5.06e+10    
+        393.8666180297137
+        159.2276600132055
+        368.4722422140579
+        26.41862927164491
+        120.6901898065875
+        369.5987779840294
+       -35.78961642325547
+        26.29308279471088
+        157.9489931949569
+        396.1990122214374
+ 5.07e+10    
+        395.0463147642786
+        159.7996301538584
+        369.4854470183816
+        26.23715642707885
+        121.0293619082557
+        370.6125038779288
+       -36.25740874572811
+        26.11124763817639
+        158.5171500422042
+        397.3850717241177
+ 5.08e+10    
+        396.2279850287745
+        160.3705018295885
+        370.4998707992835
+        26.05268091458709
+        121.3679541833415
+        371.6274596639931
+       -36.72898163381323
+        25.92640078637368
+        159.0841846427292
+        398.5730981448867
+ 5.09e+10    
+        397.4116368763511
+        160.9402689571192
+        371.5155179867471
+        25.86519935423787
+        121.7059667795999
+        372.6436495168477
+       -37.20433548229083
+        25.73853881649119
+        159.6500908942657
+        399.7630997967362
+ 5.1e+10     
+        398.5972786203234
+        161.5089260634387
+        372.5323933038924
+         25.6747088530633
+        122.0434001276355
+        373.6610778961921
+       -37.68346990420197
+        25.54765879664635
+        160.2148633092372
+         400.955085260525
+ 5.11e+10    
+        399.7849188346484
+        162.0764682909573
+        373.5505017685363
+        25.48120700922406
+        122.3802549427897
+        374.6797495483792
+       -38.16638372181339
+        25.35375829011213
+        160.7784970199319
+        402.1490633854474
+ 5.12e+10    
+        400.9745663543824
+        162.6428914025861
+         374.569848694722
+        25.28469191611502
+        122.7165322270007
+          375.69966950796
+       -38.65307495769171
+        25.15683535948383
+        161.3409877836075
+        403.3450432894913
+ 5.13e+10    
+        402.1662302761107
+        163.2081917867404
+        375.5904396942217
+        25.08516216640955
+        123.0522332706395
+        376.7208430992162
+       -39.14354082588991
+        24.95688857078501
+        161.9023319875163
+        404.5430343598692
+ 5.14e+10    
+        403.3599199583587
+        163.7723664622725
+        376.6122806780263
+        24.88261685604483
+        123.3873596543193
+        377.7432759376639
+        -39.6377777232486
+        24.75391699751287
+        162.4625266538574
+        405.7430462534267
+ 5.15e+10    
+        404.5556450219821
+        164.3354130833244
+        377.6353778578024
+        24.67705558814354
+        123.7219132506812
+        378.7669739315344
+       -40.13578122081516
+        24.54792022462174
+        163.0215694446513
+        406.9450888970318
+ 5.16e+10    
+        405.7534153505276
+        164.8973299441077
+        378.6597377473317
+        24.46847847687512
+        124.0558962261516
+        379.7919432832334
+       -40.63754605538303
+        24.33889835244378
+        163.5794586665367
+        408.1491724879376
+ 5.17e+10    
+        406.9532410905815
+        165.4581159836077
+        379.6853671639265
+        24.25688615125232
+        124.3893110426764
+        380.8181904907753
+        -41.1430661211544
+        24.12685200054647
+        164.1361932754917
+         409.355307494123
+ 5.18e+10    
+        408.1551326520843
+        166.0177707902067
+        380.7122732298104
+        24.04227975886488
+        124.7221604594257
+        381.8457223491923
+       -41.65233446152926
+        23.91178231152596
+        164.6917728814756
+        410.5635046546118
+ 5.19e+10    
+        409.3591007086272
+        166.5762946062372
+        381.7404633734996
+        23.82466096954933
+        125.0544475344783
+        382.8745459519276
+        -42.1653432610221
+        23.69369095473646
+        165.2461977529953
+        411.7737749797684
+ 5.2e+10     
+        410.5651561977279
+        167.1336883324513
+        382.7699453311328
+        23.60403197899265
+        125.3861756264738
+        383.9046686921934
+       -42.68208383731029
+         23.4725801299534
+        165.7994688215908
+         412.986129751568
+ 5.21e+10    
+        411.7733103210709
+        167.6899535324165
+        383.8007271477974
+        23.38039551227042
+        125.7173483962425
+        384.9360982643162
+       -43.20254663341717
+        23.24845257097077
+        166.3515876862426
+        414.2005805238408
+ 5.22e+10    
+        412.9835745447429
+        168.2450924368332
+        384.8328171788244
+        23.15375482731961
+        126.0479698084081
+        385.9688426650496
+       -43.72672121002994
+         23.0213115491324
+        166.9025566177025
+        415.4171391225017
+ 5.23e+10    
+        414.1959605994228
+         168.799107947772
+        385.8662240910567
+         22.9241137183427
+         126.378044132964
+        387.0029101948696
+       -44.25459623795859
+          22.791160876795
+        167.4523785627413
+         416.635817645741
+ 5.24e+10    
+        415.4104804805646
+        169.3520036428357
+        386.9009568641037
+        22.69147651914606
+        126.7075759468231
+        388.0383094592446
+       -44.78615949073487
+        22.55800491072399
+        168.0010571483192
+        417.8566284642063
+ 5.25e+10    
+        416.6271464485428
+        169.9037837792389
+         387.937024791556
+        22.45584810640803
+        127.0365701353415
+         389.075049369877
+       -45.32139783735673
+        22.32184855542005
+        168.5485966856774
+         419.079584221144
+ 5.26e+10    
+        417.8459710287844
+        170.4544532978123
+        388.9744374821958
+        22.21723390287971
+        127.3650318938151
+        390.1131391459281
+       -45.86029723517872
+        22.08269726637722
+        169.0950021743468
+        420.3046978325324
+ 5.27e+10    
+        419.0669670118645
+        171.0040178269254
+        390.0132048611672
+        21.97563988051582
+        127.6929667289505
+        391.1525883152139
+       -46.40284272295215
+        21.84055705327027
+         169.640279306079
+        421.5319824871731
+ 5.28e+10    
+        420.2901474535876
+        171.5524836863306
+         391.053337171129
+        21.73107256353514
+        128.0203804603083
+        392.1934067153783
+       -46.94901841401639
+        21.59543448307265
+        170.1844344686946
+        422.7614516467721
+ 5.29e+10    
+        421.5155256750353
+        172.0998578909275
+        392.0948449733864
+        21.48353903141101
+        128.3472792217209
+        393.2356044950421
+       -47.49880748964453
+         21.3473366831027
+        170.7274747498528
+         423.993119045984
+ 5.3e+10     
+        422.7431152625914
+        172.6461481544479
+         393.137739148992
+        21.23304692179006
+        128.6736694626823
+        394.2791921149322
+       -48.05219219254624
+        21.09627134399845
+        171.2694079407387
+        425.2269986924381
+ 5.31e+10    
+        423.9729300679458
+        173.1913628930598
+        394.1820308998296
+        20.97960443333942
+        128.9995579497117
+         395.324180348975
+       -48.60915382052794
+         20.8422467226207
+        171.8102425396696
+        426.4631048667354
+ 5.32e+10    
+        425.2049842080635
+        173.7355112288926
+         395.227731749669
+        20.72322032852207
+        129.3249517676912
+        396.3705802853831
+       -49.16967272031582
+        20.58527164488309
+        172.3499877556213
+        427.7014521224193
+ 5.33e+10    
+        426.4392920651377
+        174.2786029934806
+        396.2748535451985
+         20.4639039362992
+        129.6498583211744
+        397.4184033277002
+       -49.73372828154086
+        20.32535550850884
+        172.8886535116706
+        428.9420552859234
+ 5.34e+10    
+        427.6758682865105
+        174.8206487311287
+        397.3234084570381
+        20.20166515475886
+        129.9742853356701
+        398.4676611958337
+       -50.30129893089102
+        20.06250828571444
+        173.4262504483594
+        430.1849294564904
+ 5.35e+10    
+        428.9147277845662
+        175.3616597021923
+        398.3734089807161
+        19.93651445367171
+        130.2982408588989
+        399.5183659270607
+       -50.87236212642993
+        19.79674052581838
+        173.9627899269739
+        431.4300900060653
+ 5.36e+10    
+        430.1558857366088
+         175.901647886284
+        399.4248679376363
+         19.6684628769717
+        130.6217332620208
+         400.570529877005
+       -51.44689435208703
+        19.52806335777584
+        174.4982840327453
+        432.6775525791646
+ 5.37e+10    
+        431.3993575846964
+        176.4406259853914
+        400.4777984760133
+          19.397522045163
+         130.944771240839
+         401.624165720597
+       -52.02487111231871
+        19.25648849263765
+         175.032745577965
+        433.9273330927149
+ 5.38e+10    
+        432.6451590354682
+        176.9786074269226
+        401.5322140717856
+        19.12370415765092
+        131.2673638169741
+        402.6792864530045
+       -52.60626692694517
+        18.98202822593429
+        175.5661881050218
+         435.179447735869
+ 5.39e+10    
+        433.8933060599321
+        177.5156063666635
+        402.5881285295027
+        18.84702199499747
+        131.5895203390121
+        403.7359053905409
+        -53.1910553261623
+        18.70469543998315
+        176.0986258893541
+        436.4339129697931
+ 5.4e+10     
+        435.1438148932263
+         178.051637691658
+        403.6455559831903
+        18.56748892110147
+        131.9112504836256
+        404.7940361715482
+       -53.77920884573326
+        18.42450360611948
+        176.6300739423218
+          437.69074552743
+ 5.41e+10    
+        436.3967020343604
+        178.5867170230078
+        404.7045108971938
+        18.28511888530153
+        132.2325642566678
+        405.8536927572586
+       -54.37069902235941
+        18.14146678685102
+        177.1605480139956
+        438.9499624132284
+ 5.42e+10    
+        437.6519842459296
+        179.1208607185889
+        405.7650080669932
+        17.99992642440288
+        132.5534719942391
+        406.9148894326316
+       -54.96549638923449
+        17.85559963793413
+        177.6900645958637
+        440.2115809028574
+ 5.43e+10    
+         438.909678553794
+         179.654085875689
+        406.8270626199954
+        17.71192666462608
+        132.8739843637269
+        407.9776408071588
+       -55.56357047178249
+        17.56691741037367
+        178.2186409234588
+        441.4756185428834
+ 5.44e+10    
+        440.1698022467406
+        180.1864103335629
+        407.8906900163061
+        17.42113532347933
+        133.1941123648189
+        409.0419618156625
+       -56.16488978358184
+        17.27543595234301
+        178.7462949788994
+        442.7420931504232
+ 5.45e+10    
+        441.4323728761142
+        180.7178526759078
+        408.9559060494725
+        17.12756871155186
+        133.5138673304869
+        410.1078677190478
+       -56.76942182247713
+        16.98117171102754
+        179.2730454933526
+        444.0110228127746
+ 5.46e+10    
+        442.6974082554198
+        181.2484322332584
+        410.0227268472079
+        16.83124373423009
+        133.8332609279477
+        411.1753741050493
+       -57.37713306688123
+        16.68414173438748
+        179.7989119494131
+        445.2824258870155
+ 5.47e+10    
+        443.9649264599042
+        181.7781690852988
+        411.0911688720858
+         16.5321778933341
+        134.1523051595923
+        412.2444968889461
+       -57.98798897226791
+        16.38436367284309
+        180.3239145834008
+        446.5563209995731
+ 5.48e+10    
+        445.2349458261058
+        182.3070840630971
+        412.1612489222155
+        16.23038928867581
+        134.4710123638913
+        413.3152523142478
+       -58.60195396785808
+         16.0818557808793
+         180.848074387577
+        447.8327270457764
+ 5.49e+10    
+        446.5074849513744
+        182.8351987512562
+        413.2329841318963
+        15.92589661953821
+        134.7893952162719
+         414.387656953367
+       -59.21899145350019
+         15.7766369185715
+        181.3714131122778
+        449.1116631893709
+ 5.5e+10     
+        447.7825626933741
+        183.3625354899851
+        414.3063919722349
+        15.61871918607482
+        135.1074667299683
+        415.4617277082633
+       -59.83906379674715
+        15.46872655303009
+        181.8939532679678
+        450.3931488620113
+ 5.51e+10    
+        449.0601981695528
+         183.889117377093
+        415.3814902517597
+        15.30887689062941
+        135.4252402568445
+          416.53748181106
+       -60.46213233013079
+        15.15814475976615
+        182.4157181272105
+        451.6772037627287
+ 5.52e+10    
+        450.3404107565851
+        184.4149682698986
+        416.4582971169944
+        14.99639023897571
+        135.7427294881906
+        417.6149368246407
+       -61.08815734863552
+        14.84491222397519
+        182.9367317265584
+        452.9638478573669
+ 5.53e+10    
+        451.6232200897883
+        184.9401127870591
+        417.5368310530106
+        14.68128034147715
+        136.0599484554923
+        418.6941106432218
+       -61.71709810737247
+        14.52905024174114
+        183.4570188683619
+        454.2531013779956
+ 5.54e+10    
+        452.9086460625147
+        185.4645763103252
+        418.6171108839662
+         14.3635689141662
+        136.3769115311726
+         419.775021492903
+       -62.34891281945536
+        14.21058072115812
+        183.9766051224959
+         455.544984822291
+ 5.55e+10    
+         454.196708825515
+        185.9883849862096
+        419.6991557736145
+         14.0432782797426
+        136.6936334293073
+        420.8576879321864
+       -62.98355865408011
+        13.88952618337225
+        184.4955168280082
+        456.8395189528978
+ 5.56e+10    
+        455.4874287862747
+        186.5115657275801
+        420.7829852257855
+        13.72043136849152
+         137.010129206314
+        421.9421288524838
+       -63.62099173480838
+        13.56590976354076
+        185.0137810946851
+        458.1367247967565
+ 5.57e+10    
+        456.7808266083253
+          187.03414621517
+        421.8686190848529
+        13.39505171911987
+        137.3264142616131
+        423.0283634785915
+       -64.26116713805703
+        13.23975521171045
+        185.5314258045359
+        459.4366236444101
+ 5.58e+10    
+        458.0769232105257
+        187.5561548990136
+        422.9560775361706
+        13.06716347951246
+        137.6425043382624
+        424.1164113691418
+       -64.90403889179399
+        12.91108689361351
+        186.0484796132001
+        460.7392370492762
+ 5.59e+10    
+        459.3757397663215
+        188.0776209997971
+         424.045381106487
+        12.73679140740576
+        137.9584155235658
+         425.206292417038
+       -65.54955997444284
+        12.57992979138171
+        186.5649719512722
+         462.044586826904
+ 5.6e+10     
+        460.6772977029802
+         188.598574510138
+        425.1365506643475
+        12.40396087098134
+        138.2741642496551
+        426.2980268498592
+       -66.19768231399523
+        12.24630950417895
+        187.0809330255471
+        463.3526950541928
+ 5.61e+10    
+        461.9816187007863
+         189.119046195777
+        426.2296074204519
+        12.06869784937721
+         138.589767294043
+        427.3916352302457
+       -66.84835678733397
+         11.9102522487503
+        187.5963938201862
+        464.6635840685935
+ 5.62e+10    
+        463.2887246922292
+        189.6390675967004
+        427.3245729280108
+        11.73102893311707
+        138.9052417801535
+        428.4871384562579
+       -67.50153321976634
+         11.5717848598904
+        188.1113860978056
+         465.977276467275
+ 5.63e+10    
+        464.5986378611521
+         190.158671028179
+        428.4214690830671
+        11.39098132445923
+        139.2206051778214
+         429.584557761715
+       -68.15716038476974
+        11.23093479082786
+        188.6259424004818
+        467.2937951062736
+ 5.64e+10    
+         465.911380641876
+        190.6778895817296
+        429.5203181247939
+        11.04858283766237
+         139.535875303769
+          430.68391471651
+       -68.81518600394884
+         10.8877301135283
+        189.1400960506826
+        468.6131630996072
+ 5.65e+10    
+        467.2269757183055
+        191.1967571260031
+        430.6211426357842
+        10.70386189917011
+        139.8510703220544
+        431.7852312269011
+       -69.47555674720689
+        10.54219951891396
+        189.6538811521179
+        469.9354038183718
+ 5.66e+10    
+         468.545446022999
+        191.7153083075902
+        431.7239655422929
+        10.35684754771419
+        140.1662087444934
+        432.8885295357791
+       -70.13821823312995
+        10.19437231700164
+        190.1673325905114
+        471.2605408898033
+ 5.67e+10    
+        469.8668147362212
+        192.2335785517543
+        432.8288101144823
+        10.00756943433457
+        140.4813094310563
+        433.9938322229157
+       -70.80311502958646
+        9.844278436957154
+         190.680486034296
+        472.5885981963226
+ 5.68e+10    
+        471.1911052849649
+        192.7516040630858
+        433.9356999666296
+        9.656057822319365
+        140.7963915902384
+        435.1011622051864
+       -71.47019065454094
+        9.491948427068074
+        191.1933779352328
+        473.9195998745482
+ 5.69e+10    
+        472.5183413419501
+        193.2694218260805
+        435.0446590573137
+        9.302343587060854
+        141.1114747794019
+        436.2105427367687
+       -72.13938757708461
+        9.137413454632267
+        191.7060455289486
+        475.2535703142831
+ 5.7e+10     
+        473.8485468245962
+        193.7870696056435
+        436.1557116895881
+        8.946458215832036
+        141.4265789050961
+        437.3219974093246
+       -72.81064721867993
+        8.780705305766467
+        192.2185268354024
+        476.5905341574834
+ 5.71e+10    
+        475.1817458939729
+         194.304585947516
+        437.2688825111204
+        8.588433807479266
+        141.7417242233476
+        438.4355501521522
+       -73.48390995462374
+        8.421856385129473
+        192.7308606592718
+        477.9305162971953
+ 5.72e+10    
+        476.5179629537186
+        194.8220101786278
+         438.384196514317
+        8.228303072034723
+        142.0569313399272
+        439.5512252323224
+       -74.15911511572534
+        8.060899715564613
+        193.2430865902638
+        479.2735418764625
+ 5.73e+10    
+        477.8572226489449
+        195.3393824073766
+        439.5016790364284
+        7.866099330246806
+        142.3722212105901
+          440.66904725479
+       -74.83620099020274
+        7.697868937659319
+        193.7552450033519
+        480.6196362872253
+ 5.74e+10    
+        479.1995498651023
+        195.8567435238275
+        440.6213557596213
+        7.501856513028516
+        142.6876151412909
+        441.7890411624809
+       -75.51510482579488
+        7.332798309222625
+        194.2673770589362
+        481.9688251691761
+ 5.75e+10    
+        480.5449697268393
+        196.3741351998487
+        441.7432527110461
+        7.135609160825044
+        143.0031347883708
+        442.9112322363623
+       -76.19576283209226
+         6.96572270467998
+        194.7795247029294
+        483.3211344086019
+ 5.76e+10    
+        481.8935075968199
+        196.8915998891617
+         442.867396262861
+        6.767392422900347
+        143.3188021587243
+        444.0356460954882
+       -76.87811018308426
+        6.596677614385655
+        195.2917306667676
+        484.6765901371959
+ 5.77e+10    
+        483.2451890745276
+        197.4091808273278
+        443.9938131322589
+        6.397242056541184
+         143.634639609934
+        445.1623086970185
+       -77.56208101992353
+        6.225699143854932
+          195.80403846735
+        486.0352187308526
+ 5.78e+10    
+         484.600039995044
+        197.9269220316577
+        445.1225303814525
+        6.025194426182322
+        143.9506698503862
+        446.2912463362285
+       -78.24760845390885
+        5.852824012912166
+        196.3164924069011
+        487.3970468084311
+ 5.79e+10    
+        485.9580864278021
+        198.4448683010503
+        446.2535754176521
+        5.651286502449278
+        144.2669159393576
+         447.422485646487
+       -78.93462456968345
+        5.478089554759073
+         196.829137572763
+        488.7621012304959
+ 5.8e+10     
+        487.3193546753124
+        198.9630652157582
+        447.3869759930145
+        5.275555861120624
+        144.5834012870775
+        448.5560535992134
+       -79.62306042865227
+        5.101533714960375
+        197.3420198371147
+        490.1304090980399
+ 5.81e+10    
+        488.6838712718761
+        199.4815591370836
+         448.522760204575
+        4.898040682011093
+        144.9001496547669
+        449.6919775038179
+       -80.31284607261392
+        4.723195050348782
+        197.8551858566164
+         491.501997751177
+ 5.82e+10    
+        490.0516629822668
+        200.0003972070029
+        449.6609564941539
+        4.518779747773079
+        145.2171851546497
+        450.8302850076207
+       -81.00391052761123
+        4.343112727848965
+        198.3686830719878
+        492.8768947678153
+ 5.83e+10    
+        491.4227568003884
+        200.5196273477217
+        450.8015936482535
+         4.13781244261923
+        145.5345322499431
+        451.9710040957461
+       -81.69618180799574
+        3.961326523220613
+        198.8825597075098
+        494.2551279623058
+ 5.84e+10    
+        492.7971799479216
+        201.0392982611569
+        451.9447007979157
+        3.755178750964904
+        145.8522157548188
+        453.1141630909971
+       -82.38958692070983
+         3.57787681972038
+        199.3968647704577
+        495.6367253840696
+ 5.85e+10    
+        494.1749598729336
+        201.5594594283555
+        453.0903074185815
+        3.370919255991566
+        146.1702608343451
+        454.2597906537154
+        -83.0840518697828
+         3.19280460668481
+        199.9116480504671
+        497.0217153162014
+ 5.86e+10    
+        495.5561242484733
+        202.0801611088359
+         454.238443329909
+        2.985075138129874
+        146.4886930043984
+        455.4079157816063
+       -83.77950166104141
+        2.806151478032259
+        200.4269601188242
+        498.4101262740513
+ 5.87e+10    
+         496.940700971148
+        202.6014543398711
+          455.38913869559
+        2.597688173466718
+        146.8075381315574
+        456.5585678095644
+        -84.4758603070354
+        2.417959630685285
+        200.9428523276936
+        499.8019870037853
+ 5.88e+10    
+        498.3287181596699
+        203.1233909356948
+        456.5424240231327
+        2.208800732070236
+        147.1268224329666
+        457.7117764094578
+       -85.17305083217552
+        2.028271862913996
+        201.4593768092725
+        501.1973264809212
+ 5.89e+10    
+        499.7202041533887
+         203.646023486647
+        457.6983301636336
+         1.81845577623964
+        147.4465724761813
+        458.8675715899079
+       -85.87099527808464
+        1.637131572599975
+        201.9765864748797
+        502.5961739088469
+ 5.9e+10     
+        501.1151875107975
+        204.1694053582492
+        458.8568883115218
+        1.426696858675559
+         147.766815178985
+        460.0259836960397
+       -86.56961470915999
+        1.244582755421581
+        202.4945350139774
+        503.9985587173151
+ 5.91e+10    
+        502.5136970080251
+        204.6935906902143
+        460.0181300042917
+        1.033568120573241
+         148.087577809185
+        461.1870434092151
+       -87.26882921834653
+       0.8506700029612819
+        203.0132768931228
+        505.4045105609172
+ 5.92e+10    
+        503.9157616372977
+        205.2186343953918
+        461.1820871222125
+       0.6391142896397266
+        148.4088879843846
+        462.3507817467524
+        -87.9685579331211
+       0.4554385007344024
+        203.5328673548589
+        506.8140593175368
+ 5.93e+10    
+        505.3214106053888
+        205.7445921586466
+         462.348791888018
+       0.2433806780324339
+        148.7307736717311
+        463.5172300616154
+       -88.66871902168418
+      0.05893402614045939
+        204.0533624165349
+        508.2272350867808
+ 5.94e+10    
+        506.7306733320482
+        206.2715204356753
+        463.5182768665783
+      -0.1535868197766028
+        149.0532631876402
+        464.6864200420906
+        -89.3692296993605
+      -0.3387970536622493
+        204.5748188690624
+        509.6440681883964
+ 5.95e+10    
+        508.1435794484044
+        206.7994764517553
+        464.6905749645529
+      -0.5517417292133242
+        149.3763851974992
+        465.8583837114468
+       -90.07000623520558
+      -0.7377077839593404
+        205.0972942756104
+        511.0645891606588
+ 5.96e+10    
+        509.5601587953545
+        207.3285182004342
+        465.8657194300219
+      -0.9510369978896467
+        149.7001687153449
+        467.0331534275674
+       -90.77096395881955
+        -1.13775062475934
+        205.6208469702315
+        512.4888287587484
+ 5.97e+10    
+        510.9804414219373
+        207.8587044421548
+        467.0437438521077
+       -1.351424997966118
+        150.0246431035213
+        468.2107618825717
+       -91.47201726736334
+       -1.538877453148126
+        206.1455360564285
+        513.9168179531026
+ 5.98e+10    
+        512.4044575836764
+        208.3900947028184
+         468.224682160568
+       -1.752857528588835
+        150.3498380723119
+         469.391242102416
+       -92.17307963277906
+       -1.941039565719135
+        206.6714214056564
+        515.3485879277515
+ 5.99e+10    
+        513.8322377409113
+        208.9227492722846
+        469.4085686253712
+       -2.155285818401001
+        150.6757836795517
+        470.5746274464718
+       -92.87406360921202
+       -2.344187681078678
+        207.1985636557629
+        516.7841700786332
+ 6e+10       
+        515.2638125571175
+        209.4567292028143
+        470.5954378562674
+       -2.558660528127177
+        151.0025103302162
+        471.7609516070906
+       -93.57488084063283
+       -2.748271942425074
+        207.7270242093678
+        518.2235960118918
+ 6.01e+10    
+        516.6992128971982
+        209.9920963074481
+        471.7853248023186
+       -2.962931753231661
+        151.3300487759876
+        472.9502486091495
+       -94.27544206865863
+       -3.153241920202541
+          208.25686523218
+         519.666897542156
+ 6.02e+10    
+         518.138469825755
+        210.5289131583288
+        472.9782647514342
+       -3.368049026647629
+        151.6584301148003
+        474.1425528095756
+       -94.97565714057102
+       -3.559046614827565
+        208.7881496512581
+        521.1141066908053
+ 6.03e+10    
+        519.5816146053576
+        211.0672430849616
+        474.1742933298744
+       -3.773961321580007
+        151.9876857903636
+        475.3378988968573
+       -95.67543501753084
+       -3.965634459489447
+        209.3209411532048
+        522.5652556842028
+ 6.04e+10    
+        521.0286786947808
+        211.6071501724175
+        475.3734465017379
+        -4.18061705437839
+        152.3178475916629
+        476.5363218905359
+       -96.37468378298507
+       -4.372953323021068
+        209.8553041823101
+        524.0203769519376
+ 6.05e+10    
+         522.479693747233
+        212.1486992594799
+        476.5757605684392
+       -4.587964087481236
+        152.6489476524399
+        477.7378571406762
+       -97.07331065126826
+       -4.780950512844424
+        210.3913039386306
+        525.4795031250221
+ 6.06e+10    
+        523.9346916085649
+        212.6919559367325
+        477.7812721681656
+       -4.995949732430448
+        152.9810184506516
+        478.9425403273278
+       -97.77122197639304
+       -5.189572777983782
+        210.9290063760144
+        526.9426670340918
+ 6.07e+10    
+         525.393704315463
+        213.2369865445906
+        478.9900182753076
+       -5.404520752955356
+         153.314092807907
+        480.1504074599605
+       -98.46832326103018
+       -5.598766312153341
+        211.4684782000661
+        528.4099017075785
+ 6.08e+10    
+         526.856764093626
+        213.7838581712782
+        480.2020361998943
+       -5.813623368125599
+        153.6482038888846
+        481.3614948768907
+       -99.16451916567435
+       -6.008476756910813
+        212.0097868660588
+        529.8812403698752
+ 6.09e+10    
+         528.323903355934
+        214.3326386507495
+        481.4173635869884
+       -6.223203255572868
+        153.9833852007267
+        482.5758392446828
+       -99.85971351799701
+       -6.418649204884284
+        212.5530005767882
+        531.3567164394783
+ 6.1e+10     
+        529.7951547005856
+        214.8833965605538
+        482.6360384160809
+       -6.633205554779803
+        154.3196705924167
+        483.7934775575423
+       -100.5538093223794
+       -6.829228203064375
+        213.0981882803736
+        532.8363635271216
+ 6.11e+10    
+        531.2705509092342
+        215.4362012196484
+        483.8580990004619
+       -7.043574870436281
+        154.6570942541327
+        485.0144471366871
+       -101.2467087696294
+       -7.240157756167417
+        213.6454196680014
+        534.3202154338862
+ 6.12e+10    
+        532.7501249451084
+        215.9911226861602
+        485.0835839865828
+       -7.454255275862844
+        154.9956907165819
+        486.2387856297026
+       -101.9383132468742
+       -7.651381330063398
+        214.1947651716204
+        535.8083061493064
+ 6.13e+10    
+        534.2339099511171
+        216.5482317550916
+        486.3125323533932
+        -7.86519031649849
+        155.3354948503163
+        487.4665310098883
+       -102.6285233476329
+       -8.062841855273406
+        214.7462959615784
+         537.300669849452
+ 6.14e+10    
+        535.7219392479277
+        217.1075999559746
+        487.5449834116679
+       -8.276323013455061
+        155.6765418650255
+        488.6977215755695
+       -103.3172388820599
+        -8.47448173053079
+        215.3000839442101
+        538.7973408950013
+ 6.15e+10    
+        537.2142463320567
+        217.6692995504778
+         488.780976803321
+       -8.687595867134737
+        156.0188673088149
+        489.9323959494264
+       -104.0043588873646
+       -8.886242826409291
+        215.8562017593745
+        540.2983538293037
+ 6.16e+10    
+        538.7108648739264
+        218.2334035299581
+        490.0205525006959
+       -9.098950860912453
+        156.3625070674583
+        491.1705930777687
+       -104.6897816383971
+       -9.298066489015081
+         216.414722777937
+        541.8037433764175
+ 6.17e+10    
+        540.2118287159105
+        218.7999856129646
+        491.2637508058515
+       -9.510329464880492
+        156.7074973636362
+        492.4123522298248
+       -105.3734046584043
+        -9.70989354374308
+        216.9757210992065
+        543.3135444391492
+ 6.18e+10    
+        541.7171718703817
+        219.3691202426963
+        492.5106123498235
+       -9.921672639655807
+        157.0538747561521
+        493.6577129970032
+       -106.0551247299502
+       -10.12166429909644
+        217.5392715483197
+        544.8277920970689
+ 6.19e+10    
+        543.2269285177292
+        219.9408825844057
+        493.7611780918757
+       -10.33292084024855
+         157.401676139131
+        494.9067152921367
+       -106.7348379059978
+       -10.53331855056871
+        218.1054496735792
+          546.34652160452
+ 6.2e+10     
+        544.7411330043738
+        220.5153485227609
+        495.0154893187415
+       -10.74401401999116
+        157.7509387412007
+        496.1593993487249
+       -107.4124395211538
+       -10.94479558458754
+        218.6743317437403
+        547.8697683886119
+ 6.21e+10    
+        546.2598198407742
+        221.0925946591545
+        496.2735876438367
+       -11.15489163452897
+        158.1017001246497
+        497.4158057201446
+        -108.087824203069
+       -11.35603418251972
+        219.2459947452551
+        549.3975680472081
+ 6.22e+10    
+        547.7830236994135
+        221.6726983089733
+        497.5355150064791
+       -11.56549264586787
+        158.4539981845746
+        498.6759752788601
+       -108.7608858839939
+       -11.76697262473584
+         219.820516379466
+        550.9299563468944
+ 6.23e+10    
+        549.3107794127809
+        222.2557374988154
+        498.8013136710729
+       -11.97575552648184
+        158.8078711480012
+        499.9399492156136
+       -109.4315178124881
+        -12.1775486947353
+        220.3979750597563
+        552.4669692209419
+ 6.24e+10    
+         550.843121971341
+        222.8417909636682
+        500.0710262262956
+       -12.38561826347809
+        159.1633575729938
+        501.2077690385992
+       -110.0996125652777
+       -12.58769968332899
+        220.9784499086529
+        554.0086427672576
+ 6.25e+10    
+        552.3800865214935
+         223.430938144039
+        501.3446955842593
+       -12.79501836281875
+         159.520496347743
+        502.4794765726307
+       -110.7650620592621
+       -12.99736239288079
+        221.5620207548894
+        555.5550132463272
+ 6.26e+10    
+        553.9217083635235
+        224.0232591830425
+        502.6223649796708
+       -13.20389285359848
+         159.879326689639
+         503.755113958286
+       -111.4277575636631
+        -13.4064731416055
+        222.1487681304179
+        557.1061170791444
+ 6.27e+10    
+          555.46802294954
+        224.6188349234487
+        503.9040779689673
+       -13.61217829237806
+        160.2398881443253
+        505.0347236510519
+       -112.0875897123164
+       -13.81496776792307
+         222.738773267388
+        558.6619908451294
+ 6.28e+10    
+        557.0190658814098
+        225.2177469046833
+        505.1898784294477
+       -14.01981076757121
+         160.602220584737
+        506.3183484204375
+        -112.744448516102
+       -14.22278163486839
+        223.3321180950735
+        560.2226712800465
+ 6.29e+10    
+        558.5748729086739
+        225.8200773597923
+         506.479810558384
+        -14.4267259038868
+          160.96636421012
+        507.6060313490915
+       -113.3982233755106
+       -14.62984963455561
+        223.9288852367644
+        561.7881952739024
+ 6.3e+10     
+        560.1354799264677
+        226.4259092123625
+        507.7739188721242
+       -14.83285886682138
+        161.3323595450372
+        508.8978158318988
+       -114.0488030933416
+       -15.03610619269609
+        224.5291580066166
+        563.3585998688402
+ 6.31e+10    
+        561.7009229734256
+        227.0353260734043
+        509.0722482051864
+       -15.23814436720612
+        161.7002474383544
+        510.1937455750633
+       -114.6960758875337
+       -15.44148527316938
+        225.1330204064599
+        564.9339222570322
+ 6.32e+10    
+        563.2712382295732
+        227.6484122381944
+        510.3748437093323
+       -15.64251666580269
+        162.0700690622128
+        511.4938645951852
+       -115.3399294041197
+       -15.84592038264551
+        225.7405571225693
+        566.5141997785516
+ 6.33e+10    
+        564.8464620142245
+        228.2652526830788
+        511.6817508526336
+       -16.04590957795073
+        162.4418659109834
+         512.798217218315
+       -115.9802507303069
+       -16.24934457525962
+        226.3518535223951
+        568.0994699192443
+ 6.34e+10    
+        566.4266307838594
+        228.8859330622426
+        512.9930154185297
+       -16.44825647826368
+        162.8156798002082
+        514.1068480790127
+       -116.6169264076787
+        -16.6516904573358
+        226.9669956512575
+        569.6897703085961
+ 6.35e+10    
+        568.0117811300065
+        229.5105397044372
+        514.3086835048649
+       -16.84949030537361
+        163.1915528655219
+        515.4198021193714
+       -117.2498424455131
+        -17.0528901921604
+        227.5860702290048
+        571.2851387175888
+ 6.36e+10    
+        569.6019497771058
+        230.1391596096761
+        515.6288015229267
+       -17.24954356672291
+        163.5695275615635
+        516.7371245880576
+       -117.8788843342168
+       -17.45287550480426
+          228.20916464663
+        572.8856130565433
+ 6.37e+10    
+        571.1971735803788
+        230.7718804458907
+        516.9534161964589
+       -17.64834834340276
+        163.9496466608676
+        518.0588610393145
+       -118.5039370588697
+       -17.85157768699187
+        228.8363669628593
+        574.4912313729761
+ 6.38e+10    
+        572.7974895236817
+        231.4087905455556
+        518.2825745606749
+       -18.04583629503862
+        164.3319532527434
+        519.3850573319678
+       -119.1248851128799
+       -18.24892760201765
+        229.4677659007002
+        576.1020318494263
+ 6.39e+10    
+          574.40293471736
+         232.049978902278
+        519.6163239612547
+       -18.44193866471746
+        164.7164907421395
+        520.7157596284221
+        -119.741612511742
+       -18.64485568970778
+        230.1034508439583
+        577.7180528012959
+ 6.4e+10     
+         576.013546396097
+         232.695535167353
+        520.9547120533356
+       -18.83658628396195
+        165.1033028484929
+        522.0510143936403
+       -120.3540028068985
+       -19.03929197142653
+        230.7435118337187
+        579.3393326746719
+ 6.41e+10    
+        577.6293619167521
+        233.3455496462866
+         522.297786800484
+       -19.22970957774577
+        165.4924336045636
+         523.390868394113
+       -120.9619390996999
+       -19.43216605512663
+        231.3880395647975
+        580.9659100441543
+ 6.42e+10    
+        579.2504187562058
+        234.0001132952889
+        523.6455964736674
+       -19.62123856955117
+        165.8839273552569
+        524.7353686968218
+       -121.5653040554598
+       -19.82340714044318
+        232.0371253821581
+        582.5978236106675
+ 6.43e+10    
+        580.8767545091857
+        234.6593177177328
+        524.9981896502117
+       -20.01110288646857
+        166.2778287564286
+        526.0845626681848
+       -122.1639799176029
+       -20.21294402382789
+        232.6908612772986
+        584.2351121992815
+ 6.44e+10    
+        582.5084068861019
+        235.3232551605852
+        526.3556152127471
+       -20.39923176433427
+        166.6741827736814
+        527.4384979730066
+       -122.7578485219009
+       -20.60070510372604
+        233.3493398846078
+        585.8778147570162
+ 6.45e+10    
+        584.1454137108722
+        235.9920185108067
+        527.7179223481481
+       -20.78555405290946
+        167.0730346811429
+        528.7972225734007
+       -123.3467913107955
+       -20.98661838579277
+         234.012654477693
+        587.5259703506506
+ 6.46e+10    
+        585.7878129187405
+         236.665701291721
+        529.0851605464571
+       -21.16999822109582
+        167.4744300602338
+        530.1607847277162
+       -123.9306893478022
+        -21.3706114881486
+        234.6808989656753
+        589.1796181645258
+ 6.47e+10    
+        587.4356425541089
+        237.3443976593612
+         530.457379599811
+       -21.55249236218957
+        167.8784147984219
+        531.5292329894473
+       -124.5094233319933
+       -21.75261164667267
+        235.3541678894604
+        590.8387974983436
+ 6.48e+10    
+        589.0889407683368
+        238.0282023987816
+        531.8346296013463
+       -21.93296419917046
+         168.285035087963
+        532.9026162061388
+       -125.0828736125568
+       -22.13254572033349
+        236.0325564179805
+        592.5035477649664
+ 6.49e+10    
+        590.7477458175771
+         238.717210920348
+        533.2169609441038
+       -22.31134109002724
+        168.6943374246308
+         534.280983518278
+       -125.6509202034266
+       -22.51034019655626
+        236.7161603444065
+        594.1739084882078
+ 6.5e+10     
+        592.4120960605723
+        239.4115192559989
+        534.6044243199227
+       -22.68755003311687
+        169.1063686064319
+        535.6643843581811
+       -126.2134427979816
+       -22.88592119662471
+        237.4050760823408
+        595.8499193006344
+ 6.51e+10    
+        594.0820299564747
+        240.1112240554815
+        535.9970707183182
+       -23.06151767255728
+        169.5211757323129
+        537.0528684488722
+       -126.7703207838101
+       -23.25921448111757
+        238.0994006619764
+        597.5316199413475
+ 6.52e+10    
+        595.7575860626575
+        240.8164225825652
+        537.3949514253687
+       -23.43317030365243
+        169.9388062008509
+        538.4464858029505
+       -127.3214332575363
+       -23.63014545537852
+        238.7992317262386
+        599.2190502537791
+ 6.53e+10    
+        597.4388030325164
+        241.5272127112274
+        538.7981180225777
+       -23.80243387834857
+        170.3593077089358
+        539.8452867214492
+       -127.8666590397032
+       -23.99863917501746
+        239.5046675268966
+        600.9122501834813
+ 6.54e+10    
+        599.1257196132851
+        242.2436929218192
+        540.2066223857349
+       -24.16923401072133
+        170.7827282504392
+        541.2493217926905
+       -128.4058766897121
+       -24.36462035144443
+        240.2158069206577
+        602.6112597759104
+ 6.55e+10    
+        600.8183746438398
+        242.9659622972044
+        541.6205166837686
+       -24.53349598249221
+        171.2091161148738
+        542.6586418911285
+       -128.9389645208134
+       -24.72801335743256
+         240.932749365233
+        604.3161191742169
+ 6.56e+10    
+        602.5168070525069
+        243.6941205188821
+        543.0398533775957
+       -24.89514474857258
+        171.6385198860415
+        544.0732981761932
+       -129.4658006151433
+       -25.08874223271128
+        241.6555949153861
+        606.0268686170339
+ 6.57e+10    
+        604.2210558548704
+        244.4282678630834
+         544.464685218958
+       -25.25410494263699
+        172.0709884406685
+        545.4933420911094
+       -129.9862628388069
+       -25.44673068958705
+         242.384444218958
+        607.7435484362628
+ 6.58e+10    
+        605.9311601515819
+        245.1685051968482
+        545.8950652492524
+       -25.61030088272044
+        172.5065709470346
+        546.9188253617325
+       -130.5002288570006
+        -25.8019021185922
+        243.1193985128718
+        609.4661990548627
+ 6.59e+10    
+        607.6471591261618
+        245.9149339740838
+        547.3310467983558
+       -25.96365657684399
+        172.9453168635862
+        548.3497999953522
+       -131.0075761491726
+       -26.15417959415878
+        243.8605596191183
+        611.1948609846363
+ 6.6e+10     
+        609.3690920428182
+        246.6676562316018
+        548.7726834834439
+       -26.31409572866229
+        173.3872759375449
+        549.7863182795113
+       -131.5081820242172
+       -26.50348588031967
+        244.6080299407211
+        612.9295748240226
+ 6.61e+10    
+        611.0969982442523
+        247.4267745851397
+        550.2200292078035
+       -26.66154174313577
+        173.8324982035033
+         551.228432780804
+        -132.001923635698
+       -26.84974343643209
+        245.3619124576856
+        614.6703812558832
+ 6.62e+10    
+        612.8309171494693
+        248.1923922253609
+        551.6731381596376
+       -27.00591773222571
+        174.2810339820112
+        552.6761963436746
+       -132.4886779970995
+       -27.19287442292488
+        246.1223107229291
+        616.4173210453015
+ 6.63e+10    
+        614.5708882515906
+        248.9646129138382
+        553.1320648108602
+       -27.34714652060944
+        174.7329338781537
+        554.1296620892058
+       -132.9683219971013
+        -27.5328007070697
+        246.8893288581901
+         618.170435037365
+ 6.64e+10    
+        616.3169511156773
+        249.7435409790249
+        554.5968639158984
+       -27.68515065141799
+        175.1882487801187
+         555.588883413904
+       -133.4407324148716
+       -27.86944386877059
+        247.6630715499294
+        619.9297641549712
+ 6.65e+10    
+        618.0691453765364
+         250.529281312203
+        556.0675905104715
+       -28.01985239199058
+        175.6470298577579
+        557.0539139884804
+       -133.9057859353775
+        -28.2027252063762
+        248.4436440452086
+        621.6953493966248
+ 6.66e+10    
+        619.8275107365505
+        251.3219393634214
+        557.5442999103767
+       -28.35117373965052
+        176.1093285611347
+        558.5248077566174
+       -134.3633591647071
+       -28.53256574251077
+        249.2311521475541
+        623.4672318342278
+ 6.67e+10    
+        621.5920869634938
+        252.1216211374178
+        559.0270477102672
+       -28.67903642749647
+          176.57519661907
+         560.001618933745
+       -134.8133286454028
+       -28.85888622992232
+        250.0257022128105
+        625.2454526108959
+ 6.68e+10    
+        623.3629138883597
+        252.9284331895252
+        560.5158897824227
+       -29.00336193021092
+        177.0446860376728
+        561.4844020057963
+       -135.2555708717966
+       -29.18160715734926
+        250.8274011449777
+        627.0300529387539
+ 6.69e+10    
+        625.1400314031922
+         253.742482621568
+        562.0108822755129
+       -29.32407146988481
+        177.5178490988681
+        562.9732117279656
+        -135.689962305353
+       -29.50064875540347
+        251.6363563920336
+         628.821074096753
+ 6.7e+10     
+        626.9234794589133
+        254.5638770777423
+        563.5120816133647
+       -29.64108602185499
+        177.9947383589147
+        564.4681031234674
+       -136.1163793900045
+       -29.81593100246666
+         252.452675941748
+        630.6185574284788
+ 6.71e+10    
+        628.7132980631635
+        255.3927247404869
+        565.0195444937173
+       -29.95432632055704
+        178.4754066469153
+        565.9691314822763
+       -136.5346985674877
+       -30.12737363060383
+        253.2764683174808
+        632.4225443399686
+ 6.72e+10    
+        630.5095272781358
+        256.2291343263398
+        566.5333278869761
+       -30.26371286539025
+        178.9599070633207
+         567.476352359875
+       -136.9447962926679
+       -30.43489613148819
+        254.1078425739724
+        634.2330762975317
+ 6.73e+10    
+        632.3122072184262
+        257.0732150817871
+         568.053489034957
+        -30.5691659265925
+        179.4482929784248
+        568.9898215759936
+        -137.346549048854
+       -30.73841776233794
+        254.9469082931203
+        636.0501948255755
+ 6.74e+10    
+        634.1213780488761
+        257.9250767790986
+        569.5800854496364
+       -30.87060555112837
+        179.9406180308534
+        570.5095952133412
+       -137.7398333630967
+       -31.03785755186646
+        255.7937755797491
+        637.8739415044338
+ 6.75e+10    
+        635.9370799824266
+        258.7848297121567
+        571.1131749118913
+       -31.16795156858407
+         180.436936126049
+        572.0357296163403
+       -138.1245258214694
+       -31.33313430624032
+        256.6485550573677
+        639.7043579681973
+ 6.76e+10    
+        637.7593532779774
+        259.6525846922749
+        572.6528154702322
+        -31.4611235970737
+        180.9373014347439
+        573.5682813898546
+        -138.500503084328
+        -31.6241666150485
+         257.511357863922
+        641.5414859025569
+ 6.77e+10    
+        639.5882382382451
+        260.5284530440059
+        574.1990654395432
+       -31.75004104915119
+        181.4417683914317
+        575.1073073979117
+       -138.8676419015429
+       -31.91087285727912
+        258.3822956475352
+        643.3853670426433
+ 6.78e+10    
+        641.4237752076344
+        261.4125466009467
+        575.7519833998084
+       -32.03462313772904
+        181.9503916928308
+        576.6528647624215
+       -139.2258191277054
+       -32.19317120730295
+        259.2614805622446
+        645.2360431708782
+ 6.79e+10    
+         643.266004570109
+        262.3049777015316
+         577.311628194838
+       -32.31478888200421
+        182.4632262963418
+        578.2050108619007
+       -139.5749117373001
+       -32.47097964086481
+        260.1490252637269
+        647.0935561148244
+ 6.8e+10     
+        645.1149667470698
+        263.2058591848224
+        578.8780589309948
+       -32.59045711338717
+        182.9803274184991
+         579.763803330176
+       -139.9147968398425
+       -32.74421594107845
+        261.0450429050234
+        648.9579477450537
+ 6.81e+10    
+        646.9707021952385
+        264.1153043862902
+        580.4513349759171
+       -32.86154648143515
+        183.5017505334202
+        581.3293000551065
+       -140.2453516949794
+       -33.01279770442792
+        261.9496471322534
+        650.8292599729994
+ 6.82e+10    
+        648.8332514045476
+        265.0334271335914
+        582.0315159572308
+       -33.12797545978933
+        184.0275513712441
+        582.9015591772866
+       -140.5664537275454
+        -33.2766423467705
+        262.8629520803264
+        652.7075347488408
+ 6.83e+10    
+        650.7026548960366
+        265.9603417423423
+        583.6186617612748
+       -33.38966235211146
+        184.5577859165707
+        584.4806390887543
+       -140.8779805425757
+       -33.53566710934346
+        263.7850723686485
+        654.5928140593711
+ 6.84e+10    
+        652.5789532197548
+        266.8961630118861
+        585.2128325318084
+       -33.64652529802427
+        185.0925104068913
+        586.0665984316936
+       -141.1798099402708
+       -33.78978906477142
+        264.7161230968255
+        656.4851399258894
+ 6.85e+10    
+        654.4621869526667
+        267.8410062210555
+        586.8140886687245
+        -33.8984822790492
+         185.631781331017
+         587.659496097139
+       -141.4718199309073
+       -34.03892512307468
+        265.6562198403618
+        658.3845544020853
+ 6.86e+10    
+        656.3523966965699
+        268.7949871239364
+        588.4224908267624
+       -34.14545112454591
+        186.1756554275002
+        589.2593912236714
+       -141.7538887496986
+       -34.28299203767762
+        266.6054786463567
+        660.2910995719391
+ 6.87e+10    
+        658.2496230760185
+        269.7582219456252
+         590.038099914213
+       -34.38734951764675
+        186.7241896830564
+        590.8663431961237
+       -142.0258948715928
+       -34.52190641141528
+        267.5640160291991
+        662.2048175476248
+ 6.88e+10    
+        660.1539067362456
+        270.7308273779845
+        591.6609770916251
+       -34.62409500119108
+        187.2774413309755
+        592.4804116442642
+       -142.2877170260123
+       -34.75558470253715
+        268.5319489662598
+        664.1257504674215
+ 6.89e+10    
+        662.0652883411078
+        271.7129205753989
+        593.2911837705127
+       -34.85560498365452
+        187.8354678495367
+        594.1016564415052
+       -142.5392342115295
+       -34.98394323070887
+        269.5093948935845
+        666.0539404936337
+ 6.9e+10     
+        663.9838085710218
+         272.704619150529
+         594.928781612057
+       -35.08179674507382
+         188.398326960415
+        595.7301377035916
+       -142.7803257104745
+       -35.20689818300968
+        270.4964717015811
+        667.9894298105131
+ 6.91e+10    
+        665.9095081209157
+        273.7060411700634
+        596.5738325258097
+       -35.30258744296597
+         188.966076627085
+        597.3659157872893
+       -143.0108711034721
+        -35.4243656199235
+        271.4932977307158
+        669.9322606221978
+ 6.92e+10    
+        667.8424276981909
+        274.7173051504741
+         598.226398668396
+       -35.51789411824144
+        189.5387750532233
+        599.0090512890821
+       -143.2307502839076
+       -35.63626148132622
+        272.4999917671996
+        671.8824751506462
+ 6.93e+10    
+        669.7826080206826
+        275.7385300537684
+        599.8865424422111
+       -35.72763370110916
+        190.1164806811083
+        600.6596050438592
+       -143.4398434723142
+       -35.84250159246422
+        273.5166730386833
+        673.8401156335904
+ 6.94e+10    
+        671.7300898146359
+        276.7698352832456
+         601.554326494124
+        -35.9317230169742
+        190.6992521900132
+        602.3176381236055
+       -143.6380312306829
+       -36.04300166992591
+         274.543461209951
+        675.8052243224943
+ 6.95e+10    
+        673.6849138126897
+        277.8113406792535
+        603.2298137141798
+       -36.13007879232513
+        191.2871484946034
+        603.9832118360955
+       -143.8251944766903
+       -36.23767732760516
+        275.5804763786166
+        677.7778434805126
+ 6.96e+10    
+        675.6471207518566
+        278.8631665149464
+        604.9130672342915
+       -36.32261766061264
+        191.8802287433243
+        605.6563877235752
+       -144.0012144978395
+       -36.42644408265398
+          276.62783907082
+        679.7580153804676
+ 6.97e+10    
+        677.6167513715341
+        279.9254334920452
+        606.6041504269446
+        -36.5092561681164
+         192.478552316793
+        607.3372275614564
+       -144.1659729655173
+       -36.60921736142613
+        277.6856702369305
+        681.7457823028307
+ 6.98e+10    
+        679.5938464114988
+        280.9982627366059
+        608.3031269038962
+       -36.68991077980066
+        193.0821788261845
+        609.0257933570003
+       -144.3193519489564
+       -36.78591250540808
+        278.7540912472517
+        683.7411865337097
+ 6.99e+10    
+        681.5784466099258
+        282.0817757947825
+        610.0100605148705
+       -36.86449788515687
+        193.6911681116172
+        610.7221473480141
+        -144.461233929108
+       -36.95644477713918
+        279.8332238877294
+        685.7442703628475
+ 7e+10       
+        683.5705927014085
+        283.1760946286022
+        611.7250153462609
+       -37.03293380403266
+        194.3055802405381
+        612.4263520015319
+       -144.5915018124156
+       -37.12072936611767
+        280.9231903556666
+        687.7550760816317
* NOTE: Solution at 1e+08 Hz used as DC point.

.model l_m4lines_port_1 sp N=4 SPACING=nonuniform VALTYPE=real
+ INTERPOLATION=spline
+ INFINITY =
+    4.750572009209595e-07
+    2.002860793599409e-07
+    4.579454404695213e-07
+     6.37920267040962e-08
+    1.290978198905292e-07
+    4.575299532832819e-07
+    2.841009207981307e-08
+    6.374627613487148e-08
+    2.005831724691381e-07
+    4.751237083519819e-07
+ DATA = 700
+ 0           
+    4.161185452528795e-07
+    1.501129145652629e-07
+    4.133044816583034e-07
+    4.576475473155456e-08
+     9.33984140372853e-08
+    4.128254273149257e-07
+    2.492636456251042e-08
+    4.585388542163275e-08
+    1.505121816752186e-07
+    4.160184534840582e-07
+ 2e+08       
+    4.124674982773361e-07
+    1.498111269492382e-07
+    4.095935298607717e-07
+    4.567127792791265e-08
+    9.295302755871797e-08
+    4.090985011578709e-07
+    2.490601859685072e-08
+    4.576060695980833e-08
+    1.502229064519691e-07
+    4.123714896777287e-07
+ 3e+08       
+    4.107955828678745e-07
+    1.496806833958028e-07
+    4.079106636739773e-07
+    4.561664417113724e-08
+    9.275924621976011e-08
+    4.074090367227649e-07
+    2.488877489633768e-08
+    4.570548968373417e-08
+    1.500965059173988e-07
+    4.106993511407159e-07
+ 4e+08       
+    4.098446379977531e-07
+     1.49630887889878e-07
+    4.069532541220837e-07
+    4.558967803829978e-08
+    9.265390254351089e-08
+    4.064469168355302e-07
+    2.488286615191472e-08
+     4.56782713104685e-08
+    1.500494299889396e-07
+    4.097475895375576e-07
+ 5e+08       
+    4.091894057447739e-07
+    1.495965094554214e-07
+    4.062929526449319e-07
+    4.557360608608974e-08
+    9.258195650188645e-08
+    4.057828010897483e-07
+    2.488063100206433e-08
+    4.566206802954512e-08
+    1.500172999314607e-07
+    4.090914134825178e-07
+ 6e+08       
+    4.086904070749359e-07
+    1.495663700273411e-07
+    4.057905376850967e-07
+    4.556228585534797e-08
+    9.252733939933493e-08
+    4.052772836251412e-07
+     2.48792563611113e-08
+    4.565065125983407e-08
+    1.499889823442598e-07
+    4.085914211836883e-07
+ 7e+08       
+    4.082929694905094e-07
+    1.495404975525814e-07
+    4.053912200764045e-07
+    4.555361973622064e-08
+    9.248421046569685e-08
+     4.04875497898638e-07
+    2.487812154905077e-08
+    4.564189507479129e-08
+    1.499645919522025e-07
+    4.081929975207392e-07
+ 8e+08       
+    4.079692620040247e-07
+    1.495194200504797e-07
+    4.050666072305823e-07
+    4.554680649429544e-08
+    9.244953393711487e-08
+    4.045489169388144e-07
+    2.487725177487061e-08
+    4.563499467757789e-08
+    1.499447457797467e-07
+     4.07868348888434e-07
+ 9e+08       
+    4.077014515086331e-07
+    1.495027383425224e-07
+    4.047981432627704e-07
+    4.554144658534555e-08
+      9.2421227222706e-08
+    4.042787933542984e-07
+    2.487678339382288e-08
+    4.562955463272481e-08
+    1.499291049035168e-07
+    4.075996574219543e-07
+ 1e+09       
+    4.074765492396635e-07
+    1.494894836481794e-07
+    4.045721593763728e-07
+    4.553727075769961e-08
+     9.23976961099218e-08
+     4.04051245434181e-07
+    2.487681883883212e-08
+    4.562531108731319e-08
+     1.49916733917596e-07
+    4.073739346510244e-07
+ 1.1e+09     
+    4.072750426808511e-07
+    1.494829776718474e-07
+    4.043705915550338e-07
+    4.554007612947905e-08
+    9.238698836550983e-08
+    4.038476415211274e-07
+    2.487954351449982e-08
+    4.562794177509821e-08
+    1.499087713052823e-07
+    4.071712125605106e-07
+ 1.2e+09     
+    4.070934453823108e-07
+    1.494761713065997e-07
+    4.041883396601975e-07
+    4.554232276209583e-08
+     9.23759407379601e-08
+    4.036636249285331e-07
+    2.488256994769246e-08
+    4.563003220589512e-08
+    1.499011653337313e-07
+    4.069885611639511e-07
+ 1.3e+09     
+     4.06931002298291e-07
+    1.494694626780808e-07
+    4.040248466941724e-07
+    4.554407163035181e-08
+    9.236490159675793e-08
+    4.034986125539983e-07
+    2.488580410576813e-08
+    4.563164117621565e-08
+    1.498941489485369e-07
+     4.06825201451716e-07
+ 1.4e+09     
+    4.067863617488966e-07
+    1.494631310662023e-07
+    4.038789337365786e-07
+    4.554539452169479e-08
+    9.235413620630198e-08
+    4.033514009410969e-07
+      2.4889148462016e-08
+    4.563283861843677e-08
+    1.498878670551993e-07
+    4.066797606690226e-07
+ 1.5e+09     
+    4.066578724953411e-07
+    1.494573581659914e-07
+    4.037490906196623e-07
+    4.554636918414288e-08
+    9.234383822925318e-08
+     4.03220457571746e-07
+    2.489251136985221e-08
+    4.563370060433711e-08
+    1.498823962715307e-07
+    4.065505696513779e-07
+ 1.6e+09     
+    4.065437866894425e-07
+    1.494522521741015e-07
+    4.036336779846842e-07
+    4.554707634359468e-08
+     9.23341441615189e-08
+    4.031041227697645e-07
+    2.489581464126434e-08
+    4.563430625620271e-08
+    1.498777648454504e-07
+    4.064358655059405e-07
+ 1.7e+09     
+     4.06442389811746e-07
+    1.494478697711686e-07
+    4.035310595169822e-07
+    4.554759789694662e-08
+    9.232514732978937e-08
+    4.030007415363164e-07
+    2.489899902698746e-08
+     4.56347358845373e-08
+    1.498739698212263e-07
+    4.063339211060429e-07
+ 1.8e+09     
+    4.063520774479294e-07
+    1.494442340501823e-07
+    4.034396826076147e-07
+    4.554801579599741e-08
+    9.231690992970876e-08
+    4.029087438174014e-07
+    2.490202754028625e-08
+    4.563506985750382e-08
+    1.498709904710619e-07
+    4.062431214176051e-07
+ 1.9e+09     
+    4.062713952544132e-07
+    1.494413480848632e-07
+    4.033581227684211e-07
+    4.554841130425799e-08
+    9.230947265327252e-08
+    4.028266886259239e-07
+    2.490488674877557e-08
+    4.563538786897467e-08
+    1.498687980578901e-07
+    4.061620030754235e-07
+ 2e+09       
+    4.061990545836646e-07
+    1.494392046047644e-07
+    4.032851036648791e-07
+    4.554886443349851e-08
+    9.230286200127233e-08
+    4.027532838990365e-07
+    2.490758629343015e-08
+     4.56357683986952e-08
+    1.498673624638122e-07
+    4.060892696960652e-07
+ 2.1e+09     
+    4.061339327967622e-07
+    1.494377925161939e-07
+    4.032195014698288e-07
+    4.554945345498901e-08
+     9.22970956101784e-08
+    4.026873907763268e-07
+     2.49101569843789e-08
+    4.563628825017434e-08
+    1.498666563550123e-07
+    4.060237919491868e-07
+ 2.2e+09     
+    4.060750645433125e-07
+    1.494371010249528e-07
+    4.031603396726735e-07
+    4.555025443900841e-08
+    9.229218598579834e-08
+    4.026280184063686e-07
+    2.491264786927643e-08
+    4.563702211428777e-08
+    1.498666575239546e-07
+    4.059645986542819e-07
+ 2.3e+09     
+    4.060216282295995e-07
+    1.494371220223738e-07
+    4.031067785271397e-07
+    4.555134081201232e-08
+     9.22881430158708e-08
+    4.025743134389917e-07
+    2.491512267385752e-08
+    4.563804214521034e-08
+    1.498673499510773e-07
+    4.059108631100865e-07
+ 2.4e+09     
+    4.059729304163215e-07
+    1.494378512672061e-07
+    4.030581019014075e-07
+    4.555278293984946e-08
+    9.228497557973232e-08
+    4.025255469467247e-07
+    2.491765598174908e-08
+    4.563941755614275e-08
+    1.498687240130369e-07
+     4.05861887386363e-07
+ 2.5e+09     
+    4.059283898571924e-07
+    1.494392887695671e-07
+    4.030137032945636e-07
+    4.555464775276527e-08
+    9.228269251102242e-08
+    4.024811005247314e-07
+    2.492032946158123e-08
+    4.564121425073501e-08
+    1.498707761572994e-07
+    4.058170862803229e-07
+ 2.6e+09     
+    4.058875221911141e-07
+    1.494414386745352e-07
+    4.029730720965088e-07
+    4.555699842790502e-08
+    9.228130311111847e-08
+    4.024404526364661e-07
+    2.492322837563499e-08
+    4.564349450665869e-08
+    1.498735082728703e-07
+    4.057759719438044e-07
+ 2.7e+09     
+    4.058499258384376e-07
+    1.494443088559141e-07
+    4.029357807072766e-07
+    4.555989414098273e-08
+    9.228081736133069e-08
+    4.024031658143712e-07
+    2.492643852701067e-08
+    4.564631672397824e-08
+    1.498769269159205e-07
+    4.057381397270539e-07
+ 2.8e+09     
+     4.05815269354066e-07
+    1.494479103641072e-07
+    4.029014728290143e-07
+    4.556338989315107e-08
+    9.228124594181568e-08
+    4.023688750242667e-07
+    2.493004373073263e-08
+    4.564973524539826e-08
+    1.498810424953335e-07
+    4.057032554886147e-07
+ 2.9e+09     
+    4.057832803044905e-07
+    1.494522568227825e-07
+    4.028698530504143e-07
+    4.556753641349554e-08
+    9.228260013397902e-08
+    4.023372773096058e-07
+    2.493412383434096e-08
+    4.565380024980693e-08
+    1.498858684838919e-07
+    4.056710444361654e-07
+ 3e+09       
+     4.05753735625172e-07
+    1.494573638335853e-07
+    4.028406777238736e-07
+    4.557238013289281e-08
+    9.228489165949003e-08
+    4.023081227127073e-07
+    2.493875326820777e-08
+    4.565855771575648e-08
+    1.498914206929138e-07
+    4.056412814531665e-07
+ 3.1e+09     
+      4.0572645335335e-07
+    1.494632484233607e-07
+    4.028137470655274e-07
+    4.557796322160772e-08
+     9.22881324914801e-08
+    4.022812064000297e-07
+    2.494400007526784e-08
+    4.566404944803795e-08
+    1.498977166289473e-07
+    4.056137828052533e-07
+ 3.2e+09     
+    4.057012856016089e-07
+    1.494699285514418e-07
+    4.027888983705665e-07
+    4.558432368098457e-08
+    9.229233466071792e-08
+    4.022563618809203e-07
+    2.494992535246985e-08
+    4.567031315836564e-08
+    1.499047749383752e-07
+    4.055883990908814e-07
+ 3.3e+09     
+    4.056781126276432e-07
+    1.494774226834329e-07
+    4.027660002194031e-07
+    4.559149547875243e-08
+    9.229751007044374e-08
+    4.022334551926934e-07
+    2.495658302946121e-08
+    4.567738259022529e-08
+    1.499126149377243e-07
+    4.055650092910077e-07
+ 3.4e+09     
+    4.056568378576177e-07
+    1.494857494308877e-07
+    4.027449475466053e-07
+     4.55995087175447e-08
+    9.230367032720513e-08
+    4.022123799218079e-07
+    2.496401991095026e-08
+    4.568528767789772e-08
+      1.4992125622273e-07
+    4.055435157746471e-07
+ 3.5e+09     
+    4.056373837292035e-07
+    1.494949272521352e-07
+     4.02725657448968e-07
+    4.560838982695698e-08
+     9.23108265907757e-08
+    4.021930529362992e-07
+    2.497227591516665e-08
+     4.56940547302743e-08
+    1.499307183467947e-07
+    4.055238401259371e-07
+ 3.6e+09     
+    4.056196882324408e-07
+    1.495049742073368e-07
+    4.027080656182693e-07
+    4.561816177058461e-08
+     9.23189894435156e-08
+    4.021754107150559e-07
+    2.498138444962609e-08
+    4.570370663108243e-08
+    1.499410205586292e-07
+    4.055059196704332e-07
+ 3.7e+09     
+    4.056037020399695e-07
+    1.495159077600046e-07
+    4.026921232960331e-07
+    4.562884426079469e-08
+    9.232816877794058e-08
+    4.021594061728898e-07
+    2.499137287530321e-08
+    4.571426304834057e-08
+    1.499521815890606e-07
+    4.054897045918114e-07
+ 3.8e+09     
+    4.055893861315765e-07
+    1.495277446172376e-07
+    4.026777946605917e-07
+    4.564045397534684e-08
+     9.23383737004885e-08
+    4.021450058949781e-07
+     2.50022630201527e-08
+    4.572574064712166e-08
+    1.499642194778207e-07
+    4.054751555436008e-07
+ 3.9e+09     
+     4.05576709830821e-07
+    1.495405006014836e-07
+    4.026650545699623e-07
+    4.565300477128693e-08
+    9.234961244926299e-08
+    4.021321877091918e-07
+    2.501407171196614e-08
+    4.573815330092031e-08
+    1.499771514323435e-07
+    4.054622416734067e-07
+ 4e+09       
+    4.055656491831899e-07
+    1.495541905475092e-07
+    4.026538865969751e-07
+    4.566650789272925e-08
+    9.236189232370761e-08
+    4.021209385392135e-07
+    2.502681130842313e-08
+    4.575151229803588e-08
+    1.499909937119624e-07
+    4.054509389888493e-07
+ 4.1e+09     
+    4.055561856158301e-07
+    1.495688282192806e-07
+    4.026442813052376e-07
+    4.568097217018552e-08
+     9.23752196245589e-08
+    4.021112524946109e-07
+    2.504049020875857e-08
+     4.57658265403697e-08
+    1.500057615322985e-07
+    4.054412290050581e-07
+ 4.2e+09     
+    4.055483048282214e-07
+    1.495844262425275e-07
+    4.026362347256519e-07
+    4.569640420997545e-08
+    9.238959960293357e-08
+    4.021031291657396e-07
+    2.505511333673841e-08
+    4.578110273287683e-08
+    1.500214689859357e-07
+    4.054330976229459e-07
+ 4.3e+09     
+     4.05541995871357e-07
+    1.496009960497765e-07
+    4.026297470030284e-07
+    4.571280857296464e-08
+     9.24050364179228e-08
+    4.020965721011786e-07
+    2.507068258873489e-08
+    4.579734556261361e-08
+    1.500381289766395e-07
+    4.054265341957455e-07
+ 4.4e+09     
+    4.055372503801157e-07
+    1.496185478355845e-07
+    4.026248211907683e-07
+    4.573018794242464e-08
+    9.242153310252653e-08
+    4.020915874531292e-07
+    2.508719724377728e-08
+    4.581455786688578e-08
+    1.500557531653296e-07
+    4.054215307484615e-07
+ 4.5e+09     
+    4.055340619296817e-07
+    1.496370905204957e-07
+    4.026214621784685e-07
+    4.574854328121609e-08
+    9.243909153811975e-08
+    4.020881827818803e-07
+    2.510465433469808e-08
+    4.583274079044266e-08
+    1.500743519267562e-07
+    4.054180813211169e-07
+ 4.6e+09     
+    4.055324254921641e-07
+    1.496566317228981e-07
+    4.026196757426222e-07
+    4.576787397877099e-08
+    9.245771243786534e-08
+      4.0208636601403e-07
+    2.512304898106732e-08
+    4.585189393199003e-08
+    1.500939343163486e-07
+    4.054161814120238e-07
+ 4.7e+09     
+    4.055323369741378e-07
+    1.496771777384543e-07
+    4.026194677144147e-07
+    4.578817798851677e-08
+    9.247739533957554e-08
+    4.020861445509344e-07
+    2.514237468565431e-08
+    4.587201548052631e-08
+    1.501145080470107e-07
+     4.05415827501927e-07
+ 4.8e+09     
+    4.055337928197046e-07
+    1.496987335271088e-07
+    4.026208432609643e-07
+     4.58094519564637e-08
+    9.249813860847746e-08
+    4.020875245241307e-07
+    2.516262359680617e-08
+    4.589310234215198e-08
+     1.50136079475779e-07
+    4.054170166437733e-07
+ 4.9e+09     
+    4.055367896669856e-07
+    1.497213027078777e-07
+    4.026238062775255e-07
+    4.583169134168692e-08
+    9.251993945018089e-08
+    4.020905101935461e-07
+     2.51837867394896e-08
+    4.591515025808089e-08
+     1.50158653600247e-07
+    4.054197461062135e-07
+ 5e+09       
+    4.055413240487434e-07
+    1.497448875616925e-07
+    4.026283588882504e-07
+    4.585489052939811e-08
+    9.254279393390994e-08
+    4.020951034826628e-07
+     2.52058542178881e-08
+    4.593815391460371e-08
+    1.501822340645661e-07
+    4.054240130617367e-07
+ 5.1e+09     
+     4.05547392130136e-07
+    1.497694890425422e-07
+    4.026345010524247e-07
+     4.58790429372328e-08
+    9.256669702577156e-08
+     4.02101303642736e-07
+    2.522881539244713e-08
+    4.596210704573284e-08
+    1.502068231746641e-07
+    4.054298143126496e-07
+ 5.2e+09     
+    4.055549894785421e-07
+    1.497951067970597e-07
+    4.026422302718993e-07
+    4.590414111529778e-08
+    9.259164263153469e-08
+    4.021091070360828e-07
+    2.525265903416191e-08
+    4.598700252920934e-08
+    1.502324219221502e-07
+    4.054371460500346e-07
+ 5.3e+09     
+    4.055641108619015e-07
+    1.498217391925518e-07
+    4.026515413939704e-07
+    4.593017684043615e-08
+    9.261762364810955e-08
+    4.021185070265973e-07
+    2.527737345874283e-08
+     4.60128324764827e-08
+    1.502590300162013e-07
+    4.054460036423097e-07
+ 5.4e+09     
+    4.055747500732396e-07
+    1.498493833533022e-07
+    4.026624265024492e-07
+    4.595714120508808e-08
+    9.264463202266836e-08
+    4.021294939642206e-07
+     2.53029466430994e-08
+     4.60395883171972e-08
+    1.502866459225872e-07
+    4.054563814511968e-07
+ 5.5e+09     
+    4.055868997799314e-07
+    1.498780352048104e-07
+    4.026748748883091e-07
+    4.598502470105461e-08
+      9.2672658818164e-08
+    4.021420552492275e-07
+    2.532936632636984e-08
+    4.606726087863839e-08
+    1.503152669089012e-07
+    4.054682726737545e-07
+ 5.6e+09     
+     4.05600551396907e-07
+    1.499076895254732e-07
+    4.026888730902417e-07
+    4.601381729841835e-08
+    9.270169428388035e-08
+    4.021561754618916e-07
+    2.535662009750804e-08
+    4.609584046051993e-08
+    1.503448890950148e-07
+    4.054816692097266e-07
+ 5.7e+09     
+    4.056156949833931e-07
+    1.499383400050837e-07
+    4.027044049947201e-07
+     4.60435085198313e-08
+    9.273172792959344e-08
+     4.02171836543346e-07
+    2.538469547122522e-08
+     4.61253169054224e-08
+    1.503755075077845e-07
+    4.054965615538005e-07
+ 5.8e+09     
+    4.056323191630021e-07
+    1.499699793094224e-07
+    4.027214519848954e-07
+    4.607408751035412e-08
+     9.27627486019352e-08
+    4.021890180142275e-07
+    2.541357995388075e-08
+    4.615567966514089e-08
+    1.504071161390826e-07
+    4.055129387125279e-07
+ 5.9e+09     
+    4.056504110670012e-07
+    1.500025991501467e-07
+    4.027399931277402e-07
+    4.610554310301296e-08
+    9.279474456162008e-08
+    4.022076972188239e-07
+    2.544326110072455e-08
+    4.618691786315308e-08
+     1.50439708006309e-07
+    4.055307881456548e-07
+ 6e+09       
+    4.056699563005187e-07
+    1.500361903591441e-07
+    4.027600053892951e-07
+    4.613786388023163e-08
+    9.282770356030321e-08
+    4.022278495838356e-07
+    2.547372656571658e-08
+    4.621902035338422e-08
+    1.504732752146386e-07
+    4.055500957314572e-07
+ 6.1e+09     
+    4.056909389312295e-07
+    1.500707429664974e-07
+    4.027814638686396e-07
+     4.61710382312942e-08
+     9.28616129159886e-08
+    4.022494488824605e-07
+    2.550496414498726e-08
+    4.625197577542347e-08
+    1.505078090203848e-07
+     4.05570845755478e-07
+ 6.2e+09     
+    4.057133414998163e-07
+    1.501062462812248e-07
+    4.028043420421418e-07
+    4.620505440599282e-08
+    9.289645958606643e-08
+    4.022724674961074e-07
+    2.553696181485562e-08
+    4.628577260632788e-08
+    1.505432998949709e-07
+    4.055930209217581e-07
+ 6.3e+09     
+    4.057371450511932e-07
+     1.50142688973968e-07
+    4.028286120106842e-07
+    4.623990056461802e-08
+    9.293223023723527e-08
+     4.02296876667652e-07
+    2.556970776519073e-08
+    4.632039920914307e-08
+    1.505797375891275e-07
+    4.056166023853682e-07
+ 6.4e+09     
+    4.057623291851705e-07
+    1.501800591608463e-07
+     4.02854244743686e-07
+    4.627556482444854e-08
+    9.296891131173298e-08
+    4.023226467416278e-07
+    2.560319042878448e-08
+    4.635584387826354e-08
+    1.506171111970359e-07
+    4.056415698047224e-07
+ 6.5e+09     
+    4.057888721249456e-07
+    1.502183444877216e-07
+    4.028812103149567e-07
+     4.63120353028995e-08
+    9.300648908946769e-08
+    4.023497473881087e-07
+    2.563739850730079e-08
+    4.639209488175577e-08
+    1.506554092202389e-07
+    4.056679014118997e-07
+ 6.6e+09     
+    4.058167508015307e-07
+    1.502575322141733e-07
+     4.02909478126515e-07
+    4.634930015748495e-08
+    9.304494974578593e-08
+    4.023781478082048e-07
+    2.567232099427624e-08
+    4.642914050076761e-08
+    1.506946196312186e-07
+    4.056955740989463e-07
+ 6.7e+09     
+    4.058459409520161e-07
+    1.502976092965129e-07
+    4.029390171175572e-07
+    4.638734762274847e-08
+    9.308427940474724e-08
+    4.024078169200891e-07
+    2.570794719556802e-08
+    4.646696906614917e-08
+    1.507347299366067e-07
+    4.057245635179481e-07
+ 6.8e+09     
+    4.058764172294032e-07
+    1.503385624692257e-07
+    4.029697959566716e-07
+    4.642616604431009e-08
+    9.312446418788376e-08
+    4.024387235252814e-07
+     2.57442667475795e-08
+    4.650556899241272e-08
+    1.507757272400473e-07
+    4.057548441925562e-07
+ 6.9e+09     
+    4.059081533216461e-07
+    1.503803783242562e-07
+    4.030017832162049e-07
+    4.646574391017284e-08
+    9.316549025851692e-08
+    4.024708364555474e-07
+    2.578126963353544e-08
+    4.654492880916057e-08
+    1.508175983047622e-07
+    4.057863896385814e-07
+ 7e+09       
+    4.059411220774994e-07
+    1.504230433876102e-07
+    4.030349475283434e-07
+    4.650606987942439e-08
+    9.320734386177116e-08
+     4.02504124701244e-07
+    2.581894619803236e-08
+    4.658503719011012e-08
+    1.508603296158949e-07
+    4.058191724912845e-07
+ 7.1e+09     
+      4.0597529563681e-07
+    1.504665441927818e-07
+    4.030692577230099e-07
+    4.654713280846355e-08
+    9.325001136048059e-08
+    4.025385575222799e-07
+    2.585728716004935e-08
+    4.662588297984634e-08
+    1.509039074427179e-07
+    4.058531646370687e-07
+ 7.2e+09     
+    4.060106455629624e-07
+    1.505108673505608e-07
+    4.031046829480907e-07
+    4.658892177487367e-08
+    9.329347926721983e-08
+    4.025741045430751e-07
+     2.58962836245728e-08
+    4.666745521842838e-08
+    1.509483179007844e-07
+    4.058883373473818e-07
+ 7.3e+09     
+    4.060471429753422e-07
+    1.505559996148284e-07
+    4.031411927728246e-07
+    4.663142609905908e-08
+    9.333773427271516e-08
+      4.0261073583302e-07
+    2.593592709296222e-08
+    4.670974316397706e-08
+    1.509935470140936e-07
+    4.059246614128194e-07
+ 7.4e+09     
+      4.0608475867984e-07
+    1.506019279439872e-07
+    4.031787572753918e-07
+     4.66746353637538e-08
+    9.338276327090204e-08
+    4.026484219739771e-07
+    2.597620947216364e-08
+    4.675273631336394e-08
+    1.510395807773173e-07
+    4.059621072756021e-07
+ 7.5e+09     
+    4.061234632956512e-07
+     1.50648639557735e-07
+      4.0321734711588e-07
+    4.671853943150861e-08
+    9.342855338090053e-08
+    4.026871341163489e-07
+    2.601712308286077e-08
+     4.67964244211193e-08
+    1.510864052181012e-07
+    4.060006451588214e-07
+ 7.6e+09     
+    4.061632273768335e-07
+    1.506961219889353e-07
+    4.032569335958794e-07
+    4.676312846025545e-08
+    9.347509196617166e-08
+     4.02726844025166e-07
+    2.605866066664132e-08
+    4.684079751667044e-08
+    1.511340064594199e-07
+    4.060402451910829e-07
+ 7.7e+09     
+    4.062040215273558e-07
+    1.507443631304012e-07
+    4.032974887059797e-07
+    4.680839291704727e-08
+    9.352236665111109e-08
+    4.027675241175539e-07
+    2.610081539224645e-08
+    4.688584592001437e-08
+     1.51182370781915e-07
+    4.060808775254046e-07
+ 7.8e+09     
+    4.062458165085974e-07
+    1.507933512764616e-07
+    4.033389851624266e-07
+    4.685432359006642e-08
+    9.357036533532058e-08
+    4.028091474928249e-07
+    2.614358086096326e-08
+    4.693156025592245e-08
+    1.512314846860956e-07
+    4.061225124514537e-07
+ 7.9e+09     
+    4.062885833385163e-07
+    1.508430751592366e-07
+    4.033813964341393e-07
+    4.690091159899328e-08
+    9.361907620577898e-08
+    4.028516879562908e-07
+    2.618695111121498e-08
+     4.69779314667651e-08
+    1.512813349542247e-07
+    4.061651205004209e-07
+ 8e+09       
+    4.063322933819314e-07
+    1.508935239796145e-07
+    4.034246967612531e-07
+    4.694814840382548e-08
+    9.366848774712257e-08
+    4.028951200377851e-07
+    2.623092062239917e-08
+    4.702495082403835e-08
+     1.51331908711658e-07
+    4.062086725420414e-07
+ 8.1e+09     
+    4.063769184315786e-07
+    1.509446874329649e-07
+      4.0346886116624e-07
+    4.699602581223456e-08
+     9.37185887502164e-08
+    4.029394190057164e-07
+    2.627548431802013e-08
+    4.707260993866201e-08
+     1.51383193487337e-07
+    4.062531398734266e-07
+ 8.2e+09     
+    4.064224307798099e-07
+    1.509965557296933e-07
+    4.035138654586006e-07
+    4.704453598554802e-08
+    9.376936831918816e-08
+    4.029845608773693e-07
+     2.63206375681595e-08
+    4.712090077011286e-08
+    1.514351772730843e-07
+    4.062984942995492e-07
+ 8.3e+09     
+    4.064688032809642e-07
+    1.510491196107826e-07
+    4.035596862340378e-07
+    4.709367144344115e-08
+    9.382081587707225e-08
+    4.030305224260249e-07
+    2.636637619132635e-08
+    4.716981563444638e-08
+    1.514878485812893e-07
+    4.063447082053425e-07
+ 8.4e+09     
+    4.065160094046032e-07
+    1.511023703585193e-07
+    4.036063008689114e-07
+    4.714342506742312e-08
+    9.387292117019556e-08
+    4.030772811853672e-07
+    2.641269645572596e-08
+    4.721934721125105e-08
+    1.515411965005232e-07
+    4.063917546194892e-07
+ 8.5e+09     
+    4.065640232799267e-07
+    1.511562998026445e-07
+    4.036536875107251e-07
+     4.71937901031997e-08
+    9.392567427142235e-08
+    4.031248154515428e-07
+    2.645959507998445e-08
+    4.726948854957265e-08
+    1.515952107485765e-07
+    4.064396072700609e-07
+ 8.6e+09     
+    4.066128197317816e-07
+    1.512109003222048e-07
+    4.037018250652889e-07
+    4.724476016199305e-08
+    9.397906558235657e-08
+    4.031731042831332e-07
+    2.650706923336505e-08
+    4.732023307283769e-08
+    1.516498817223801e-07
+    4.064882406322407e-07
+ 8.7e+09     
+    4.066623743087717e-07
+     1.51266164843413e-07
+    4.037506931811552e-07
+    4.729632922089847e-08
+    9.403308583459257e-08
+    4.032221274992401e-07
+    2.655511653550972e-08
+     4.73715745827992e-08
+    1.517052005442479e-07
+    4.065376299684061e-07
+ 8.8e+09     
+    4.067126633040172e-07
+    1.513220868338507e-07
+    4.038002722318362e-07
+    4.734849162235426e-08
+    9.408772609008717e-08
+    4.032718656758019e-07
+    2.660373505573906e-08
+    4.742350726252293e-08
+    1.517611591038696e-07
+    4.065877513608937e-07
+ 8.9e+09     
+     4.06763663769168e-07
+    1.513786602933626e-07
+    4.038505432962634e-07
+    4.740124207279995e-08
+     9.41429777407212e-08
+    4.033223001402152e-07
+    2.665292331194149e-08
+    4.747602567842821e-08
+    1.518177500954894e-07
+    4.066385817377843e-07
+ 9e+09       
+    4.068153535222893e-07
+    1.514358797420088e-07
+    4.039014881378967e-07
+    4.745457564059558e-08
+    9.419883250710815e-08
+    4.033734129642953e-07
+    2.670268026908274e-08
+    4.752912478139572e-08
+    1.518749670497301e-07
+    4.066900988920678e-07
+ 9.1e+09     
+    4.068677111502479e-07
+     1.51493740205441e-07
+    4.039530891828273e-07
+    4.750848775327178e-08
+    9.425528243670033e-08
+    4.034251869555694e-07
+    2.675300533736518e-08
+    4.758279990695371e-08
+    1.519328043595587e-07
+    4.067422814945568e-07
+ 9.2e+09     
+    4.069207160062218e-07
+    1.515522371980734e-07
+    4.040053294971889e-07
+    4.756297419417847e-08
+    9.431231990123951e-08
+    4.034776056468982e-07
+    2.680389837006687e-08
+     4.76370467745547e-08
+    1.519912572999497e-07
+     4.06795109100913e-07
+ 9.3e+09     
+    4.069743482029453e-07
+    1.516113667044123e-07
+    4.040581927641414e-07
+    4.761803109859719e-08
+    9.436993759359372e-08
+    4.035306532843972e-07
+    2.685535966109021e-08
+    4.769186148595802e-08
+    1.520503220408702e-07
+      4.0684856215317e-07
+ 9.4e+09     
+    4.070285886022654e-07
+    1.516711251588945e-07
+     4.04111663260661e-07
+    4.767365494937947e-08
+    9.442812852402021e-08
+    4.035843148136416e-07
+    2.690738994225006e-08
+    4.774724052273673e-08
+    1.521099956533011e-07
+    4.069026219761189e-07
+ 9.5e+09     
+    4.070834188015754e-07
+    1.517315094245755e-07
+    4.041657258343326e-07
+    4.772984257217139e-08
+    9.448688601589308e-08
+    4.036385758641447e-07
+     2.69599903803329e-08
+    4.780318074293328e-08
+    1.521702761081067e-07
+    4.069572707689414e-07
+ 9.6e+09     
+    4.071388211176375e-07
+    1.517925167709856e-07
+    4.042203658803196e-07
+    4.778659113028162e-08
+    9.454620370093383e-08
+    4.036934227321202e-07
+    2.701316257395853e-08
+    4.785967937689413e-08
+    1.522311622676714e-07
+    4.070124915924582e-07
+ 9.7e+09     
+    4.071947785682723e-07
+    1.518541448514523e-07
+    4.042755693186501e-07
+    4.784389811924805e-08
+    9.460607551398305e-08
+    4.037488423615589e-07
+    2.706690855027815e-08
+    4.791673402232077e-08
+    1.522926538703445e-07
+    4.070682683523807e-07
+ 9.8e+09     
+    4.072512748523676e-07
+    1.519163916801641e-07
+    4.043313225719483e-07
+      4.7901761361156e-08
+    9.466649568735348e-08
+    4.038048223236783e-07
+    2.712123076154362e-08
+    4.797434263858312e-08
+    1.523547515078484e-07
+    4.071245857789493e-07
+ 9.9e+09     
+    4.073082943285951e-07
+    1.519792556092254e-07
+    4.043876125437022e-07
+    4.796017899875798e-08
+    9.472745874480501e-08
+    4.038613507948299e-07
+    2.717613208158424e-08
+    4.803250354034752e-08
+    1.524174565959267e-07
+    4.071814294033397e-07
+ 1e+10       
+    4.073658219931997e-07
+     1.52042735305925e-07
+    4.044444265971605e-07
+    4.801914948944354e-08
+    9.478895949518508e-08
+     4.03918416532984e-07
+    2.723161580222911e-08
+    4.809121539058081e-08
+    1.524807713386255e-07
+    4.072387855312354e-07
+ 1.01e+10    
+    4.074291518940316e-07
+    1.521093693555264e-07
+    4.045066328904309e-07
+    4.808043371133499e-08
+    9.485439787315414e-08
+    4.039806693815412e-07
+    2.728878695400085e-08
+    4.815228227855506e-08
+     1.52547377810851e-07
+    4.073020165720528e-07
+ 1.02e+10    
+    4.074926954905424e-07
+    1.521761034243912e-07
+    4.045689387804566e-07
+    4.814174348781137e-08
+    9.491982463860424e-08
+    4.040430279264992e-07
+     2.73459525230823e-08
+    4.821337436912494e-08
+    1.526140833057561e-07
+    4.073654610943146e-07
+ 1.03e+10    
+    4.075564490882994e-07
+    1.522429324583086e-07
+    4.046313407029074e-07
+    4.820307225915832e-08
+    9.498523511922253e-08
+    4.041054884697791e-07
+    2.740310560309693e-08
+     4.82744851260369e-08
+    1.526808827688975e-07
+    4.074291154329677e-07
+ 1.04e+10    
+    4.076204091131647e-07
+    1.523098515772779e-07
+    4.046938352295498e-07
+    4.826441364171484e-08
+    9.505062484558628e-08
+    4.041680474488048e-07
+    2.746023944509962e-08
+    4.833560818835864e-08
+    1.527477713203002e-07
+    4.074929760432182e-07
+ 1.05e+10    
+    4.076845721080951e-07
+     1.52376856071769e-07
+    4.047564190638383e-07
+    4.832576142535423e-08
+    9.511598954564429e-08
+    4.042307014322394e-07
+    2.751734745546999e-08
+    4.839673736796687e-08
+     1.52814744250701e-07
+    4.075570394973355e-07
+ 1.06e+10    
+    4.077489347299521e-07
+    1.524439413989866e-07
+    4.048190890366213e-07
+    4.838710957091927e-08
+     9.51813251392593e-08
+    4.042934471158178e-07
+    2.757442319377544e-08
+    4.845786664698999e-08
+    1.528817970177964e-07
+    4.076213024814678e-07
+ 1.07e+10    
+    4.078134937463301e-07
+    1.525111031791418e-07
+    4.048818421019482e-07
+    4.844845220761711e-08
+    9.524662773281535e-08
+    4.043562813182768e-07
+    2.763146037060829e-08
+    4.851899017521092e-08
+       1.529489252425e-07
+    4.076857617924767e-07
+ 1.08e+10    
+    4.078782460323978e-07
+    1.525783371917382e-07
+     4.04944675332988e-07
+    4.850978363037862e-08
+     9.53118936138957e-08
+    4.044192009773936e-07
+     2.76884528454006e-08
+    4.858010226743547e-08
+    1.530161247052143e-07
+    4.077504143347906e-07
+ 1.09e+10    
+    4.079431885677712e-07
+    1.526456393718765e-07
+    4.050075859180622e-07
+    4.857109829718793e-08
+    9.537711924603495e-08
+    4.044822031461222e-07
+    2.774539462422083e-08
+    4.864119740083069e-08
+    1.530833913421196e-07
+    4.078152571172808e-07
+ 1.1e+10     
+    4.080083184334058e-07
+    1.527130058065807e-07
+    4.050705711567826e-07
+    4.863239082638559e-08
+    9.544230126354888e-08
+    4.045452849888373e-07
+    2.780227985755561e-08
+    4.870227021223784e-08
+    1.531507212414879e-07
+    4.078802872501661e-07
+ 1.11e+10    
+     4.08073632808524e-07
+    1.527804327311517e-07
+    4.051336284563069e-07
+    4.869365599395076e-08
+    9.550743646644581e-08
+    4.046084437776854e-07
+    2.785910283808004e-08
+    4.876331549546458e-08
+    1.532181106400232e-07
+    4.079455019419494e-07
+ 1.12e+10    
+    4.081391289675748e-07
+    1.528479165255515e-07
+    4.051967553277059e-07
+    4.875488873076638e-08
+    9.557252181542271e-08
+    4.046716768890432e-07
+    2.791585799841973e-08
+     4.88243281985607e-08
+    1.532855559192329e-07
+    4.080108984963867e-07
+ 1.13e+10    
+    4.082048042772292e-07
+    1.529154537108202e-07
+    4.052599493824416e-07
+    4.881608411987092e-08
+     9.56375544269474e-08
+    4.047349818000816e-07
+    2.797253990890729e-08
+    4.888530342108059e-08
+     1.53353053601834e-07
+    4.080764743094929e-07
+ 1.14e+10    
+    4.082706561934165e-07
+    1.529830409455311e-07
+    4.053232083289571e-07
+    4.887723739370115e-08
+    9.570253156843013e-08
+    4.047983560854389e-07
+    2.802914327533645e-08
+    4.894623641133719e-08
+    1.534206003481963e-07
+    4.081422268665897e-07
+ 1.15e+10    
+    4.083366822584017e-07
+    1.530506750222856e-07
+    4.053865299693842e-07
+    4.893834393132911e-08
+    9.576745065348664e-08
+    4.048617974140023e-07
+    2.808566293671587e-08
+    4.900712256365029e-08
+    1.534881929528269e-07
+    4.082081537393912e-07
+ 1.16e+10    
+    4.084028800979069e-07
+    1.531183528642501e-07
+    4.054499121963529e-07
+    4.899939925569685e-08
+    9.583230923729308e-08
+    4.049253035457942e-07
+    2.814209386302562e-08
+    4.906795741559279e-08
+    1.535558283408971e-07
+    4.082742525831383e-07
+ 1.17e+10    
+    4.084692474182818e-07
+    1.531860715217379e-07
+    4.055133529899184e-07
+    4.906039903085159e-08
+    9.589710501203511e-08
+    4.049888723289657e-07
+    2.819843115297806e-08
+    4.912873664523805e-08
+     1.53623503564816e-07
+    4.083405211337782e-07
+ 1.18e+10    
+    4.085357820037193e-07
+    1.532538281688396e-07
+    4.055768504145924e-07
+    4.912133905918602e-08
+    9.596183580245231e-08
+    4.050525016968979e-07
+    2.825467003178575e-08
+    4.918945606841155e-08
+    1.536912158008511e-07
+    4.084069572051902e-07
+ 1.19e+10    
+    4.086024817135251e-07
+    1.533216201001007e-07
+    4.056404026164835e-07
+    4.918221527868401e-08
+    9.602649956147772e-08
+    4.051161896654037e-07
+    2.831080584893791e-08
+    4.925011163594933e-08
+    1.537589623457988e-07
+    4.084735586864667e-07
+ 1.2e+10     
+    4.086693444794405e-07
+     1.53389444727252e-07
+    4.057040078205445e-07
+    4.924302376017685e-08
+    9.609109436597401e-08
+    4.051799343300353e-07
+    2.836683407598759e-08
+    4.931069943096594e-08
+    1.538267406137065e-07
+    4.085403235392416e-07
+ 1.21e+10    
+     4.08736368303014e-07
+    1.534572995759907e-07
+    4.057676643279192e-07
+    4.930376070461121e-08
+    9.615561841256641e-08
+    4.052437338634943e-07
+    2.842275030435103e-08
+    4.937121566613493e-08
+    1.538945481326487e-07
+    4.086072497950771e-07
+ 1.22e+10    
+    4.088035512530363e-07
+    1.535251822828169e-07
+     4.05831370513396e-07
+    4.936442244033099e-08
+    9.622007001357164e-08
+    4.053075865131361e-07
+     2.84785502431208e-08
+    4.943165668098307e-08
+    1.539623825415555e-07
+    4.086743355529019e-07
+ 1.23e+10    
+    4.088708914630275e-07
+    1.535930905919243e-07
+    4.058951248229599e-07
+    4.942500542037689e-08
+    9.628444759302461e-08
+    4.053714905985798e-07
+    2.853422971689446e-08
+    4.949201893920203e-08
+    1.540302415870987e-07
+    4.087415789765071e-07
+ 1.24e+10    
+     4.08938387128784e-07
+    1.536610223521467e-07
+    4.059589257714398e-07
+    4.948550621980355e-08
+    9.634874968280055e-08
+      4.0543544450941e-07
+    2.858978466361952e-08
+    4.955229902597774e-08
+    1.540981231206334e-07
+    4.088089782921016e-07
+ 1.25e+10    
+    4.090060365059859e-07
+    1.537289755139626e-07
+    4.060227719402558e-07
+    4.954592153301787e-08
+    9.641297491883384e-08
+     4.05499446702973e-07
+    2.864521113245659e-08
+    4.961249364534138e-08
+     1.54166025095198e-07
+    4.088765317859252e-07
+ 1.26e+10    
+    4.090738379078647e-07
+     1.53796948126556e-07
+    4.060866619752566e-07
+    4.960624817113939e-08
+    9.647712203743195e-08
+    4.055634957022654e-07
+    2.870050528166118e-08
+    4.967259961754173e-08
+    1.542339455625712e-07
+    4.089442378019211e-07
+ 1.27e+10    
+    4.091417897029345e-07
+    1.538649383349364e-07
+    4.061505945846477e-07
+    4.966648305938507e-08
+    9.654118987168416e-08
+    4.056275900939129e-07
+     2.87556633764858e-08
+    4.973261387644197e-08
+    1.543018826703885e-07
+    4.090120947394694e-07
+ 1.28e+10    
+    4.092098903127806e-07
+    1.539329443771172e-07
+    4.062145685370098e-07
+    4.972662323447919e-08
+    9.660517734796455e-08
+    4.056917285262356e-07
+    2.881068178710277e-08
+    4.979253346694192e-08
+     1.54369834659318e-07
+    4.090801010511829e-07
+ 1.29e+10    
+      4.0927813820992e-07
+    1.540009645813531e-07
+    4.062785826594017e-07
+    4.978666584209059e-08
+    9.666908348252779e-08
+    4.057559097073988e-07
+    2.886555698654896e-08
+    4.985235554242681e-08
+    1.544377998602952e-07
+     4.09148255240766e-07
+ 1.3e+10     
+    4.093465319157182e-07
+    1.540689973634365e-07
+    4.063426358355454e-07
+    4.984660813429783e-08
+    9.673290737819687e-08
+    4.058201324036449e-07
+    2.892028554869311e-08
+    4.991207736224447e-08
+    1.545057766918176e-07
+    4.092165558609328e-07
+ 1.31e+10    
+    4.094150699983769e-07
+    1.541370412240535e-07
+     4.06406727004095e-07
+    4.990644746708391e-08
+    9.679664822114193e-08
+    4.058843954376069e-07
+    2.897486414622629e-08
+     4.99716962892118e-08
+    1.545737636572989e-07
+    4.092850015113951e-07
+ 1.32e+10    
+    4.094837510709808e-07
+    1.542050947461989e-07
+    4.064708551569779e-07
+    4.996618129786164e-08
+    9.686030527774838e-08
+    4.059486976866972e-07
+    2.902928954867632e-08
+    5.003120978715128e-08
+    1.546417593424838e-07
+    4.093535908369075e-07
+ 1.33e+10    
+    4.095525737896169e-07
+    1.542731565926509e-07
+    4.065350193378175e-07
+    5.002580718303024e-08
+    9.692387789157397e-08
+    4.060130380815724e-07
+    2.908355862044658e-08
+    5.009061541845899e-08
+    1.547097624129201e-07
+    4.094223225253816e-07
+ 1.34e+10    
+    4.096215368515563e-07
+    1.543412255035038e-07
+    4.065992186404229e-07
+    5.008532277556438e-08
+    9.698736548039191e-08
+     4.06077415604668e-07
+     2.91376683188798e-08
+    5.014991084170494e-08
+     1.54777771611493e-07
+    4.094911953060631e-07
+ 1.35e+10    
+    4.096906389935005e-07
+    1.544093002937605e-07
+    4.066634522073504e-07
+    5.014472582263645e-08
+    9.705076753332056e-08
+    4.061418292888037e-07
+    2.919161569234711e-08
+    5.020909380926599e-08
+    1.548457857560163e-07
+    4.095602079477748e-07
+ 1.36e+10    
+    4.097598789899012e-07
+    1.544773798509834e-07
+    4.067277192285337e-07
+    5.020401416327264e-08
+    9.711408360803642e-08
+    4.062062782158544e-07
+    2.924539787836286e-08
+    5.026816216499266e-08
+    1.549138037368834e-07
+    4.096293592572231e-07
+ 1.37e+10    
+     4.09829255651339e-07
+    1.545454631330019e-07
+    4.067920189399738e-07
+    5.026318572604343e-08
+    9.717731332807024e-08
+    4.062707615154863e-07
+    2.929901210172538e-08
+    5.032711384191031e-08
+    1.549818245147756e-07
+    4.096986480773722e-07
+ 1.38e+10    
+    4.098987678229736e-07
+    1.546135491656789e-07
+    4.068563506224953e-07
+    5.032223852678896e-08
+    9.724045638018373e-08
+    4.063352783639489e-07
+    2.935245567268415e-08
+    5.038594685995463e-08
+    1.550498471184294e-07
+    4.097680732858808e-07
+ 1.39e+10    
+    4.099684143830613e-07
+    1.546816370407338e-07
+    4.069207136005571e-07
+    5.038117066638036e-08
+    9.730351251182568e-08
+    4.063998279829319e-07
+    2.940572598513338e-08
+    5.044465932374289e-08
+    1.551178706424594e-07
+    4.098376337936052e-07
+ 1.4e+10     
+    4.100381942415367e-07
+    1.547497259136217e-07
+    4.069851072411222e-07
+     5.04399803285163e-08
+    9.736648152866616e-08
+    4.064644096384716e-07
+    2.945882051483235e-08
+    5.050324942038056e-08
+    1.551858942452392e-07
+    4.099073285431708e-07
+ 1.41e+10    
+    4.101081063386629e-07
+    1.548178150014681e-07
+    4.070495309525788e-07
+    5.049866577755605e-08
+     9.74293632922062e-08
+    4.065290226399138e-07
+    2.951173681765254e-08
+    5.056171541730382e-08
+    1.552539171468372e-07
+    4.099771565076029e-07
+ 1.42e+10    
+    4.101781496437477e-07
+    1.548859035810596e-07
+    4.071139841837145e-07
+    5.055722535638927e-08
+    9.749215771746304e-08
+    4.065936663389239e-07
+    2.956447252785161e-08
+    5.062005566015855e-08
+    1.553219386270079e-07
+    4.100471166890261e-07
+ 1.43e+10    
+    4.102483231539267e-07
+    1.549539909868877e-07
+    4.071784664227358e-07
+    5.061565748434168e-08
+    9.755486477072666e-08
+    4.066583401285465e-07
+    2.961702535637449e-08
+    5.067826857071556e-08
+    1.553899580232376e-07
+    4.101172081174272e-07
+ 1.44e+10    
+    4.103186258930109e-07
+    1.550220766092474e-07
+    4.072429771963368e-07
+    5.067396065511856e-08
+    9.761748446738872e-08
+    4.067230434423079e-07
+    2.966939308918142e-08
+     5.07363526448224e-08
+    1.554579747288433e-07
+    4.101874298494842e-07
+ 1.45e+10    
+    4.103890569104009e-07
+    1.550901598923872e-07
+    4.073075160688068e-07
+    5.073213343478419e-08
+    9.768001686983988e-08
+    4.067877757533619e-07
+    2.972157358560286e-08
+    5.079430645039178e-08
+    1.555259881911251e-07
+    4.102577809674552e-07
+ 1.46e+10    
+    4.104596152800665e-07
+    1.551582403327121e-07
+    4.073720826411824e-07
+    5.079017445977876e-08
+    9.774246208543553e-08
+    4.068525365736738e-07
+     2.97735647767216e-08
+    5.085212862542701e-08
+    1.555939979095701e-07
+    4.103282605781346e-07
+ 1.47e+10    
+    4.105303000995887e-07
+    1.552263174770375e-07
+    4.074366765504354e-07
+    5.084808243497238e-08
+    9.780482026452707e-08
+    4.069173254532447e-07
+    2.982536466378155e-08
+    5.090981787608369e-08
+     1.55662003434107e-07
+    4.103988678118698e-07
+ 1.48e+10    
+    4.106011104892672e-07
+    1.552943909208925e-07
+     4.07501297468698e-07
+    5.090585613175523e-08
+    9.786709159855767e-08
+    4.069821419793648e-07
+    2.987697131662344e-08
+    5.096737297476838e-08
+    1.557300043634115e-07
+    4.104696018216416e-07
+ 1.49e+10    
+    4.106720455912909e-07
+    1.553624603068735e-07
+    4.075659451025227e-07
+    5.096349438616543e-08
+    9.792927631822052e-08
+    4.070469857759045e-07
+    2.992838287214731e-08
+     5.10247927582738e-08
+    1.557980003432602e-07
+    4.105404617822044e-07
+ 1.5e+10     
+    4.107431045689701e-07
+    1.554305253230454e-07
+    4.076306191921698e-07
+    5.102099609705282e-08
+     9.79913746916784e-08
+    4.071118565026323e-07
+    2.997959753280129e-08
+    5.108207612595041e-08
+    1.558659910649336e-07
+    4.106114468892896e-07
+ 1.51e+10    
+     4.10814286606029e-07
+    1.554985857013908e-07
+    4.076953195109291e-07
+    5.107836022427983e-08
+      9.8053387022842e-08
+    4.071767538545615e-07
+    3.003061356509717e-08
+    5.113922203791432e-08
+    1.559339762636651e-07
+    4.106825563588673e-07
+ 1.52e+10    
+    4.108855909059621e-07
+     1.55566641216305e-07
+    4.077600458644659e-07
+    5.113558578695822e-08
+    9.811531364970671e-08
+    4.072416775613231e-07
+    3.008142929815184e-08
+    5.119622951329127e-08
+    1.560019557171382e-07
+    4.107537894264675e-07
+ 1.53e+10    
+    4.109570166914463e-07
+     1.55634691683137e-07
+    4.078247980901908e-07
+    5.119267186172211e-08
+    9.817715494274422e-08
+    4.073066273865593e-07
+    3.013204312225511e-08
+    5.125309762849652e-08
+    1.560699292440269e-07
+    4.108251453465599e-07
+ 1.54e+10    
+    4.110285632038131e-07
+    1.557027369567748e-07
+    4.078895760566594e-07
+    5.124961758103686e-08
+     9.82389113033506e-08
+    4.073716031273428e-07
+    3.018245348746307e-08
+    5.130982551555048e-08
+    1.561378967025822e-07
+     4.10896623391992e-07
+ 1.55e+10    
+    4.111002297025776e-07
+    1.557707769302742e-07
+    4.079543796629841e-07
+    5.130642213154326e-08
+    9.830058316234482e-08
+    4.074366046136115e-07
+    3.023265890221728e-08
+     5.13664123604292e-08
+    1.562058579892608e-07
+    4.109682228534799e-07
+ 1.56e+10    
+    4.111720154650247e-07
+    1.558388115335301e-07
+    4.080192088382738e-07
+    5.136308475243708e-08
+    9.836217097852062e-08
+    4.075016317076219e-07
+    3.028265793198923e-08
+    5.142285740145049e-08
+    1.562738130373964e-07
+    4.110399430391586e-07
+ 1.57e+10    
+    4.112439197858474e-07
+    1.559068407319898e-07
+    4.080840635410858e-07
+    5.141960473388357e-08
+    9.842367523724758e-08
+    4.075666843034207e-07
+    3.033244919795004e-08
+    5.147915992769443e-08
+    1.563417618159135e-07
+    4.111117832741837e-07
+ 1.58e+10    
+    4.113159419768416e-07
+     1.55974864525406e-07
+    4.081489437588968e-07
+    5.147598141546619e-08
+    9.848509644911991e-08
+    4.076317623263269e-07
+    3.038203137566484e-08
+    5.153531927745817e-08
+    1.564097043280793e-07
+    4.111837429003858e-07
+ 1.59e+10    
+    4.113880813666487e-07
+    1.560428829466297e-07
+    4.082138495075892e-07
+    5.153221418466968e-08
+    9.854643514865335e-08
+    4.076968657324276e-07
+    3.043140319381189e-08
+    5.159133483674479e-08
+    1.564776406102965e-07
+    4.112558212759756e-07
+ 1.6e+10     
+    4.114603373005522e-07
+    1.561108960604419e-07
+    4.082787808309462e-07
+    5.158830247539687e-08
+    9.860769189302616e-08
+    4.077619945080866e-07
+    3.048056343292607e-08
+    5.164720603778568e-08
+    1.565455707309346e-07
+    4.113280177753014e-07
+ 1.61e+10    
+    4.115327091403205e-07
+    1.561789039624224e-07
+    4.083437378001634e-07
+    5.164424576651853e-08
+    9.866886726086521e-08
+    4.078271486694571e-07
+    3.052951092416608e-08
+    5.170293235759622e-08
+    1.566134947891973e-07
+    4.114003317886517e-07
+ 1.62e+10    
+    4.116051962640989e-07
+    1.562469067778556e-07
+    4.084087205133704e-07
+    5.170004358045649e-08
+    9.872996185107449e-08
+    4.078923282620095e-07
+    3.057824454810575e-08
+    5.175851331656397e-08
+    1.566814129140271e-07
+     4.11472762722106e-07
+ 1.63e+10    
+    4.116777980663422e-07
+    1.563149046606712e-07
+    4.084737290951559e-07
+     5.17556954817987e-08
+    9.879097628170441e-08
+    4.079575333600605e-07
+    3.062676323354833e-08
+     5.18139484770693e-08
+    1.567493252630449e-07
+    4.115453099974314e-07
+ 1.64e+10    
+    4.117505139577979e-07
+    1.563828977924196e-07
+    4.085387636961087e-07
+    5.181120107594681e-08
+    9.885191118886172e-08
+    4.080227640663076e-07
+    3.067506595636428e-08
+    5.186923744213796e-08
+    1.568172320215238e-07
+    4.116179730520209e-07
+ 1.65e+10    
+    4.118233433655216e-07
+    1.564508863812811e-07
+    4.086038244923582e-07
+    5.186656000779464e-08
+    9.891276722565775e-08
+    4.080880205113712e-07
+    3.072315173835144e-08
+    5.192437985412477e-08
+    1.568851334013966e-07
+    4.116907513388769e-07
+ 1.66e+10    
+    4.118962857329419e-07
+    1.565188706611078e-07
+    4.086689116851257e-07
+    5.192177196043811e-08
+     9.89735450611946e-08
+    4.081533028533374e-07
+    3.077101964611782e-08
+     5.19793753934284e-08
+    1.569530296402956e-07
+    4.117636443266283e-07
+ 1.67e+10    
+    4.119693405199547e-07
+    1.565868508904958e-07
+     4.08734025500278e-07
+    5.197683665391555e-08
+     9.90342453795868e-08
+    4.082186112773032e-07
+     3.08186687899865e-08
+    5.203422377723662e-08
+     1.57020921000623e-07
+     4.11836651499593e-07
+ 1.68e+10    
+    4.120425072030566e-07
+    1.566548273518904e-07
+    4.087991661878852e-07
+    5.203175384397791e-08
+    9.909486887901899e-08
+    4.082839459949229e-07
+    3.086609832292209e-08
+    5.208892475830142e-08
+    1.570888077686528e-07
+    4.119097723578714e-07
+ 1.69e+10    
+     4.12115785275511e-07
+    1.567228003507181e-07
+    4.088643340217805e-07
+    5.208652332088864e-08
+    9.915541627083643e-08
+    4.083493072439557e-07
+    3.091330743947877e-08
+    5.214347812374345e-08
+    1.571566902536617e-07
+    4.119830064174757e-07
+ 1.7e+10     
+     4.12189174247546e-07
+     1.56790770214549e-07
+    4.089295292991229e-07
+    5.214114490825247e-08
+    9.921588827866952e-08
+    4.084146952878117e-07
+    3.096029537476922e-08
+    5.219788369388566e-08
+    1.572245687870884e-07
+    4.120563532104915e-07
+ 1.71e+10    
+     4.12262673646578e-07
+    1.568587372922874e-07
+    4.089947523399643e-07
+    5.219561846187277e-08
+    9.927628563758897e-08
+    4.084801104150986e-07
+     3.10070614034544e-08
+    5.225214132111512e-08
+    1.572924437217203e-07
+    4.121298122852683e-07
+ 1.72e+10    
+    4.123362830174678e-07
+    1.569267019533873e-07
+    4.090600034868094e-07
+    5.224994386863669e-08
+    9.933660909329186e-08
+    4.085455529391641e-07
+    3.105360483875352e-08
+    5.230625088877284e-08
+    1.573603154309081e-07
+    4.122033832066419e-07
+ 1.73e+10    
+    4.124100019227933e-07
+    1.569946645870953e-07
+    4.091252831041849e-07
+    5.230412104542788e-08
+    9.939685940131795e-08
+    4.086110231976389e-07
+    3.109992503147401e-08
+    5.236021231007114e-08
+    1.574281843078041e-07
+    4.122770655561747e-07
+ 1.74e+10    
+    4.124838299431518e-07
+    1.570626256017186e-07
+    4.091905915782037e-07
+    5.235814993806627e-08
+    9.945703732629389e-08
+    4.086765215519746e-07
+    3.114602136906122e-08
+    5.241402552703772e-08
+    1.574960507646278e-07
+    4.123508589324274e-07
+ 1.75e+10    
+    4.125577666774767e-07
+    1.571305854239155e-07
+    4.092559293161275e-07
+    5.241203052027386e-08
+    9.951714364120501e-08
+    4.087420483869802e-07
+    3.119189327466717e-08
+    5.246769050948609e-08
+    1.575639152319531e-07
+    4.124247629512485e-07
+ 1.76e+10    
+    4.126318117433738e-07
+    1.571985444980111e-07
+    4.093212967459296e-07
+    5.246576279266667e-08
+    9.957717912669463e-08
+    4.088076041103544e-07
+     3.12375402062384e-08
+    5.252120725401188e-08
+    1.576317781580206e-07
+    4.124987772460831e-07
+ 1.77e+10    
+    4.127059647774704e-07
+    1.572665032853338e-07
+     4.09386694315858e-07
+      5.2519346781772e-08
+    9.963714457038852e-08
+    4.088731891522145e-07
+    3.128296165562216e-08
+    5.257457578301458e-08
+    1.576996400080715e-07
+    4.125729014682989e-07
+ 1.78e+10    
+    4.127802254357795e-07
+     1.57334462263574e-07
+    4.094521224939938e-07
+    5.257278253907022e-08
+    9.969704076624421e-08
+    4.089388039646212e-07
+    3.132815714769092e-08
+    5.262779614374403e-08
+     1.57767501263702e-07
+     4.12647135287525e-07
+ 1.79e+10    
+    4.128545933940734e-07
+    1.574024219261638e-07
+    4.095175817678084e-07
+    5.262607014006138e-08
+    9.975686851392499e-08
+    4.090044490210992e-07
+    3.137312623948462e-08
+    5.268086840737106e-08
+    1.578353624222402e-07
+    4.127214783920092e-07
+ 1.8e+10     
+    4.129290683482631e-07
+     1.57470382781675e-07
+    4.095830726437194e-07
+    5.267920968335495e-08
+    9.981662861819663e-08
+    4.090701248161533e-07
+    3.141786851937022e-08
+    5.273379266808191e-08
+    1.579032239961411e-07
+    4.127959304889736e-07
+ 1.81e+10    
+    4.130036500147843e-07
+    1.575383453532385e-07
+    4.096485956466434e-07
+    5.273220128978332e-08
+    9.987632188834687e-08
+    4.091358318647811e-07
+    3.146238360621866e-08
+    5.278656904219628e-08
+    1.579710865124018e-07
+    4.128704913049936e-07
+ 1.82e+10    
+    4.130783381309871e-07
+    1.576063101779792e-07
+    4.097141513195454e-07
+    5.278504510153777e-08
+    9.993594913762662e-08
+    4.092015707019819e-07
+    3.150667114859819e-08
+    5.283919766730755e-08
+    1.580389505119944e-07
+    4.129451605863656e-07
+ 1.83e+10    
+    4.131531324555255e-07
+     1.57674277806471e-07
+    4.097797402229892e-07
+    5.283774128132675e-08
+    9.999551118271209e-08
+    4.092673418822587e-07
+    3.155073082398437e-08
+    5.289167870144565e-08
+    1.581068165493169e-07
+    4.130199380994919e-07
+ 1.84e+10    
+    4.132280327687445e-07
+    1.577422488022065e-07
+    4.098453629346784e-07
+    5.289029001155582e-08
+    1.000550088431869e-07
+    4.093331459791201e-07
+     3.15945623379858e-08
+    5.294401232226147e-08
+    1.581746851916598e-07
+    4.130948236312581e-07
+ 1.85e+10    
+    4.133030388730648e-07
+    1.578102237410838e-07
+    4.099110200490056e-07
+    5.294269149352882e-08
+    1.001144429410448e-07
+    4.093989835845738e-07
+    3.163816542358579e-08
+    5.299619872623263e-08
+    1.582425570186908e-07
+    4.131698169894126e-07
+ 1.86e+10    
+    4.133781505933597e-07
+    1.578782032109078e-07
+    4.099767121765866e-07
+    5.299494594666979e-08
+    1.001738143002096e-07
+    4.094648553086203e-07
+    3.168153984039914e-08
+    5.304823812788982e-08
+    1.583104326219523e-07
+    4.132449180029415e-07
+ 1.87e+10    
+    4.134533677773254e-07
+    1.579461878109075e-07
+    4.100424399438031e-07
+    5.304705360776519e-08
+    1.002331237460753e-07
+    4.095307617787415e-07
+    3.172468537394406e-08
+    5.310013075906361e-08
+    1.583783126043758e-07
+    4.133201265224393e-07
+ 1.88e+10    
+    4.135286902958391e-07
+    1.580141781512648e-07
+    4.101082039923363e-07
+    5.309901473022556e-08
+    1.002923721050625e-07
+    4.095967036393833e-07
+    3.176760183492859e-08
+    5.315187686815077e-08
+    1.584461975798088e-07
+    4.133954424204696e-07
+ 1.89e+10    
+    4.136041180433072e-07
+    1.580821748526594e-07
+     4.10174004978702e-07
+    5.315082958336699e-08
+    1.003515602041929e-07
+    4.096626815514414e-07
+    3.181028905855151e-08
+    5.320347671940014e-08
+    1.585140881725573e-07
+    4.134708655919205e-07
+ 1.9e+10     
+    4.136796509379951e-07
+    1.581501785458238e-07
+    4.102398435737826e-07
+    5.320249845171075e-08
+    1.004106888706789e-07
+    4.097286961917369e-07
+    3.185274690381702e-08
+    5.325493059221723e-08
+    1.585819850169371e-07
+    4.135463959543419e-07
+ 1.91e+10    
+    4.137552889223444e-07
+    1.582181898711121e-07
+    4.103057204623576e-07
+     5.32540216343019e-08
+    1.004697589315313e-07
+     4.09794748252495e-07
+    3.189497525286327e-08
+    5.330623878048702e-08
+    1.586498887568419e-07
+    4.136220334482761e-07
+ 1.92e+10    
+    4.138310319632699e-07
+    1.582862094780786e-07
+    4.103716363426318e-07
+     5.33053994440451e-08
+      1.0052877121318e-07
+    4.098608384408185e-07
+    3.193697401030406e-08
+     5.33574015919149e-08
+    1.587178000453195e-07
+    4.136977780375679e-07
+ 1.93e+10    
+    4.139068800524391e-07
+    1.583542380250696e-07
+    4.104375919257663e-07
+    5.335663220705879e-08
+     1.00587726541112e-07
+    4.099269674781622e-07
+     3.19787431025838e-08
+    5.340841934738513e-08
+    1.587857195441612e-07
+    4.137736297096607e-07
+ 1.94e+10    
+    4.139828332065264e-07
+    1.584222761788227e-07
+    4.105035879354021e-07
+    5.340772026204527e-08
+     1.00646625739522e-07
+    4.099931360998022e-07
+    3.202028247734498e-08
+    5.345929238033591e-08
+       1.588536479235e-07
+    4.138495884758717e-07
+ 1.95e+10    
+    4.140588914674462e-07
+    1.584903246140779e-07
+    4.105696251071884e-07
+    5.345866395967835e-08
+    1.007054696309779e-07
+    4.100593450543087e-07
+    3.206159210280816e-08
+    5.351002103615155e-08
+    1.589215858614207e-07
+    4.139256543716499e-07
+ 1.96e+10    
+    4.141350549025655e-07
+    1.585583840131975e-07
+    4.106357041883098e-07
+    5.350946366200661e-08
+    1.007642590360997e-07
+    4.101255951030139e-07
+    3.210267196716417e-08
+    5.356060567157058e-08
+    1.589895340435772e-07
+    4.140018274568074e-07
+ 1.97e+10    
+    4.142113236048822e-07
+    1.586264550657942e-07
+    4.107018259370112e-07
+     5.35601197418726e-08
+    1.008229947732511e-07
+    4.101918870194831e-07
+    3.214352207797804e-08
+    5.361104665410948e-08
+    1.590574931628212e-07
+    4.140781078157316e-07
+ 1.98e+10    
+    4.142876976931857e-07
+    1.586945384683683e-07
+    4.107679911221252e-07
+    5.361063258234727e-08
+    1.008816776582444e-07
+    4.102582215889849e-07
+    3.218414246160459e-08
+    5.366134436150214e-08
+    1.591254639188377e-07
+     4.14154495557573e-07
+ 1.99e+10    
+    4.143641773121821e-07
+    1.587626349239526e-07
+    4.108342005225991e-07
+    5.366100257617963e-08
+    1.009403085040572e-07
+      4.1032459960796e-07
+    3.222453316261528e-08
+    5.371149918115386e-08
+     1.59193447017789e-07
+    4.142309908164023e-07
+ 2e+10       
+    4.144407626325954e-07
+    1.588307451417648e-07
+     4.10900454927026e-07
+    5.371123012526064e-08
+    1.009988881205609e-07
+    4.103910218834954e-07
+    3.226469424323622e-08
+    5.376151150961047e-08
+    1.592614431719675e-07
+    4.143075937513472e-07
+ 2.01e+10    
+    4.145174538512357e-07
+    1.588988698368665e-07
+    4.109667551331693e-07
+    5.376131564010183e-08
+    1.010574173142609e-07
+    4.104574892327971e-07
+    3.230462578279681e-08
+    5.381138175204097e-08
+     1.59329453099454e-07
+    4.143843045466966e-07
+ 2.02e+10    
+    4.145942511910376e-07
+      1.5896700972983e-07
+    4.110331019475003e-07
+    5.381125953932704e-08
+    1.011158968880481e-07
+     4.10524002482666e-07
+    3.234432787718904e-08
+    5.386111032173464e-08
+    1.593974775237849e-07
+    4.144611234119795e-07
+ 2.03e+10    
+    4.146711549010699e-07
+    1.590351655464106e-07
+    4.110994961847262e-07
+    5.386106224917848e-08
+    1.011743276409607e-07
+    4.105905624689742e-07
+    3.238380063833707e-08
+    5.391069763961125e-08
+    1.594655171736242e-07
+    4.145380505820102e-07
+ 2.04e+10    
+    4.147481652565086e-07
+    1.591033380172263e-07
+    4.111659386673323e-07
+    5.391072420303536e-08
+    1.012327103679566e-07
+    4.106571700361477e-07
+    3.242304419367688e-08
+    5.396014413374472e-08
+    1.595335727824434e-07
+     4.14615086316909e-07
+ 2.05e+10    
+    4.148252825585812e-07
+    1.591715278774404e-07
+    4.112324302251156e-07
+    5.396024584094556e-08
+    1.012910458596965e-07
+    4.107238260366505e-07
+    3.246205868564576e-08
+    5.400945023889908e-08
+    1.596016450882059e-07
+    4.146922309020868e-07
+ 2.06e+10    
+    4.149025071344792e-07
+    1.592397358664539e-07
+    4.112989716947284e-07
+    5.400962760917001e-08
+    1.013493349023355e-07
+    4.107905313304711e-07
+     3.25008442711815e-08
+    5.405861639607751e-08
+    1.596697348330587e-07
+    4.147694846482029e-07
+ 2.07e+10    
+    4.149798393372348e-07
+    1.593079627275994e-07
+    4.113655639192254e-07
+    5.405886995973877e-08
+    1.014075782773259e-07
+    4.108572867846163e-07
+    3.253940112123093e-08
+    5.410764305208316e-08
+    1.597378427630281e-07
+     4.14846847891089e-07
+ 2.08e+10    
+     4.15057279545567e-07
+     1.59376209207842e-07
+    4.114322077476097e-07
+    5.410797335001972e-08
+    1.014657767612275e-07
+     4.10924093272607e-07
+    3.257772942026774e-08
+    5.415653065909184e-08
+    1.598059696277211e-07
+    4.149243209916419e-07
+ 2.09e+10    
+    4.151348281636961e-07
+    1.594444760574841e-07
+     4.11498904034388e-07
+     5.41569382422979e-08
+    1.015239311255279e-07
+    4.109909516739783e-07
+    3.261582936581934e-08
+    5.420527967423639e-08
+    1.598741161800323e-07
+    4.150019043356864e-07
+ 2.1e+10     
+    4.152124856211237e-07
+    1.595127640298763e-07
+    4.115656536391291e-07
+    5.420576510336742e-08
+    1.015820421364714e-07
+    4.110578628737897e-07
+    3.265370116800256e-08
+    5.425389055920223e-08
+    1.599422831758547e-07
+    4.150795983338037e-07
+ 2.11e+10    
+    4.152902523723816e-07
+    1.595810738811305e-07
+    4.116324574260235e-07
+    5.425445440413307e-08
+    1.016401105548959e-07
+    4.111248277621346e-07
+    3.269134504906804e-08
+    5.430236377983389e-08
+    1.600104713737957e-07
+    4.151574034211306e-07
+ 2.12e+10    
+    4.153681288967489e-07
+    1.596494063698389e-07
+    4.116993162634517e-07
+    5.430300661922378e-08
+    1.016981371360778e-07
+     4.11191847233661e-07
+    3.272876124295312e-08
+    5.435069980575222e-08
+    1.600786815348972e-07
+    4.152353200571272e-07
+ 2.13e+10    
+    4.154461156979372e-07
+    1.597177622567968e-07
+    4.117662310235587e-07
+    5.435142222661595e-08
+    1.017561226295855e-07
+    4.112589221870948e-07
+    3.276594999484307e-08
+    5.439889910998211e-08
+    1.601469144223599e-07
+    4.153133487253122e-07
+ 2.14e+10    
+    4.155242133037505e-07
+    1.597861423047296e-07
+    4.118332025818296e-07
+    5.439970170726756e-08
+    1.018140677791398e-07
+    4.113260535247726e-07
+    3.280291156074068e-08
+    5.444696216859045e-08
+     1.60215170801272e-07
+    4.153914899329696e-07
+ 2.15e+10    
+    4.156024222657033e-07
+    1.598545472780225e-07
+    4.119002318166748e-07
+    5.444784554476173e-08
+    1.018719733224822e-07
+    4.113932421521807e-07
+    3.283964620704355e-08
+     5.44948894603338e-08
+    1.602834514383416e-07
+     4.15469744210825e-07
+ 2.16e+10    
+    4.156807431586243e-07
+     1.59922977942456e-07
+    4.119673196090205e-07
+    5.449585422496064e-08
+    1.019298399912501e-07
+    4.114604889774993e-07
+    3.287615421012966e-08
+    5.454268146631601e-08
+    1.603517571016331e-07
+    4.155481121126917e-07
+ 2.17e+10    
+    4.157591765802209e-07
+    1.599914350649434e-07
+    4.120344668419044e-07
+    5.454372823566871e-08
+    1.019876685108595e-07
+    4.115277949111596e-07
+    3.291243585595048e-08
+    5.459033866965519e-08
+    1.604200885603072e-07
+    4.156265942150884e-07
+ 2.18e+10    
+    4.158377231506213e-07
+    1.600599194132729e-07
+    4.121016744000796e-07
+    5.459146806630531e-08
+    1.020454596003935e-07
+    4.115951608654014e-07
+    3.294849143963185e-08
+    5.463786155516001e-08
+    1.604884465843652e-07
+    4.157051911168316e-07
+ 2.19e+10    
+    4.159163835118892e-07
+    1.601284317558529e-07
+    4.121689431696235e-07
+     5.46390742075864e-08
+    1.021032139724982e-07
+    4.116625877538448e-07
+    3.298432126508236e-08
+    5.468525060901506e-08
+     1.60556831944396e-07
+    4.157839034385971e-07
+ 2.2e+10     
+     4.15995158327514e-07
+     1.60196972861461e-07
+    4.122362740375554e-07
+    5.468654715121552e-08
+    1.021609323332847e-07
+    4.117300764910694e-07
+    3.301992564460905e-08
+    5.473250631847486e-08
+    1.606252454113278e-07
+    4.158627318224591e-07
+ 2.21e+10    
+    4.160740482818764e-07
+    1.602655434989973e-07
+    4.123036678914613e-07
+     5.47338873895831e-08
+    1.022186153822377e-07
+    4.117976279921981e-07
+    3.305530489854059e-08
+    5.477962917156681e-08
+    1.606936877561822e-07
+    4.159416769314027e-07
+ 2.22e+10    
+    4.161530540796911e-07
+    1.603341444372392e-07
+    4.123711256191236e-07
+    5.478109541547468e-08
+    1.022762638121287e-07
+    4.118652431724941e-07
+    3.309045935485762e-08
+    5.482661965680244e-08
+    1.607621597498331e-07
+    4.160207394488129e-07
+ 2.23e+10    
+    4.162321764454299e-07
+     1.60402776444602e-07
+    4.124386481081611e-07
+     5.48281717217874e-08
+    1.023338783089369e-07
+     4.11932922946964e-07
+    3.312538934882993e-08
+    5.487347826289673e-08
+     1.60830662162767e-07
+    4.160999200779395e-07
+ 2.24e+10    
+    4.163114161227201e-07
+    1.604714402889022e-07
+    4.125062362456763e-07
+    5.487511680125469e-08
+    1.023914595517742e-07
+    4.120006682299735e-07
+    3.316009522266117e-08
+      5.4920205478496e-08
+    1.608991957648508e-07
+    4.161792195413451e-07
+ 2.25e+10    
+    4.163907738737297e-07
+    1.605401367371233e-07
+    4.125738909179103e-07
+      5.4921931146179e-08
+    1.024490082128169e-07
+    4.120684799348661e-07
+     3.31945773251399e-08
+    5.496680179191332e-08
+    1.609677613250975e-07
+    4.162586385803273e-07
+ 2.26e+10    
+     4.16470250478531e-07
+    1.606088665551869e-07
+    4.126416130099019e-07
+    5.496861524817261e-08
+    1.025065249572413e-07
+    4.121363589735988e-07
+    3.322883601129796e-08
+     5.50132676908717e-08
+    1.610363596114407e-07
+     4.16338177954325e-07
+ 2.27e+10    
+    4.165498467344509e-07
+    1.606776305077263e-07
+    4.127094034051641e-07
+    5.501516959790599e-08
+    1.025640104431658e-07
+    4.122043062563808e-07
+    3.326287164207532e-08
+    5.505960366225523e-08
+    1.611049913905092e-07
+    4.164178384403076e-07
+ 2.28e+10    
+     4.16629563455403e-07
+    1.607464293578634e-07
+    4.127772629853574e-07
+    5.506159468486355e-08
+    1.026214653215968e-07
+    4.122723226913259e-07
+    3.329668458399155e-08
+    5.510581019186705e-08
+    1.611736574274067e-07
+    4.164976208321431e-07
+ 2.29e+10    
+    4.167094014712117e-07
+    1.608152638669912e-07
+    4.128451926299806e-07
+    5.510789099710755e-08
+    1.026788902363809e-07
+    4.123404091841125e-07
+    3.333027520882434e-08
+    5.515188776419533e-08
+    1.612423584854946e-07
+    4.165775259399613e-07
+ 2.3e+10     
+    4.167893616269171e-07
+    1.608841347945562e-07
+    4.129131932160635e-07
+    5.515405902104819e-08
+    1.027362858241595e-07
+     4.12408566637653e-07
+    3.336364389329387e-08
+    5.519783686218568e-08
+    1.613110953261781e-07
+    4.166575545894907e-07
+ 2.31e+10    
+    4.168694447820797e-07
+      1.6095304289785e-07
+    4.129812656178743e-07
+    5.520009924122208e-08
+    1.027936527143306e-07
+    4.124767959517763e-07
+    3.339679101875431e-08
+    5.524365796702135e-08
+     1.61379868708697e-07
+    4.167377076213939e-07
+ 2.32e+10    
+    4.169496518100661e-07
+    1.610219889317986e-07
+    4.130494107066276e-07
+     5.52460121400767e-08
+    1.028509915290126e-07
+    4.125450980229136e-07
+    3.342971697089128e-08
+    5.528935155790932e-08
+    1.614486793899188e-07
+    4.168179858905866e-07
+ 2.33e+10    
+    4.170299835973339e-07
+    1.610909736487604e-07
+    4.131176293502081e-07
+    5.529179819776238e-08
+    1.029083028830143e-07
+    4.126134737438038e-07
+    3.346242213942582e-08
+    5.533491811187425e-08
+    1.615175281241367e-07
+    4.168983902655488e-07
+ 2.34e+10    
+    4.171104410427063e-07
+    1.611599977983249e-07
+    4.131859224128991e-07
+    5.533745789193064e-08
+    1.029655873838071e-07
+    4.126819240031964e-07
+    3.349490691782459e-08
+    5.538035810355803e-08
+    1.615864156628705e-07
+    4.169789216276283e-07
+ 2.35e+10    
+    4.171910250566482e-07
+    1.612290621271176e-07
+    4.132542907551196e-07
+    5.538299169753959e-08
+    1.030228456315029e-07
+    4.127504496855755e-07
+    3.352717170301637e-08
+    5.542567200502648e-08
+    1.616553427546717e-07
+    4.170595808703369e-07
+ 2.36e+10    
+    4.172717365605319e-07
+    1.612981673786073e-07
+    4.133227352331726e-07
+    5.542840008666531e-08
+    1.030800782188348e-07
+    4.128190516708865e-07
+    3.355921689511462e-08
+    5.547086028558222e-08
+    1.617243101449322e-07
+    4.171403688986417e-07
+ 2.37e+10    
+    4.173525764859046e-07
+    1.613673142929179e-07
+    4.133912566989975e-07
+    5.547368352832026e-08
+    1.031372857311418e-07
+    4.128877308342763e-07
+    3.359104289714625e-08
+    5.551592341158375e-08
+    1.617933185756981e-07
+    4.172212866282563e-07
+ 2.38e+10    
+    4.174335457737572e-07
+     1.61436503606644e-07
+    4.134598559999344e-07
+    5.551884248827729e-08
+    1.031944687463571e-07
+    4.129564880458402e-07
+    3.362265011478622e-08
+    5.556086184627049e-08
+    1.618623687854851e-07
+    4.173023349849197e-07
+ 2.39e+10    
+    4.175146453737904e-07
+    1.615057360526718e-07
+    4.135285339784966e-07
+    5.556387742890031e-08
+    1.032516278349998e-07
+    4.130253241703812e-07
+    3.365403895609846e-08
+    5.560567604959439e-08
+       1.619314615091e-07
+     4.17383514903686e-07
+ 2.4e+10     
+    4.175958762436852e-07
+    1.615750123600022e-07
+    4.135972914721498e-07
+    5.560878880898082e-08
+      1.0330876356017e-07
+    4.130942400671767e-07
+    3.368520983128248e-08
+    5.565036647805691e-08
+    1.620005974774654e-07
+    4.174648273282064e-07
+ 2.41e+10    
+     4.17677239348374e-07
+    1.616443332535799e-07
+    4.136661293131011e-07
+    5.565357708358037e-08
+    1.033658764775473e-07
+    4.131632365897572e-07
+    3.371616315242597e-08
+    5.569493358455201e-08
+    1.620697774174486e-07
+    4.175462732100163e-07
+ 2.42e+10    
+    4.177587356593226e-07
+    1.617136994541253e-07
+    4.137350483280952e-07
+    5.569824270387898e-08
+    1.034229671353918e-07
+    4.132323145856906e-07
+     3.37468993332632e-08
+    5.573937781821493e-08
+    1.621390020516943e-07
+    4.176278535078221e-07
+ 2.43e+10    
+    4.178403661538089e-07
+    1.617831116779721e-07
+    4.138040493382212e-07
+    5.574278611702905e-08
+    1.034800360745492e-07
+    4.133014748963801e-07
+    3.377741878893922e-08
+    5.578369962427637e-08
+    1.622082720984619e-07
+    4.177095691867946e-07
+ 2.44e+10    
+    4.179221318142155e-07
+    1.618525706369078e-07
+    4.138731331587241e-07
+     5.57872077660152e-08
+    1.035370838284575e-07
+    4.133707183568691e-07
+    3.380772193577984e-08
+    5.582789944392246e-08
+    1.622775882714671e-07
+    4.177914212178658e-07
+ 2.45e+10    
+    4.180040336273279e-07
+    1.619220770380196e-07
+    4.139423005988266e-07
+    5.583150808951935e-08
+    1.035941109231576e-07
+    4.134400457956536e-07
+    3.383780919106718e-08
+    5.587197771415988e-08
+    1.623469512797269e-07
+    4.178734105770328e-07
+ 2.46e+10    
+    4.180860725836414e-07
+    1.619916315835438e-07
+    4.140115524615583e-07
+    5.587568752179145e-08
+    1.036511178773059e-07
+     4.13509458034507e-07
+    3.386768097282094e-08
+    5.591593486768622e-08
+    1.624163618274101e-07
+    4.179555382446671e-07
+ 2.47e+10    
+    4.181682496766753e-07
+    1.620612349707207e-07
+    4.140808895435954e-07
+    5.591974649252529e-08
+    1.037081052021897e-07
+    4.135789558883119e-07
+    3.389733769958516e-08
+    5.595977133276597e-08
+    1.624858206136906e-07
+    4.180378052048347e-07
+ 2.48e+10    
+    4.182505659023043e-07
+    1.621308878916527e-07
+    4.141503126351009e-07
+    5.596368542673986e-08
+    1.037650734017454e-07
+    4.136485401649013e-07
+    3.392677979022056e-08
+    5.600348753311104e-08
+    1.625553283326067e-07
+    4.181202124446206e-07
+ 2.49e+10    
+    4.183330222580947e-07
+    1.622005910331671e-07
+    4.142198225195819e-07
+    5.600750474466537e-08
+    1.038220229725785e-07
+    4.137182116649055e-07
+    3.395600766370238e-08
+    5.604708388776679e-08
+    1.626248856729229e-07
+     4.18202760953471e-07
+ 2.5e+10     
+    4.184156197426552e-07
+    1.622703450766847e-07
+     4.14289419973748e-07
+    5.605120486163487e-08
+    1.038789544039862e-07
+    4.137879711816119e-07
+    3.398502173892349e-08
+    5.609056081100283e-08
+    1.626944933179978e-07
+    4.182854517225375e-07
+ 2.51e+10    
+    4.184983593550049e-07
+    1.623401506980905e-07
+     4.14359105767379e-07
+    5.609478618798021e-08
+    1.039358681779826e-07
+    4.138578195008319e-07
+    3.401382243450301e-08
+    5.613391871220835e-08
+     1.62764151945655e-07
+     4.18368285744039e-07
+ 2.52e+10    
+    4.185812420939463e-07
+    1.624100085676108e-07
+    4.144288806632006e-07
+    5.613824912893322e-08
+    1.039927647693254e-07
+    4.139277574007716e-07
+    3.404241016860006e-08
+    5.617715799579283e-08
+    1.628338622280591e-07
+    4.184512640106346e-07
+ 2.53e+10    
+    4.186642689574619e-07
+    1.624799193496937e-07
+    4.144987454167654e-07
+    5.618159408453166e-08
+    1.040496446455447e-07
+    4.139977856519166e-07
+    3.407078535873293e-08
+    5.622027906109053e-08
+    1.629036248315955e-07
+    4.185343875148069e-07
+ 2.54e+10    
+    4.187474409421197e-07
+    1.625498837028942e-07
+    4.145687007763449e-07
+    5.622482144952941e-08
+    1.041065082669742e-07
+    4.140679050169206e-07
+    3.409894842160328e-08
+    5.626328230227055e-08
+    1.629734404167553e-07
+    4.186176572482633e-07
+ 2.55e+10    
+    4.188307590424963e-07
+    1.626199022797643e-07
+    4.146387474828234e-07
+    5.626793161331158e-08
+    1.041633560867839e-07
+    4.141381162505032e-07
+    3.412689977292555e-08
+    5.630616810825042e-08
+    1.630433096380238e-07
+    4.187010742013485e-07
+ 2.56e+10    
+    4.189142242506166e-07
+    1.626899757267462e-07
+    4.147088862696016e-07
+    5.631092495981417e-08
+    1.042201885510146e-07
+    4.142084200993544e-07
+     3.41546398272614e-08
+     5.63489368626147e-08
+    1.631132331437739e-07
+    4.187846393624728e-07
+ 2.57e+10    
+    4.189978375554058e-07
+    1.627601046840712e-07
+    4.147791178625077e-07
+    5.635380186744745e-08
+    1.042770060986144e-07
+    4.142788173020467e-07
+    3.418216899785905e-08
+    5.639158894353758e-08
+    1.631832115761628e-07
+    4.188683537175552e-07
+ 2.58e+10    
+    4.190815999421674e-07
+    1.628302897856631e-07
+     4.14849442979713e-07
+     5.63965627090246e-08
+    1.043338091614764e-07
+    4.143493085889552e-07
+    3.420948769649791e-08
+    5.643412472370989e-08
+     1.63253245571035e-07
+    4.189522182494847e-07
+ 2.59e+10    
+    4.191655123920641e-07
+    1.629005316590431e-07
+    4.149198623316533e-07
+     5.64392078516934e-08
+     1.04390598164478e-07
+    4.144198946821819e-07
+     3.42365963333375e-08
+    5.647654457026983e-08
+    1.633233357578269e-07
+    4.190362339375929e-07
+ 2.6e+10     
+    4.192495758816306e-07
+    1.629708309252434e-07
+    4.149903766209601e-07
+    5.648173765687319e-08
+    1.044473735255224e-07
+    4.144905762954902e-07
+    3.426349531677178e-08
+    5.651884884473834e-08
+     1.63393482759478e-07
+    4.191204017571487e-07
+ 2.61e+10    
+    4.193337913822935e-07
+    1.630411881987214e-07
+    4.150609865423937e-07
+    5.652415248019478e-08
+    1.045041356555803e-07
+    4.145613541342438e-07
+    3.429018505328782e-08
+    5.656103790295784e-08
+    1.634636871923453e-07
+    4.192047226788647e-07
+ 2.62e+10    
+    4.194181598599134e-07
+    1.631116040872797e-07
+     4.15131692782786e-07
+    5.656645267144491e-08
+     1.04560884958734e-07
+    4.146322288953522e-07
+    3.431666594732939e-08
+    5.660311209503519e-08
+    1.635339496661209e-07
+    4.192891976684246e-07
+ 2.63e+10    
+    4.195026822743448e-07
+    1.631820791919901e-07
+    4.152024960209839e-07
+    5.660863857451453e-08
+    1.046176218322221e-07
+    4.147032012672232e-07
+      3.4342938401165e-08
+    5.664507176528827e-08
+    1.636042707837558e-07
+    4.193738276860252e-07
+ 2.64e+10    
+    4.195873595790114e-07
+    1.632526141071215e-07
+    4.152733969278066e-07
+    5.665071052735023e-08
+    1.046743466664857e-07
+    4.147742719297198e-07
+    3.436900281476062e-08
+     5.66869172521964e-08
+    1.636746511413863e-07
+    4.194586136859374e-07
+ 2.65e+10    
+    4.196721927204999e-07
+    1.633232094200714e-07
+    4.153443961659986e-07
+     5.66926688619101e-08
+    1.047310598452158e-07
+    4.148454415541261e-07
+    3.439485958565673e-08
+    5.672864888835401e-08
+    1.637450913282644e-07
+    4.195435566160825e-07
+ 2.66e+10    
+    4.197571826381775e-07
+     1.63393865711303e-07
+    4.154154943901961e-07
+    5.673451390412272e-08
+    1.047877617454015e-07
+    4.149167108031149e-07
+    3.442050910885007e-08
+    5.677026700042845e-08
+    1.638155919266934e-07
+    4.196286574176289e-07
+ 2.67e+10    
+    4.198423302638159e-07
+    1.634645835542838e-07
+    4.154866922468928e-07
+     5.67762459738495e-08
+    1.048444527373795e-07
+    4.149880803307239e-07
+    3.444595177667935e-08
+     5.68117719091206e-08
+    1.638861535119657e-07
+    4.197139170246036e-07
+ 2.68e+10    
+    4.199276365212447e-07
+    1.635353635154301e-07
+    4.155579903744156e-07
+    5.681786538485076e-08
+    1.049011331848844e-07
+    4.150595507823352e-07
+    3.447118797871557e-08
+    5.685316392912924e-08
+    1.639567766523058e-07
+    4.197993363635225e-07
+ 2.69e+10    
+    4.200131023260127e-07
+    1.636062061540544e-07
+    4.156293894029006e-07
+    5.685937244475497e-08
+    1.049578034450996e-07
+     4.15131122794661e-07
+    3.449621810165637e-08
+    5.689444336911867e-08
+    1.640274619088167e-07
+    4.198849163530393e-07
+ 2.7e+10     
+    4.200987285850749e-07
+    1.636771120223164e-07
+    4.157008899542766e-07
+    5.690076745503106e-08
+    1.050144638687099e-07
+     4.15202796995735e-07
+    3.452104252922458e-08
+    5.693561053168933e-08
+    1.640982098354297e-07
+    4.199706579036086e-07
+ 2.71e+10    
+    4.201845161964928e-07
+    1.637480816651785e-07
+    4.157724926422546e-07
+    5.694205071096421e-08
+    1.050711147999539e-07
+    4.152745740049058e-07
+    3.454566164207083e-08
+    5.697666571335164e-08
+    1.641690209788582e-07
+    4.200565619171695e-07
+ 2.72e+10    
+    4.202704660491493e-07
+    1.638191156203635e-07
+    4.158441980723167e-07
+    5.698322250163427e-08
+     1.05127756576678e-07
+    4.153464544328387e-07
+    3.457007581768019e-08
+    5.701760920450317e-08
+    1.642398958785553e-07
+    4.201426292868448e-07
+ 2.73e+10    
+    4.203565790224867e-07
+    1.638902144183172e-07
+     4.15916006841713e-07
+     5.70242831098975e-08
+      1.0518438953039e-07
+    4.154184388815186e-07
+    3.459428543028267e-08
+    5.705844128940822e-08
+    1.643108350666744e-07
+    4.202288608966578e-07
+ 2.74e+10    
+    4.204428559862563e-07
+    1.639613785821736e-07
+    4.159879195394634e-07
+    5.706523281237112e-08
+    1.052410139863149e-07
+    4.154905279442592e-07
+    3.461829085076759e-08
+    5.709916224618068e-08
+    1.643818390680332e-07
+    4.203152576212623e-07
+ 2.75e+10    
+    4.205292978002882e-07
+    1.640326086277239e-07
+    4.160599367463591e-07
+    5.710607187942062e-08
+    1.052976302634494e-07
+    4.155627222057146e-07
+    3.464209244660192e-08
+    5.713977234676967e-08
+    1.644529084000821e-07
+    4.204018203256977e-07
+ 2.76e+10    
+    4.206159053142725e-07
+    1.641039050633879e-07
+    4.161320590349735e-07
+    5.714680057514967e-08
+    1.053542386746188e-07
+    4.156350222418987e-07
+    3.466569058175198e-08
+    5.718027185694777e-08
+    1.645240435728744e-07
+    4.204885498651501e-07
+ 2.77e+10    
+    4.207026793675612e-07
+    1.641752683901903e-07
+    4.162042869696728e-07
+    5.718741915739309e-08
+     1.05410839526533e-07
+    4.157074286202024e-07
+    3.468908561660915e-08
+    5.722066103630205e-08
+    1.645952450890414e-07
+    4.205754470847353e-07
+ 2.78e+10    
+    4.207896207889837e-07
+    1.642466991017379e-07
+    4.162766211066301e-07
+    5.722792787771203e-08
+    1.054674331198433e-07
+    4.157799418994195e-07
+    3.471227790791895e-08
+    5.726094013822754e-08
+    1.646665134437687e-07
+    4.206625128192982e-07
+ 2.79e+10    
+    4.208767303966756e-07
+    1.643181976842019e-07
+    4.163490619938456e-07
+    5.726832698139177e-08
+    1.055240197492005e-07
+    4.158525626297742e-07
+    3.473526780871367e-08
+    5.730110940992339e-08
+    1.647378491247775e-07
+    4.207497478932238e-07
+ 2.8e+10     
+    4.209640089979246e-07
+    1.643897646163018e-07
+    4.164216101711688e-07
+    5.730861670744199e-08
+    1.055805997033118e-07
+    4.159252913529514e-07
+    3.475805566824843e-08
+    5.734116909239121e-08
+    1.648092526123074e-07
+    4.208371531202652e-07
+ 2.81e+10    
+    4.210514573890319e-07
+    1.644614003692928e-07
+    4.164942661703223e-07
+    5.734879728859955e-08
+    1.056371732649994e-07
+    4.159981286021323e-07
+    3.478064183194074e-08
+    5.738111942043614e-08
+    1.648807243791032e-07
+    4.209247293033875e-07
+ 2.82e+10    
+    4.211390763551829e-07
+    1.645331054069556e-07
+     4.16567030514931e-07
+    5.738886895133303e-08
+    1.056937407112588e-07
+    4.160710749020285e-07
+     3.48030266413131e-08
+    5.742096062266993e-08
+    1.649522648904036e-07
+    4.210124772346248e-07
+ 2.83e+10    
+    4.212268666703365e-07
+     1.64604880185589e-07
+     4.16639903720553e-07
+    5.742883191585026e-08
+    1.057503023133172e-07
+    4.161441307689265e-07
+    3.482521043393908e-08
+    5.746069292151632e-08
+    1.650238746039334e-07
+    4.211003976949497e-07
+ 2.84e+10    
+    4.213148290971251e-07
+    1.646767251540059e-07
+     4.16712886294713e-07
+    5.746868639610724e-08
+    1.058068583366922e-07
+    4.162172967107269e-07
+    3.484719354339237e-08
+    5.750031653321854e-08
+    1.650955539698978e-07
+    4.211884914541603e-07
+ 2.85e+10    
+    4.214029643867686e-07
+      1.6474864075353e-07
+    4.167859787369389e-07
+    5.750843259981977e-08
+    1.058634090412513e-07
+    4.162905732269915e-07
+    3.486897629919909e-08
+    5.753983166784904e-08
+    1.651673034309796e-07
+    4.212767592707758e-07
+ 2.86e+10    
+    4.214912732790004e-07
+    1.648206274179975e-07
+    4.168591815388026e-07
+    5.754807072847658e-08
+    1.059199546812708e-07
+    4.163639608089911e-07
+    3.489055902679307e-08
+    5.757923852932124e-08
+    1.652391234223387e-07
+    4.213652018919499e-07
+ 2.87e+10    
+    4.215797565020041e-07
+    1.648926855737582e-07
+    4.169324951839578e-07
+    5.758760097735468e-08
+    1.059764955054947e-07
+    4.164374599397557e-07
+    3.491194204747394e-08
+    5.761853731540296e-08
+    1.653110143716145e-07
+    4.214538200533928e-07
+ 2.88e+10    
+    4.216684147723647e-07
+    1.649648156396822e-07
+    4.170059201481875e-07
+    5.762702353553677e-08
+     1.06033031757195e-07
+    4.165110710941281e-07
+    3.493312567836844e-08
+    5.765772821773215e-08
+    1.653829766989299e-07
+    4.215426144793074e-07
+ 2.89e+10    
+    4.217572487950293e-07
+    1.650370180271656e-07
+    4.170794568994476e-07
+    5.766633858592987e-08
+    1.060895636742298e-07
+     4.16584794738817e-07
+    3.495411023239418e-08
+    5.769681142183418e-08
+    1.654550108168982e-07
+    4.216315858823354e-07
+ 2.9e+10     
+    4.218462592632783e-07
+    1.651092931401407e-07
+    4.171531058979153e-07
+    5.770554630528635e-08
+    1.061460914891039e-07
+    4.166586313324551e-07
+    3.497489601822648e-08
+    5.773578710714086e-08
+    1.655271171306314e-07
+    4.217207349635161e-07
+ 2.91e+10    
+    4.219354468587069e-07
+     1.65181641375087e-07
+    4.172268675960401e-07
+    5.774464686422623e-08
+    1.062026154290279e-07
+    4.167325813256582e-07
+    3.499548334026773e-08
+    5.777465544701164e-08
+    1.655992960377521e-07
+    4.218100624122579e-07
+ 2.92e+10    
+    4.220248122512192e-07
+    1.652540631210444e-07
+    4.173007424385923e-07
+    5.778364042726136e-08
+     1.06259135715977e-07
+    4.168066451610838e-07
+    3.501587249861945e-08
+    5.781341660875557e-08
+    1.656715479284051e-07
+     4.21899568906313e-07
+ 2.93e+10    
+    4.221143560990282e-07
+    1.653265587596295e-07
+    4.173747308627238e-07
+    5.782252715282096e-08
+    1.063156525667517e-07
+    4.168808232734953e-07
+    3.503606378905698e-08
+    5.785207075365609e-08
+    1.657438731852737e-07
+    4.219892551117748e-07
+ 2.94e+10    
+    4.222040790486668e-07
+    1.653991286650511e-07
+    4.174488332980131e-07
+    5.786130719327883e-08
+    1.063721661930355e-07
+    4.169551160898245e-07
+    3.505605750300647e-08
+    5.789061803699601e-08
+    1.658162721835952e-07
+    4.220791216830692e-07
+ 2.95e+10    
+    4.222939817350097e-07
+    1.654717732041306e-07
+    4.175230501665318e-07
+    5.789998069498209e-08
+    1.064286768014554e-07
+    4.170295240292368e-07
+    3.507585392752475e-08
+    5.792905860808516e-08
+    1.658887452911804e-07
+    4.221691692629707e-07
+ 2.96e+10    
+    4.223840647812986e-07
+     1.65544492736321e-07
+    4.175973818828964e-07
+    5.793854779828096e-08
+    1.064851845936404e-07
+    4.171040475031993e-07
+      3.5095453345281e-08
+    5.796739261028852e-08
+    1.659612928684332e-07
+    4.222593984826139e-07
+ 2.97e+10    
+    4.224743287991795e-07
+    1.656172876137309e-07
+    4.176718288543318e-07
+    5.797700863756048e-08
+    1.065416897662806e-07
+    4.171786869155464e-07
+    3.511485603454143e-08
+     5.80056201810565e-08
+    1.660339152683732e-07
+     4.22349809961525e-07
+ 2.98e+10    
+    4.225647743887475e-07
+    1.656901581811459e-07
+    4.177463914807282e-07
+     5.80153633412728e-08
+    1.065981925111857e-07
+    4.172534426625504e-07
+    3.513406226915558e-08
+    5.804374145195592e-08
+    1.661066128366584e-07
+    4.224404043076525e-07
+ 2.99e+10    
+    4.226554021385962e-07
+    1.657631047760559e-07
+    4.178210701547084e-07
+    5.805361203197143e-08
+    1.066546930153442e-07
+    4.173283151329918e-07
+    3.515307231854544e-08
+    5.808175654870276e-08
+    1.661793859116112e-07
+     4.22531182117411e-07
+ 3e+10       
+    4.227462126258772e-07
+    1.658361277286808e-07
+    4.178958652616878e-07
+    5.809175482634633e-08
+    1.067111914609813e-07
+     4.17403304708229e-07
+     3.51718864476963e-08
+    5.811966559119571e-08
+    1.662522348242441e-07
+    4.226221439757304e-07
+ 3.01e+10    
+    4.228372064163622e-07
+    1.659092273619978e-07
+    4.179707771799374e-07
+    5.812979183525991e-08
+    1.067676880256172e-07
+    4.174784117622712e-07
+    3.519050491714987e-08
+     5.81574686935512e-08
+    1.663251598982876e-07
+    4.227132904561101e-07
+ 3.02e+10    
+    4.229283840645168e-07
+    1.659824039917715e-07
+    4.180458062806534e-07
+    5.816772316378488e-08
+    1.068241828821254e-07
+    4.175536366618529e-07
+     3.52089279829996e-08
+     5.81951659641395e-08
+    1.663981614502203e-07
+    4.228046221206867e-07
+ 3.03e+10    
+    4.230197461135737e-07
+    1.660556579265842e-07
+    4.181209529280197e-07
+    5.820554891124219e-08
+    1.068806761987898e-07
+    4.176289797665035e-07
+    3.522715589688776e-08
+    5.823275750562157e-08
+    1.664712397892979e-07
+    4.228961395202977e-07
+ 3.04e+10    
+    4.231112930956173e-07
+    1.661289894678667e-07
+    4.181962174792763e-07
+    5.824326917124083e-08
+    1.069371681393628e-07
+    4.177044414286257e-07
+     3.52451889060046e-08
+    5.827024341498763e-08
+    1.665443952175861e-07
+      4.2298784319456e-07
+ 3.05e+10    
+    4.232030255316677e-07
+    1.662023989099322e-07
+    4.182716002847874e-07
+    5.828088403171814e-08
+    1.069936588631222e-07
+    4.177800219935689e-07
+    3.526302725308952e-08
+    5.830762378359599e-08
+    1.666176280299926e-07
+    4.230797336719507e-07
+ 3.06e+10    
+    4.232949439317765e-07
+    1.662758865400089e-07
+    4.183471016881093e-07
+    5.831839357498115e-08
+    1.070501485249281e-07
+    4.178557217997048e-07
+    3.528067117643378e-08
+    5.834489869721325e-08
+    1.666909385143014e-07
+    4.231718114698904e-07
+ 3.07e+10    
+      4.2338704879512e-07
+    1.663494526382754e-07
+    4.184227220260585e-07
+    5.835579787774877e-08
+    1.071066372752793e-07
+     4.17931541178502e-07
+    3.529812090988551e-08
+    5.838206823605539e-08
+    1.667643269512073e-07
+    4.232640770948384e-07
+ 3.08e+10    
+    4.234793406101003e-07
+    1.664230974778961e-07
+    4.184984616287836e-07
+    5.839309701119488e-08
+    1.071631252603702e-07
+    4.180074804546055e-07
+    3.531537668285592e-08
+    5.841913247482952e-08
+    1.668377936143518e-07
+    4.233565310423835e-07
+ 3.09e+10    
+    4.235718198544508e-07
+    1.664968213250575e-07
+    4.185743208198332e-07
+     5.84302910409923e-08
+    1.072196126221461e-07
+    4.180835399459102e-07
+    3.533243872032767e-08
+    5.845609148277669e-08
+    1.669113387703602e-07
+    4.234491737973468e-07
+ 3.1e+10     
+    4.236644869953452e-07
+    1.665706244390061e-07
+    4.186502999162281e-07
+    5.846738002735731e-08
+    1.072760994983591e-07
+    4.181597199636409e-07
+    3.534930724286471e-08
+    5.849294532371531e-08
+    1.669849626788787e-07
+    4.235420058338851e-07
+ 3.11e+10    
+    4.237573424895063e-07
+    1.666445070720861e-07
+    4.187263992285304e-07
+     5.85043640250951e-08
+    1.073325860226234e-07
+    4.182360208124265e-07
+    3.536598246662371e-08
+    5.852969405608539e-08
+    1.670586655926129e-07
+    4.236350276155973e-07
+ 3.12e+10    
+    4.238503867833219e-07
+    1.667184694697784e-07
+    4.188026190609162e-07
+    5.854124308364579e-08
+    1.073890723244702e-07
+    4.183124427903801e-07
+    3.538246460336723e-08
+    5.856633773299361e-08
+    1.671324477573674e-07
+    4.237282395956372e-07
+ 3.13e+10    
+     4.23943620312963e-07
+    1.667925118707403e-07
+    4.188789597112473e-07
+    5.857801724713115e-08
+     1.07445558529402e-07
+     4.18388986189175e-07
+    3.539875386047823e-08
+    5.860287640225889e-08
+    1.672063094120851e-07
+    4.238216422168261e-07
+ 3.14e+10    
+    4.240370435045042e-07
+    1.668666345068455e-07
+    4.189554214711405e-07
+    5.861468655440207e-08
+    1.075020447589473e-07
+    4.184656512941239e-07
+    3.541485044097629e-08
+     5.86393101064586e-08
+    1.672802507888881e-07
+    4.239152359117705e-07
+ 3.15e+10    
+    4.241306567740437e-07
+    1.669408376032254e-07
+    4.190320046260427e-07
+    5.865125103908637e-08
+     1.07558531130714e-07
+     4.18542438384254e-07
+    3.543075454353515e-08
+    5.867563888297572e-08
+    1.673542721131189e-07
+    4.240090211029816e-07
+ 3.16e+10    
+    4.242244605278303e-07
+    1.670151213783095e-07
+    4.191087094553008e-07
+    5.868771072963739e-08
+     1.07615017758443e-07
+    4.186193477323878e-07
+    3.544646636250161e-08
+    5.871186276404604e-08
+    1.674283736033822e-07
+    4.241029982029993e-07
+ 3.17e+10    
+    4.243184551623883e-07
+    1.670894860438685e-07
+    4.191855362322333e-07
+    5.872406564938304e-08
+    1.076715047520609e-07
+    4.186963796052189e-07
+    3.546198608791598e-08
+    5.874798177680633e-08
+    1.675025554715866e-07
+    4.241971676145128e-07
+ 3.18e+10    
+     4.24412641064647e-07
+    1.671639318050564e-07
+    4.192624852242059e-07
+    5.876031581657533e-08
+    1.077279922177331e-07
+    4.187735342633891e-07
+    3.547731390553377e-08
+    5.878399594334305e-08
+    1.675768179229884e-07
+    4.242915297304913e-07
+ 3.19e+10    
+    4.245070186120685e-07
+    1.672384588604525e-07
+    4.193395566926989e-07
+    5.879646124444034e-08
+    1.077844802579157e-07
+    4.188508119615678e-07
+    3.549244999684864e-08
+    5.881990528074113e-08
+     1.67651161156234e-07
+    4.243860849343085e-07
+ 3.2e+10     
+    4.246015881727809e-07
+    1.673130674021062e-07
+    4.194167508933824e-07
+    5.883250194122885e-08
+    1.078409689714074e-07
+    4.189282129485271e-07
+    3.550739453911685e-08
+     5.88557098011338e-08
+    1.677255853634045e-07
+    4.244808335998764e-07
+ 3.21e+10    
+    4.246963501057078e-07
+    1.673877576155789e-07
+    4.194940680761876e-07
+    5.886843791026693e-08
+    1.078974584534007e-07
+    4.190057374672195e-07
+    3.552214770538243e-08
+    5.889140951175224e-08
+    1.678000907300589e-07
+    4.245757760917707e-07
+ 3.22e+10    
+     4.24791304760704e-07
+    1.674625296799897e-07
+    4.195715084853777e-07
+     5.89042691500077e-08
+    1.079539487955332e-07
+    4.190833857548558e-07
+    3.553670966450427e-08
+    5.892700441497625e-08
+    1.678746774352793e-07
+    4.246709127653688e-07
+ 3.23e+10    
+    4.248864524786863e-07
+    1.675373837680588e-07
+     4.19649072359622e-07
+    5.893999565408248e-08
+     1.08010440085938e-07
+    4.191611580429805e-07
+    3.555108058118373e-08
+    5.896249450838488e-08
+    1.679493456517153e-07
+    4.247662439669796e-07
+ 3.24e+10    
+    4.249817935917702e-07
+    1.676123200461524e-07
+    4.197267599320645e-07
+    5.897561741135317e-08
+    1.080669324092936e-07
+    4.192390545575477e-07
+    3.556526061599373e-08
+    5.899787978480745e-08
+    1.680240955456294e-07
+    4.248617700339783e-07
+ 3.25e+10    
+    4.250773284234039e-07
+    1.676873386743276e-07
+    4.198045714303967e-07
+    5.901113440596422e-08
+    1.081234258468737e-07
+    4.193170755189966e-07
+    3.557924992540883e-08
+    5.903316023237527e-08
+     1.68098927276942e-07
+    4.249574912949412e-07
+ 3.26e+10    
+    4.251730572885031e-07
+    1.677624398063776e-07
+    4.198825070769301e-07
+     5.90465466173957e-08
+    1.081799204765969e-07
+    4.193952211423301e-07
+    3.559304866183645e-08
+    5.906833583457331e-08
+    1.681738409992777e-07
+    4.250534080697809e-07
+ 3.27e+10    
+    4.252689804935858e-07
+    1.678376235898769e-07
+    4.199605670886644e-07
+    5.908185402051579e-08
+    1.082364163730746e-07
+    4.194734916371849e-07
+    3.560665697364904e-08
+     5.91034065702921e-08
+    1.682488368600107e-07
+    4.251495206698833e-07
+ 3.28e+10    
+    4.253650983369099e-07
+    1.679128901662272e-07
+    4.200387516773602e-07
+    5.911705658563418e-08
+    1.082929136076604e-07
+    4.195518872079107e-07
+    3.562007500521724e-08
+    5.913837241388039e-08
+    1.683239150003106e-07
+    4.252458293982399e-07
+ 3.29e+10    
+    4.254614111086052e-07
+    1.679882396707029e-07
+     4.20117061049608e-07
+    5.915215427855535e-08
+     1.08349412248497e-07
+    4.196304080536414e-07
+    3.563330289694423e-08
+    5.917323333519757e-08
+    1.683990755551895e-07
+    4.253423345495866e-07
+ 3.3e+10     
+     4.25557919090811e-07
+    1.680636722324968e-07
+     4.20195495406898e-07
+    5.918714706063222e-08
+    1.084059123605645e-07
+    4.197090543683715e-07
+    3.564634078530077e-08
+    5.920798929966653e-08
+    1.684743186535478e-07
+    4.254390364105396e-07
+ 3.31e+10    
+    4.256546225578086e-07
+    1.681391879747664e-07
+    4.202740549456911e-07
+       5.922203488882e-08
+    1.084624140057271e-07
+    4.197878263410257e-07
+    3.565918880286125e-08
+    5.924264026832666e-08
+    1.685496444182204e-07
+    4.255359352597277e-07
+ 3.32e+10    
+    4.257515217761585e-07
+    1.682147870146801e-07
+    4.203527398574871e-07
+    5.925681771573011e-08
+    1.085189172427799e-07
+    4.198667241555364e-07
+    3.567184707834081e-08
+    5.927718619788728e-08
+    1.686250529660241e-07
+    4.256330313679321e-07
+ 3.33e+10    
+    4.258486170048312e-07
+     1.68290469463463e-07
+    4.204315503288924e-07
+    5.929149548968443e-08
+    1.085754221274947e-07
+     4.19945747990912e-07
+    3.568431573663312e-08
+    5.931162704078086e-08
+     1.68700544407804e-07
+    4.257303249982186e-07
+ 3.34e+10    
+    4.259459084953421e-07
+    1.683662354264437e-07
+    4.205104865416919e-07
+    5.932606815476948e-08
+    1.086319287126662e-07
+    4.200248980213108e-07
+    3.569659489884898e-08
+    5.934596274521666e-08
+    1.687761188484799e-07
+    4.258278164060719e-07
+ 3.35e+10    
+    4.260433964918829e-07
+    1.684420850030999e-07
+    4.205895486729118e-07
+    5.936053565089097e-08
+    1.086884370481566e-07
+    4.201041744161117e-07
+    3.570868468235603e-08
+    5.938019325523451e-08
+    1.688517763870938e-07
+    4.259255058395314e-07
+ 3.36e+10    
+    4.261410812314542e-07
+    1.685180182871049e-07
+    4.206687368948913e-07
+    5.939489791382825e-08
+    1.087449471809413e-07
+    4.201835773399846e-07
+    3.572058520081895e-08
+    5.941431851075861e-08
+    1.689275171168561e-07
+    4.260233935393222e-07
+ 3.37e+10    
+     4.26238962943996e-07
+    1.685940353663753e-07
+    4.207480513753483e-07
+    5.942915487528908e-08
+    1.088014591551528e-07
+     4.20263106952961e-07
+     3.57322965642406e-08
+    5.944833844765148e-08
+    1.690033411251928e-07
+    4.261214797389887e-07
+ 3.38e+10    
+     4.26337041852518e-07
+    1.686701363231152e-07
+    4.208274922774454e-07
+    5.946330646296433e-08
+    1.088579730121243e-07
+    4.203427634105036e-07
+    3.574381887900389e-08
+     5.94822529977681e-08
+    1.690792484937929e-07
+    4.262197646650265e-07
+ 3.39e+10    
+    4.264353181732262e-07
+    1.687463212338641e-07
+    4.209070597598567e-07
+    5.949735260058262e-08
+    1.089144887904341e-07
+    4.204225468635742e-07
+    3.575515224791433e-08
+    5.951606208901005e-08
+    1.691552392986545e-07
+    4.263182485370132e-07
+ 3.4e+10     
+    4.265337921156556e-07
+     1.68822590169543e-07
+    4.209867539768325e-07
+    5.953129320796545e-08
+    1.089710065259478e-07
+    4.205024574587036e-07
+    3.576629677024337e-08
+     5.95497656453795e-08
+    1.692313136101315e-07
+    4.264169315677358e-07
+ 3.41e+10    
+    4.266324638827918e-07
+    1.688989431955001e-07
+    4.210665750782649e-07
+    5.956512820108199e-08
+    1.090275262518616e-07
+    4.205824953380574e-07
+    3.577725254177236e-08
+    5.958336358703387e-08
+    1.693074714929817e-07
+    4.265158139633228e-07
+ 3.42e+10    
+    4.267313336711991e-07
+    1.689753803715577e-07
+    4.211465232097522e-07
+    5.959885749210387e-08
+    1.090840479987437e-07
+    4.206626606395049e-07
+    3.578801965483712e-08
+    5.961685583033972e-08
+    1.693837130064119e-07
+    4.266148959233686e-07
+ 3.43e+10    
+    4.268304016711462e-07
+    1.690519017520586e-07
+    4.212265985126643e-07
+    5.963248098946055e-08
+    1.091405717945772e-07
+    4.207429534966848e-07
+    3.579859819837356e-08
+    5.965024228792757e-08
+    1.694600382041262e-07
+    4.267141776410638e-07
+ 3.44e+10    
+    4.269296680667267e-07
+    1.691285073859114e-07
+     4.21306801124202e-07
+    5.966599859789391e-08
+    1.091970976648003e-07
+    4.208233740390712e-07
+    3.580898825796318e-08
+    5.968352286874582e-08
+    1.695364471343716e-07
+    4.268136593033156e-07
+ 3.45e+10    
+    4.270291330359819e-07
+    1.692051973166375e-07
+     4.21387131177465e-07
+    5.969941021851335e-08
+    1.092536256323475e-07
+    4.209039223920383e-07
+    3.581918991587993e-08
+    5.971669747811545e-08
+     1.69612939839985e-07
+    4.269133410908764e-07
+ 3.46e+10    
+    4.271287967510228e-07
+    1.692819715824164e-07
+    4.214675888015108e-07
+    5.973271574885089e-08
+    1.093101557176908e-07
+    4.209845986769255e-07
+    3.582920325113719e-08
+    5.974976601778419e-08
+    1.696895163584396e-07
+    4.270132231784629e-07
+ 3.47e+10    
+    4.272286593781473e-07
+    1.693588302161321e-07
+    4.215481741214167e-07
+    5.976591508291597e-08
+    1.093666879388786e-07
+    4.210654030111008e-07
+    3.583902833953556e-08
+      5.9782728385981e-08
+    1.697661767218913e-07
+    4.271133057348801e-07
+ 3.48e+10    
+    4.273287210779598e-07
+    1.694357732454189e-07
+    4.216288872583437e-07
+    5.979900811125041e-08
+    1.094232223115761e-07
+    4.211463355080254e-07
+    3.584866525371109e-08
+    5.981558447747035e-08
+     1.69842920957225e-07
+    4.272135889231401e-07
+ 3.49e+10    
+    4.274289820054857e-07
+     1.69512800692707e-07
+    4.217097283295937e-07
+     5.98319947209833e-08
+    1.094797588491042e-07
+    4.212273962773139e-07
+    3.585811406318408e-08
+    5.984833418360665e-08
+     1.69919749086101e-07
+    4.273140729005806e-07
+ 3.5e+10     
+    4.275294423102896e-07
+    1.695899125752679e-07
+    4.217906974486716e-07
+    5.986487479588593e-08
+    1.095362975624782e-07
+    4.213085854247992e-07
+    3.586737483440843e-08
+    5.988097739238836e-08
+    1.699966611250009e-07
+    4.274147578189832e-07
+ 3.51e+10    
+    4.276301021365837e-07
+    1.696671089052603e-07
+    4.218717947253431e-07
+    5.989764821642616e-08
+    1.095928384604463e-07
+    4.213899030525903e-07
+    3.587644763082139e-08
+    5.991351398851229e-08
+    1.700736570852732e-07
+    4.275156438246885e-07
+ 3.52e+10    
+    4.277309616233466e-07
+    1.697443896897755e-07
+    4.219530202656959e-07
+    5.993031485982387e-08
+    1.096493815495275e-07
+    4.214713492591365e-07
+    3.588533251289405e-08
+    5.994594385342783e-08
+    1.701507369731799e-07
+    4.276167310587102e-07
+ 3.53e+10    
+    4.278320209044281e-07
+    1.698217549308823e-07
+    4.220343741721957e-07
+    5.996287460010484e-08
+    1.097059268340491e-07
+    4.215529241392855e-07
+    3.589402953818195e-08
+    5.997826686539095e-08
+    1.702279007899419e-07
+    4.277180196568494e-07
+ 3.54e+10    
+    4.279332801086617e-07
+    1.698992046256725e-07
+    4.221158565437463e-07
+    5.999532730815575e-08
+    1.097624743161839e-07
+    4.216346277843418e-07
+    3.590253876137642e-08
+    6.001048289951828e-08
+    1.703051485317841e-07
+    4.278195097498035e-07
+ 3.55e+10    
+    4.280347393599704e-07
+    1.699767387663054e-07
+    4.221974674757424e-07
+    6.002767285177846e-08
+    1.098190239959865e-07
+    4.217164602821278e-07
+    3.591086023435628e-08
+    6.004259182784096e-08
+    1.703824801899816e-07
+    4.279212014632788e-07
+ 3.56e+10    
+    4.281363987774748e-07
+    1.700543573400537e-07
+    4.222792070601321e-07
+    6.005991109574452e-08
+    1.098755758714303e-07
+    4.217984217170399e-07
+    3.591899400623996e-08
+    6.007459351935877e-08
+    1.704598957509043e-07
+    4.280230949180976e-07
+ 3.57e+10    
+     4.28238258475596e-07
+    1.701320603293469e-07
+    4.223610753854673e-07
+    6.009204190184941e-08
+    1.099321299384429e-07
+    4.218805121701061e-07
+    3.592694012343799e-08
+    6.010648784009349e-08
+    1.705373951960626e-07
+    4.281251902303053e-07
+ 3.58e+10    
+    4.283403185641594e-07
+     1.70209847711817e-07
+    4.224430725369618e-07
+    6.012406512896654e-08
+    1.099886861909416e-07
+    4.219627317190435e-07
+    3.593469862970604e-08
+      6.0138274653143e-08
+    1.706149785021521e-07
+    4.282274875112753e-07
+ 3.59e+10    
+    4.284425791484967e-07
+    1.702877194603421e-07
+    4.225251985965457e-07
+    6.015598063310153e-08
+    1.100452446208689e-07
+    4.220450804383128e-07
+    3.594226956619815e-08
+    6.016995381873444e-08
+    1.706926456410983e-07
+     4.28329986867814e-07
+ 3.6e+10     
+    4.285450403295446e-07
+    1.703656755430917e-07
+    4.226074536429206e-07
+    6.018778826744607e-08
+     1.10101805218227e-07
+    4.221275583991758e-07
+    3.594965297152043e-08
+    6.020152519427796e-08
+    1.707703965801018e-07
+    4.284326884022613e-07
+ 3.61e+10    
+    4.286477022039464e-07
+    1.704437159235698e-07
+     4.22689837751609e-07
+    6.021948788243176e-08
+     1.10158367971112e-07
+    4.222101656697487e-07
+    3.595684888178531e-08
+    6.023298863441995e-08
+    1.708482312816826e-07
+    4.285355922125948e-07
+ 3.62e+10    
+    4.287505648641448e-07
+    1.705218405606594e-07
+    4.227723509950123e-07
+    6.025107932578353e-08
+    1.102149328657482e-07
+    4.222929023150551e-07
+    3.596385733066562e-08
+    6.026434399109608e-08
+     1.70926149703724e-07
+    4.286386983925241e-07
+ 3.63e+10    
+    4.288536283984812e-07
+    1.706000494086664e-07
+    4.228549934424593e-07
+    6.028256244257361e-08
+    1.102714998865213e-07
+    4.223757683970823e-07
+    3.597067834944961e-08
+    6.029559111358464e-08
+    1.710041517995173e-07
+    4.287420070315926e-07
+ 3.64e+10    
+    4.289568928912872e-07
+     1.70678342417363e-07
+    4.229377651602611e-07
+    6.031393707527468e-08
+    1.103280690160122e-07
+    4.224587639748317e-07
+    3.597731196709592e-08
+    6.032672984855932e-08
+    1.710822375178062e-07
+    4.288455182152722e-07
+ 3.65e+10    
+    4.290603584229796e-07
+    1.707567195320317e-07
+     4.23020666211759e-07
+    6.034520306381308e-08
+     1.10384640235029e-07
+    4.225418891043719e-07
+    3.598375821028892e-08
+    6.035776004014198e-08
+    1.711604068028297e-07
+    4.289492320250579e-07
+ 3.66e+10    
+    4.291640250701497e-07
+    1.708351806935084e-07
+    4.231036966573779e-07
+    6.037636024562218e-08
+    1.104412135226404e-07
+    4.226251438388899e-07
+     3.59900171034945e-08
+    6.038868152995551e-08
+    1.712386595943669e-07
+    4.290531485385615e-07
+ 3.67e+10    
+    4.292678929056527e-07
+    1.709137258382254e-07
+    4.231868565546745e-07
+    6.040740845569498e-08
+     1.10497788856207e-07
+    4.227085282287418e-07
+    3.599608866901589e-08
+    6.041949415717604e-08
+    1.713169958277796e-07
+    4.291572678296028e-07
+ 3.68e+10    
+    4.293719619986968e-07
+     1.70992354898255e-07
+    4.232701459583879e-07
+    6.043834752663729e-08
+    1.105543662114138e-07
+     4.22792042321504e-07
+    3.600197292704998e-08
+    6.045019775858558e-08
+    1.713954154340566e-07
+    4.292615899682995e-07
+ 3.69e+10    
+    4.294762324149312e-07
+    1.710710678013519e-07
+    4.233535649204861e-07
+    6.046917728872002e-08
+     1.10610945562301e-07
+    4.228756861620217e-07
+     3.60076698957439e-08
+    6.048079216862399e-08
+    1.714739183398562e-07
+    4.293661150211584e-07
+ 3.7e+10     
+    4.295807042165279e-07
+    1.711498644709962e-07
+     4.23437113490218e-07
+    6.049989756993193e-08
+    1.106675268812952e-07
+    4.229594597924584e-07
+    3.601317959125161e-08
+    6.051127721944116e-08
+    1.715525044675496e-07
+    4.294708430511574e-07
+ 3.71e+10    
+     4.29685377462269e-07
+    1.712287448264362e-07
+     4.23520791714158e-07
+    6.053050819603179e-08
+    1.107241101392404e-07
+    4.230433632523441e-07
+    3.601850202779102e-08
+    6.054165274094884e-08
+    1.716311737352642e-07
+    4.295757741178376e-07
+ 3.72e+10    
+    4.297902522076264e-07
+    1.713077087827305e-07
+    4.236045996362541e-07
+    6.056100899060054e-08
+    1.107806953054281e-07
+    4.231273965786237e-07
+    3.602363721770122e-08
+    6.057191856087237e-08
+    1.717099260569253e-07
+    4.296809082773828e-07
+ 3.73e+10    
+    4.298953285048446e-07
+    1.713867562507903e-07
+    4.236885372978747e-07
+     6.05913997750932e-08
+    1.108372823476271e-07
+    4.232115598057035e-07
+    3.602858517149989e-08
+    6.060207450480217e-08
+    1.717887613423001e-07
+     4.29786245582706e-07
+ 3.74e+10    
+    4.300006064030205e-07
+    1.714658871374218e-07
+     4.23772604737855e-07
+    6.062168036889079e-08
+    1.108938712321138e-07
+    4.232958529654979e-07
+    3.603334589794102e-08
+    6.063212039624514e-08
+    1.718676794970386e-07
+    4.298917860835265e-07
+ 3.75e+10    
+    4.301060859481803e-07
+    1.715451013453678e-07
+    4.238568019925404e-07
+    6.065185058935175e-08
+     1.10950461923701e-07
+    4.233802760874761e-07
+    3.603791940407272e-08
+     6.06620560566758e-08
+     1.71946680422717e-07
+     4.29997529826455e-07
+ 3.76e+10    
+    4.302117671833575e-07
+    1.716243987733499e-07
+    4.239411290958344e-07
+    6.068191025186353e-08
+     1.11007054385767e-07
+    4.234648291987064e-07
+    3.604230569529537e-08
+    6.069188130558734e-08
+    1.720257640168795e-07
+    4.301034768550688e-07
+ 3.77e+10    
+    4.303176501486684e-07
+    1.717037793161104e-07
+    4.240255860792402e-07
+    6.071185916989365e-08
+    1.110636485802846e-07
+    4.235495123239021e-07
+     3.60465047754198e-08
+     6.07215959605425e-08
+    1.721049301730801e-07
+    4.302096272099915e-07
+ 3.78e+10    
+    4.304237348813855e-07
+    1.717832428644524e-07
+    4.241101729719066e-07
+    6.074169715504077e-08
+    1.111202444678489e-07
+    4.236343254854648e-07
+    3.605051664672568e-08
+    6.075119983722401e-08
+    1.721841787809243e-07
+    4.303159809289662e-07
+ 3.79e+10    
+    4.305300214160121e-07
+    1.718627893052829e-07
+    4.241948898006692e-07
+    6.077142401708565e-08
+    1.111768420077062e-07
+    4.237192687035291e-07
+    3.605434131002023e-08
+    6.078069274948519e-08
+     1.72263509726111e-07
+    4.304225380469325e-07
+ 3.8e+10     
+     4.30636509784352e-07
+    1.719424185216532e-07
+    4.242797365900958e-07
+    6.080103956404165e-08
+    1.112334411577809e-07
+    4.238043419960053e-07
+    3.605797876469682e-08
+    6.081007450940023e-08
+    1.723429228904737e-07
+    4.305292985961003e-07
+ 3.81e+10    
+    4.307432000155819e-07
+    1.720221303927996e-07
+    4.243647133625263e-07
+    6.083054360220528e-08
+    1.112900418747033e-07
+    4.238895453786215e-07
+     3.60614290087939e-08
+    6.083934492731416e-08
+     1.72422418152022e-07
+    4.306362626060193e-07
+ 3.82e+10    
+    4.308500921363197e-07
+    1.721019247941852e-07
+    4.244498201381143e-07
+    6.085993593620639e-08
+    1.113466441138369e-07
+    4.239748788649667e-07
+    3.606469203905403e-08
+    6.086850381189267e-08
+    1.725019953849827e-07
+    4.307434301036512e-07
+ 3.83e+10    
+    4.309571861706919e-07
+    1.721818015975397e-07
+    4.245350569348709e-07
+    6.088921636905817e-08
+    1.114032478293046e-07
+    4.240603424665309e-07
+    3.606776785098305e-08
+    6.089755097017202e-08
+    1.725816544598409e-07
+    4.308508011134403e-07
+ 3.84e+10    
+    4.310644821404012e-07
+    1.722617606709009e-07
+    4.246204237687031e-07
+    6.091838470220715e-08
+    1.114598529740162e-07
+    4.241459361927484e-07
+    3.607065643890924e-08
+    6.092648620760823e-08
+    1.726613952433804e-07
+    4.309583756573797e-07
+ 3.85e+10    
+    4.311719800647925e-07
+    1.723418018786544e-07
+    4.247059206534548e-07
+    6.094744073558271e-08
+    1.115164594996935e-07
+    4.242316600510352e-07
+    3.607335779604279e-08
+    6.095530932812644e-08
+    1.727412175987249e-07
+    4.310661537550793e-07
+ 3.86e+10    
+    4.312796799609153e-07
+    1.724219250815741e-07
+     4.24791547600944e-07
+     6.09763842676465e-08
+    1.115730673568971e-07
+    4.243175140468307e-07
+    3.607587191453525e-08
+    6.098402013417008e-08
+    1.728211213853782e-07
+    4.311741354238322e-07
+ 3.87e+10    
+    4.313875818435898e-07
+    1.725021301368629e-07
+    4.248773046210074e-07
+    6.100521509544172e-08
+    1.116296764950516e-07
+    4.244034981836381e-07
+    3.607819878553903e-08
+    6.101261842674951e-08
+    1.729011064592651e-07
+    4.312823206786782e-07
+ 3.88e+10    
+    4.314956857254654e-07
+    1.725824168981919e-07
+    4.249631917215337e-07
+    6.103393301464213e-08
+    1.116862868624711e-07
+    4.244896124630606e-07
+    3.608033839926708e-08
+    6.104110400549095e-08
+    1.729811726727708e-07
+    4.313907095324679e-07
+ 3.89e+10    
+    4.316039916170859e-07
+     1.72662785215741e-07
+    4.250492089085052e-07
+    6.106253781960078e-08
+    1.117428984063844e-07
+    4.245758568848418e-07
+    3.608229074505269e-08
+    6.106947666868469e-08
+    1.730613198747817e-07
+     4.31499301995926e-07
+ 3.9e+10     
+    4.317124995269461e-07
+    1.727432349362377e-07
+    4.251353561860326e-07
+    6.109102930339861e-08
+    1.117995110729592e-07
+    4.246622314469026e-07
+    3.608405581140915e-08
+    6.109773621333336e-08
+    1.731415479107252e-07
+    4.316080980777093e-07
+ 3.91e+10    
+    4.318212094615519e-07
+    1.728237659029982e-07
+    4.252216335563966e-07
+    6.111940725789285e-08
+    1.118561248073277e-07
+    4.247487361453799e-07
+     3.60856335860897e-08
+    6.112588243519998e-08
+    1.732218566226091e-07
+    4.317170977844705e-07
+ 3.92e+10    
+    4.319301214254778e-07
+    1.729043779559649e-07
+    4.253080410200781e-07
+    6.114767147376518e-08
+    1.119127395536095e-07
+    4.248353709746619e-07
+    3.608702405614737e-08
+    6.115391512885583e-08
+     1.73302245849062e-07
+    4.318263011209158e-07
+ 3.93e+10    
+    4.320392354214228e-07
+    1.729850709317477e-07
+    4.253945785758031e-07
+    6.117582174056953e-08
+    1.119693552549371e-07
+    4.249221359274257e-07
+    3.608822720799489e-08
+    6.118183408772788e-08
+     1.73382715425372e-07
+    4.319357080898609e-07
+ 3.94e+10    
+    4.321485514502691e-07
+    1.730658446636617e-07
+    4.254812462205695e-07
+     6.12038578467799e-08
+    1.120259718534782e-07
+    4.250090309946715e-07
+    3.608924302746478e-08
+    6.120963910414627e-08
+    1.734632651835267e-07
+    4.320453186922913e-07
+ 3.95e+10    
+    4.322580695111328e-07
+    1.731466989817667e-07
+    4.255680439496898e-07
+    6.123177957983784e-08
+    1.120825892904599e-07
+    4.250960561657612e-07
+    3.609007149986925e-08
+    6.123732996939141e-08
+    1.735438949522522e-07
+    4.321551329274149e-07
+ 3.96e+10    
+    4.323677896014196e-07
+    1.732276337129064e-07
+    4.256549717568216e-07
+    6.125958672619964e-08
+    1.121392075061921e-07
+    4.251832114284505e-07
+    3.609071261006025e-08
+    6.126490647374092e-08
+    1.736246045570519e-07
+    4.322651507927192e-07
+ 3.97e+10    
+    4.324777117168778e-07
+    1.733086486807467e-07
+    4.257420296340043e-07
+    6.128727907138334e-08
+    1.121958264400897e-07
+    4.252704967689244e-07
+     3.60911663424895e-08
+    6.129236840651635e-08
+    1.737053938202462e-07
+    4.323753722840229e-07
+ 3.98e+10    
+    4.325878358516488e-07
+    1.733897437058151e-07
+    4.258292175716926e-07
+     6.13148564000157e-08
+    1.122524460306959e-07
+    4.253579121718323e-07
+    3.609143268126857e-08
+    6.131971555612967e-08
+    1.737862625610106e-07
+    4.324857973955313e-07
+ 3.99e+10    
+    4.326981619983195e-07
+    1.734709186055377e-07
+    4.259165355587891e-07
+    6.134231849587861e-08
+    1.123090662157046e-07
+    4.254454576203203e-07
+     3.60915116102289e-08
+    6.134694771012949e-08
+    1.738672105954149e-07
+    4.325964261198859e-07
+ 4e+10       
+    4.328086901479701e-07
+    1.735521731942796e-07
+    4.260039835826806e-07
+    6.136966514195547e-08
+    1.123656869319824e-07
+    4.255331330960647e-07
+     3.60914031129817e-08
+     6.13740646552471e-08
+    1.739482377364611e-07
+    4.327072584482151e-07
+ 4.01e+10    
+    4.329194202902256e-07
+    1.736335072833815e-07
+    4.260915616292667e-07
+    6.139689612047737e-08
+    1.124223081155906e-07
+    4.256209385793058e-07
+    3.609110717297818e-08
+    6.140106617744233e-08
+    1.740293437941227e-07
+    4.328182943701865e-07
+ 4.02e+10    
+    4.330303524133023e-07
+    1.737149206811984e-07
+    4.261792696829955e-07
+    6.142401121296901e-08
+    1.124789297018068e-07
+    4.257088740488794e-07
+    3.609062377356938e-08
+    6.142795206194917e-08
+    1.741105285753826e-07
+    4.329295338740547e-07
+ 4.03e+10    
+     4.33141486504055e-07
+    1.737964131931376e-07
+     4.26267107726894e-07
+    6.145101020029414e-08
+    1.125355516251468e-07
+    4.257969394822483e-07
+    3.608995289806611e-08
+    6.145472209332092e-08
+    1.741917918842709e-07
+    4.330409769467076e-07
+ 4.04e+10    
+    4.332528225480231e-07
+    1.738779846216967e-07
+    4.263550757426008e-07
+    6.147789286270128e-08
+    1.125921738193855e-07
+    4.258851348555354e-07
+    3.608909452979889e-08
+    6.148137605547552e-08
+    1.742731335219033e-07
+    4.331526235737166e-07
+ 4.05e+10    
+     4.33364360529478e-07
+    1.739596347665009e-07
+     4.26443173710396e-07
+    6.150465897986864e-08
+    1.126487962175781e-07
+    4.259734601435533e-07
+    3.608804865217786e-08
+    6.150791373174034e-08
+     1.74354553286519e-07
+    4.332644737393813e-07
+ 4.06e+10    
+    4.334761004314661e-07
+    1.740413634243411e-07
+    4.265314016092327e-07
+    6.153130833094935e-08
+    1.127054187520808e-07
+    4.260619153198362e-07
+    3.608681524875246e-08
+    6.153433490489699e-08
+    1.744360509735185e-07
+    4.333765274267751e-07
+ 4.07e+10    
+    4.335880422358539e-07
+    1.741231703892113e-07
+    4.266197594167679e-07
+    6.155784069461596e-08
+    1.127620413545713e-07
+    4.261505003566692e-07
+    3.608539430327138e-08
+    6.156063935722554e-08
+    1.745176263755013e-07
+    4.334887846177919e-07
+ 4.08e+10    
+    4.337001859233682e-07
+    1.742050554523451e-07
+    4.267082471093911e-07
+    6.158425584910492e-08
+    1.128186639560693e-07
+    4.262392152251191e-07
+    3.608378579974192e-08
+     6.15868268705488e-08
+     1.74599279282303e-07
+    4.336012452931858e-07
+ 4.09e+10    
+    4.338125314736434e-07
+    1.742870184022542e-07
+    4.267968646622557e-07
+    6.161055357226095e-08
+    1.128752864869568e-07
+    4.263280598950633e-07
+    3.608198972248985e-08
+    6.161289722627636e-08
+     1.74681009481033e-07
+    4.337139094326183e-07
+ 4.1e+10     
+    4.339250788652596e-07
+    1.743690590247649e-07
+    4.268856120493077e-07
+    6.163673364158113e-08
+    1.129319088769977e-07
+    4.264170343352205e-07
+    3.608000605621889e-08
+     6.16388502054483e-08
+    1.747628167561123e-07
+    4.338267770146991e-07
+ 4.11e+10    
+    4.340378280757836e-07
+    1.744511771030548e-07
+    4.269744892433124e-07
+    6.166279583425823e-08
+    1.129885310553575e-07
+    4.265061385131764e-07
+    3.607783478606996e-08
+    6.166468558877852e-08
+    1.748447008893094e-07
+    4.339398480170276e-07
+ 4.12e+10    
+    4.341507790818107e-07
+    1.745333724176904e-07
+    4.270634962158883e-07
+    6.168873992722491e-08
+    1.130451529506232e-07
+    4.265953723954164e-07
+    3.607547589768073e-08
+    6.169040315669821e-08
+    1.749266616597786e-07
+    4.340531224162333e-07
+ 4.13e+10    
+    4.342639318590026e-07
+     1.74615644746663e-07
+    4.271526329375283e-07
+    6.171456569719625e-08
+     1.13101774490822e-07
+     4.26684735947349e-07
+    3.607292937724465e-08
+    6.171600268939872e-08
+    1.750086988440961e-07
+    4.341666001880165e-07
+ 4.14e+10    
+    4.343772863821267e-07
+     1.74697993865426e-07
+    4.272418993776348e-07
+    6.174027292071347e-08
+    1.131583956034414e-07
+    4.267742291333382e-07
+    3.607019521157018e-08
+    6.174148396687447e-08
+    1.750908122162972e-07
+    4.342802813071873e-07
+ 4.15e+10    
+    4.344908426250947e-07
+    1.747804195469311e-07
+    4.273312955045404e-07
+    6.176586137418629e-08
+    1.132150162154466e-07
+    4.268638519167277e-07
+    3.606727338813981e-08
+    6.176684676896536e-08
+    1.751730015479129e-07
+     4.34394165747706e-07
+ 4.16e+10    
+    4.346046005609989e-07
+    1.748629215616643e-07
+      4.2742082128554e-07
+    6.179133083393559e-08
+    1.132716362533004e-07
+    4.269536042598676e-07
+    3.606416389516874e-08
+    6.179209087539913e-08
+    1.752552666080061e-07
+    4.345082534827174e-07
+ 4.17e+10    
+    4.347185601621496e-07
+    1.749454996776834e-07
+     4.27510476686916e-07
+    6.181668107623586e-08
+    1.133282556429814e-07
+    4.270434861241449e-07
+    3.606086672166384e-08
+    6.181721606583342e-08
+    1.753376071632084e-07
+    4.346225444845902e-07
+ 4.18e+10    
+     4.34832721400111e-07
+    1.750281536606526e-07
+    4.276002616739642e-07
+    6.184191187735707e-08
+    1.133848743100022e-07
+    4.271334974700048e-07
+    3.605738185748213e-08
+    6.184222211989762e-08
+    1.754200229777563e-07
+    4.347370387249561e-07
+ 4.19e+10    
+    4.349470842457366e-07
+    1.751108832738795e-07
+    4.276901762110201e-07
+    6.186702301360667e-08
+    1.134414921794274e-07
+    4.272236382569806e-07
+    3.605370929338923e-08
+    6.186710881723433e-08
+    1.755025138135275e-07
+    4.348517361747402e-07
+ 4.2e+10     
+    4.350616486692044e-07
+    1.751936882783506e-07
+    4.277802202614867e-07
+    6.189201426137095e-08
+    1.134981091758917e-07
+    4.273139084437183e-07
+    3.604984902111773e-08
+    6.189187593754085e-08
+    1.755850794300767e-07
+    4.349666368042015e-07
+ 4.21e+10    
+    4.351764146400503e-07
+    1.752765684327674e-07
+    4.278703937878568e-07
+    6.191688539715663e-08
+    1.135547252236174e-07
+    4.274043079879998e-07
+    3.604580103342527e-08
+    6.191652326061008e-08
+    1.756677195846715e-07
+    4.350817405829636e-07
+ 4.22e+10    
+    4.352913821272026e-07
+    1.753595234935818e-07
+      4.2796069675174e-07
+    6.194163619763165e-08
+    1.136113402464326e-07
+    4.274948368467721e-07
+    3.604156532415256e-08
+    6.194105056637165e-08
+     1.75750434032329e-07
+    4.351970474800529e-07
+ 4.23e+10    
+    4.354065510990139e-07
+    1.754425532150316e-07
+    4.280511291138894e-07
+    6.196626643966621e-08
+    1.136679541677877e-07
+    4.275854949761687e-07
+    3.603714188828116e-08
+    6.196545763493211e-08
+    1.758332225258502e-07
+    4.353125574639271e-07
+ 4.24e+10    
+    4.355219215232952e-07
+    1.755256573491764e-07
+    4.281416908342219e-07
+    6.199077590037324e-08
+     1.13724566910773e-07
+    4.276762823315345e-07
+    3.603253072199112e-08
+    6.198974424661564e-08
+    1.759160848158568e-07
+    4.354282705025133e-07
+ 4.25e+10    
+    4.356374933673462e-07
+    1.756088356459322e-07
+    4.282323818718461e-07
+    6.201516435714874e-08
+    1.137811783981357e-07
+    4.277671988674511e-07
+    3.602773182271846e-08
+    6.201391018200399e-08
+    1.759990206508262e-07
+    4.355441865632366e-07
+ 4.26e+10    
+    4.357532665979879e-07
+    1.756920878531072e-07
+    4.283232021850852e-07
+    6.203943158771194e-08
+    1.138377885522971e-07
+    4.278582445377604e-07
+    3.602274518921237e-08
+    6.203795522197635e-08
+    1.760820297771266e-07
+     4.35660305613053e-07
+ 4.27e+10    
+    4.358692411815925e-07
+    1.757754137164363e-07
+    4.284141517314996e-07
+    6.206357737014492e-08
+    1.138943972953684e-07
+    4.279494192955873e-07
+    3.601757082159233e-08
+    6.206187914774896e-08
+    1.761651119390525e-07
+    4.357766276184807e-07
+ 4.28e+10    
+    4.359854170841141e-07
+    1.758588129796169e-07
+    4.285052304679129e-07
+     6.20876014829325e-08
+    1.139510045491681e-07
+    4.280407230933637e-07
+    3.601220872140492e-08
+    6.208568174091457e-08
+    1.762482668788601e-07
+    4.358931525456315e-07
+ 4.29e+10    
+     4.36101794271118e-07
+    1.759422853843428e-07
+     4.28596438350432e-07
+    6.211150370500109e-08
+    1.140076102352374e-07
+      4.2813215588285e-07
+    3.600665889168043e-08
+    6.210936278348126e-08
+    1.763314943368017e-07
+    4.360098803602389e-07
+ 4.3e+10     
+    4.362183727078114e-07
+    1.760258306703394e-07
+     4.28687775334472e-07
+    6.213528381575824e-08
+    1.140642142748575e-07
+    4.282237176151607e-07
+    3.600092133698942e-08
+    6.213292205791162e-08
+     1.76414794051161e-07
+    4.361268110276907e-07
+ 4.31e+10    
+    4.363351523590705e-07
+    1.761094485753984e-07
+    4.287792413747785e-07
+     6.21589415951311e-08
+    1.141208165890644e-07
+    4.283154082407832e-07
+    3.599499606349878e-08
+    6.215635934716125e-08
+    1.764981657582876e-07
+    4.362439445130542e-07
+ 4.32e+10    
+    4.364521331894693e-07
+    1.761931388354122e-07
+    4.288708364254499e-07
+    6.218247682360521e-08
+    1.141774170986656e-07
+    4.284072277096038e-07
+    3.598888307902777e-08
+    6.217967443471704e-08
+    1.765816091926323e-07
+    4.363612807811086e-07
+ 4.33e+10    
+    4.365693151633076e-07
+    1.762769011844076e-07
+    4.289625604399567e-07
+     6.22058892822624e-08
+    1.142340157242552e-07
+    4.284991759709255e-07
+    3.598258239310376e-08
+    6.220286710463522e-08
+    1.766651240867803e-07
+    4.364788197963709e-07
+ 4.34e+10    
+    4.366866982446383e-07
+    1.763607353545812e-07
+    4.290544133711693e-07
+    6.222917875281941e-08
+      1.1429061238623e-07
+    4.285912529734922e-07
+    3.597609401701771e-08
+    6.222593714157945e-08
+    1.767487101714873e-07
+     4.36596561523124e-07
+ 4.35e+10    
+    4.368042823972952e-07
+    1.764446410763329e-07
+    4.291463951713731e-07
+    6.225234501766514e-08
+     1.14347207004804e-07
+    4.286834586655097e-07
+    3.596941796387947e-08
+    6.224888433085818e-08
+    1.768323671757121e-07
+    4.367145059254441e-07
+ 4.36e+10    
+    4.369220675849171e-07
+    1.765286180782996e-07
+     4.29238505792295e-07
+    6.227538785989845e-08
+    1.144037995000246e-07
+    4.287757929946663e-07
+    3.596255424867271e-08
+    6.227170845846209e-08
+    1.769160948266524e-07
+    4.368326529672275e-07
+ 4.37e+10    
+    4.370400537709764e-07
+    1.766126660873896e-07
+    4.293307451851189e-07
+     6.22983070633653e-08
+    1.144603897917868e-07
+    4.288682559081534e-07
+    3.595550288830968e-08
+    6.229440931110114e-08
+    1.769998928497773e-07
+    4.369510026122158e-07
+ 4.38e+10    
+    4.371582409188017e-07
+    1.766967848288162e-07
+    4.294231133005129e-07
+    6.232110241269574e-08
+    1.145169777998483e-07
+    4.289608473526863e-07
+    3.594826390168566e-08
+    6.231698667624138e-08
+    1.770837609688622e-07
+    4.370695548240236e-07
+ 4.39e+10    
+    4.372766289916077e-07
+    1.767809740261311e-07
+    4.295156100886434e-07
+    6.234377369334081e-08
+    1.145735634438448e-07
+    4.290535672745252e-07
+     3.59408373097332e-08
+    6.233944034214151e-08
+    1.771676989060228e-07
+    4.371883095661619e-07
+ 4.4e+10     
+    4.373952179525143e-07
+    1.768652334012586e-07
+     4.29608235499201e-07
+    6.236632069160879e-08
+    1.146301466433038e-07
+    4.291464156194945e-07
+    3.593322313547599e-08
+    6.236177009788935e-08
+    1.772517063817477e-07
+    4.373072668020643e-07
+ 4.41e+10    
+    4.375140077645738e-07
+    1.769495626745278e-07
+    4.297009894814163e-07
+    6.238874319470143e-08
+    1.146867273176593e-07
+    4.292393923330013e-07
+    3.592542140408246e-08
+    6.238397573343754e-08
+    1.773357831149328e-07
+    4.374264264951105e-07
+ 4.42e+10    
+    4.376329983907959e-07
+    1.770339615647068e-07
+    4.297938719840811e-07
+    6.241104099075014e-08
+    1.147433053862663e-07
+    4.293324973600585e-07
+    3.591743214291924e-08
+    6.240605703963974e-08
+    1.774199288229148e-07
+    4.375457886086521e-07
+ 4.43e+10    
+    4.377521897941691e-07
+    1.771184297890362e-07
+    4.298868829555695e-07
+    6.243321386885145e-08
+    1.147998807684149e-07
+    4.294257306453009e-07
+    3.590925538160407e-08
+    6.242801380828582e-08
+    1.775041432215037e-07
+    4.376653531060345e-07
+ 4.44e+10    
+     4.37871581937685e-07
+    1.772029670632605e-07
+    4.299800223438545e-07
+    6.245526161910241e-08
+    1.148564533833441e-07
+     4.29519092133006e-07
+    3.590089115205858e-08
+    6.244984583213738e-08
+    1.775884260250174e-07
+    4.377851199506218e-07
+ 4.45e+10    
+    4.379911747843599e-07
+    1.772875731016628e-07
+    4.300732900965294e-07
+    6.247718403263585e-08
+    1.149130231502557e-07
+    4.296125817671115e-07
+    3.589233948856071e-08
+    6.247155290496249e-08
+    1.776727769463128e-07
+    4.379050891058168e-07
+ 4.46e+10    
+    4.381109682972586e-07
+    1.773722476170962e-07
+     4.30166686160825e-07
+    6.249898090165521e-08
+    1.149695899883282e-07
+    4.297061994912353e-07
+    3.588360042779683e-08
+    6.249313482157074e-08
+    1.777571956968208e-07
+    4.380252605350884e-07
+ 4.47e+10    
+    4.382309624395165e-07
+    1.774569903210176e-07
+    4.302602104836293e-07
+    6.252065201946925e-08
+    1.150261538167303e-07
+    4.297999452486935e-07
+    3.587467400891357e-08
+    6.251459137784751e-08
+    1.778416819865776e-07
+    4.381456342019899e-07
+ 4.48e+10    
+    4.383511571743592e-07
+    1.775418009235189e-07
+    4.303538630115051e-07
+    6.254219718052623e-08
+    1.150827145546342e-07
+    4.298938189825191e-07
+    3.586556027356919e-08
+    6.253592237078827e-08
+    1.779262355242581e-07
+    4.382662100701819e-07
+ 4.49e+10    
+    4.384715524651261e-07
+    1.776266791333606e-07
+    4.304476436907095e-07
+    6.256361618044811e-08
+    1.151392721212293e-07
+    4.299878206354784e-07
+    3.585625926598472e-08
+    6.255712759853248e-08
+    1.780108560172083e-07
+    4.383869881034534e-07
+ 4.5e+10     
+    4.385921482752906e-07
+    1.777116246580034e-07
+    4.305415524672099e-07
+    6.258490881606445e-08
+    1.151958264357351e-07
+    4.300819501500908e-07
+    3.584677103299485e-08
+     6.25782068603973e-08
+    1.780955431714778e-07
+    4.385079682657443e-07
+ 4.51e+10    
+    4.387129445684801e-07
+    1.777966372036401e-07
+    4.306355892867039e-07
+    6.260607488544558e-08
+    1.152523774174139e-07
+    4.301762074686445e-07
+    3.583709562409825e-08
+    6.259915995691107e-08
+    1.781802966918517e-07
+    4.386291505211646e-07
+ 4.52e+10    
+    4.388339413084971e-07
+    1.778817164752286e-07
+    4.307297540946358e-07
+    6.262711418793645e-08
+    1.153089249855846e-07
+    4.302705925332157e-07
+     3.58272330915077e-08
+     6.26199866898464e-08
+    1.782651162818834e-07
+    4.387505348340158e-07
+ 4.53e+10    
+    4.389551384593392e-07
+    1.779668621765225e-07
+    4.308240468362138e-07
+    6.264802652418913e-08
+    1.153654690596348e-07
+    4.303651052856845e-07
+    3.581718349019987e-08
+    6.264068686225305e-08
+    1.783500016439262e-07
+    4.388721211688101e-07
+ 4.54e+10    
+    4.390765359852183e-07
+    1.780520740101036e-07
+     4.30918467456427e-07
+    6.266881169619572e-08
+    1.154220095590334e-07
+    4.304597456677528e-07
+    3.580694687796461e-08
+    6.266126027849056e-08
+    1.784349524791652e-07
+    4.389939094902914e-07
+ 4.55e+10    
+    4.391981338505804e-07
+    1.781373516774131e-07
+    4.310130159000631e-07
+    6.268946950732087e-08
+    1.154785464033438e-07
+     4.30554513620959e-07
+    3.579652331545397e-08
+    6.268170674426061e-08
+    1.785199684876492e-07
+    4.391158997634535e-07
+ 4.56e+10    
+    4.393199320201239e-07
+    1.782226948787834e-07
+    4.311076921117259e-07
+    6.270999976233397e-08
+    1.155350795122357e-07
+    4.306494090866983e-07
+     3.57859128662309e-08
+    6.270202606663921e-08
+    1.786050493683227e-07
+    4.392380919535604e-07
+ 4.57e+10    
+    4.394419304588198e-07
+    1.783081033134696e-07
+    4.312024960358491e-07
+    6.273040226744084e-08
+    1.155916088054973e-07
+    4.307444320062348e-07
+    3.577511559681745e-08
+    6.272221805410826e-08
+    1.786901948190564e-07
+    4.393604860261642e-07
+ 4.58e+10    
+     4.39564129131928e-07
+    1.783935766796795e-07
+    4.312974276167162e-07
+    6.275067683031558e-08
+    1.156481342030482e-07
+    4.308395823207214e-07
+    3.576413157674248e-08
+     6.27422825165873e-08
+    1.787754045366796e-07
+    4.394830819471236e-07
+ 4.59e+10    
+    4.396865280050171e-07
+     1.78479114674606e-07
+    4.313924867984727e-07
+    6.277082326013191e-08
+    1.157046556249504e-07
+    4.309348599712129e-07
+    3.575296087858947e-08
+    6.276221926546472e-08
+    1.788606782170109e-07
+    4.396058796826233e-07
+ 4.6e+10     
+    4.398091270439825e-07
+    1.785647169944574e-07
+    4.314876735251469e-07
+    6.279084136759412e-08
+    1.157611729914212e-07
+    4.310302648986842e-07
+    3.574160357804323e-08
+    6.278202811362866e-08
+    1.789460155548892e-07
+    4.397288791991901e-07
+ 4.61e+10    
+    4.399319262150624e-07
+    1.786503833344881e-07
+     4.31582987740661e-07
+    6.281073096496806e-08
+    1.158176862228443e-07
+    4.311257970440442e-07
+    3.573005975393686e-08
+    6.280170887549799e-08
+    1.790314162442051e-07
+    4.398520804637127e-07
+ 4.62e+10    
+    4.400549254848563e-07
+    1.787361133890293e-07
+    4.316784293888503e-07
+    6.283049186611151e-08
+    1.158741952397817e-07
+    4.312214563481517e-07
+    3.571832948829778e-08
+    6.282126136705243e-08
+    1.791168799779313e-07
+    4.399754834434568e-07
+ 4.63e+10    
+    4.401781248203414e-07
+    1.788219068515199e-07
+    4.317739984134767e-07
+    6.285012388650444e-08
+    1.159306999629854e-07
+    4.313172427518308e-07
+     3.57064128663937e-08
+    6.284068540586294e-08
+    1.792024064481533e-07
+    4.400990881060838e-07
+ 4.64e+10    
+    4.403015241888904e-07
+    1.789077634145356e-07
+    4.318696947582442e-07
+     6.28696268432791e-08
+    1.159872003134084e-07
+    4.314131561958861e-07
+    3.569430997677808e-08
+    6.285998081112157e-08
+    1.792879953461003e-07
+    4.402228944196676e-07
+ 4.65e+10    
+    4.404251235582861e-07
+    1.789936827698208e-07
+    4.319655183668152e-07
+    6.288900055524961e-08
+    1.160436962122167e-07
+    4.315091966211194e-07
+    3.568202091133502e-08
+      6.2879147403671e-08
+     1.79373646362175e-07
+    4.403469023527092e-07
+ 4.66e+10    
+    4.405489228967399e-07
+    1.790796646083172e-07
+    4.320614691828232e-07
+    6.290824484294134e-08
+    1.161001875807996e-07
+     4.31605363968339e-07
+    3.566954576532396e-08
+    6.289818500603406e-08
+    1.794593591859842e-07
+    4.404711118741565e-07
+ 4.67e+10    
+    4.406729221729063e-07
+    1.791657086201944e-07
+    4.321575471498902e-07
+    6.292735952862022e-08
+    1.161566743407817e-07
+    4.317016581783805e-07
+    3.565688463742371e-08
+    6.291709344244266e-08
+    1.795451335063689e-07
+    4.405955229534159e-07
+ 4.68e+10    
+    4.407971213558977e-07
+    1.792518144948795e-07
+    4.322537522116396e-07
+    6.294634443632126e-08
+    1.162131564140332e-07
+    4.317980791921179e-07
+    3.564403762977622e-08
+    6.293587253886651e-08
+    1.796309690114341e-07
+    4.407201355603716e-07
+ 4.69e+10    
+     4.40921520415303e-07
+    1.793379819210868e-07
+    4.323500843117105e-07
+    6.296519939187747e-08
+     1.16269633722681e-07
+    4.318946269504778e-07
+     3.56310048480298e-08
+    6.295452212304191e-08
+    1.797168653885785e-07
+    4.408449496654002e-07
+ 4.7e+10     
+    4.410461193211995e-07
+    1.794242105868468e-07
+    4.324465433937733e-07
+    6.298392422294789e-08
+    1.163261061891194e-07
+     4.31991301394455e-07
+    3.561778640138195e-08
+     6.29730420244997e-08
+    1.798028223245245e-07
+    4.409699652393849e-07
+ 4.71e+10    
+    4.411709180441705e-07
+    1.795105001795362e-07
+    4.325431294015418e-07
+    6.300251875904569e-08
+     1.16382573736021e-07
+    4.320881024651249e-07
+    3.560438240262171e-08
+    6.299143207459334e-08
+    1.798888395053473e-07
+    4.410951822537316e-07
+ 4.72e+10    
+    4.412959165553175e-07
+    1.795968503859065e-07
+    4.326398422787898e-07
+    6.302098283156591e-08
+    1.164390362863468e-07
+    4.321850301036588e-07
+    3.559079296817147e-08
+    6.300969210652654e-08
+    1.799749166165044e-07
+    4.412206006803822e-07
+ 4.73e+10    
+    4.414211148262771e-07
+    1.796832608921132e-07
+    4.327366819693619e-07
+    6.303931627381273e-08
+    1.164954937633567e-07
+    4.322820842513356e-07
+    3.557701821812848e-08
+    6.302782195538077e-08
+    1.800610533428648e-07
+    4.413462204918324e-07
+ 4.74e+10    
+    4.415465128292334e-07
+    1.797697313837444e-07
+    4.328336484171895e-07
+    6.305751892102681e-08
+    1.165519460906201e-07
+    4.323792648495563e-07
+    3.556305827630579e-08
+    6.304582145814217e-08
+    1.801472493687381e-07
+    4.414720416611415e-07
+ 4.75e+10    
+    4.416721105369328e-07
+    1.798562615458497e-07
+    4.329307415663025e-07
+    6.307559061041196e-08
+    1.166083931920255e-07
+    4.324765718398576e-07
+    3.554891327027263e-08
+    6.306369045372842e-08
+     1.80233504377903e-07
+    4.415980641619497e-07
+ 4.76e+10    
+    4.417979079226991e-07
+     1.79942851062969e-07
+    4.330279613608435e-07
+    6.309353118116186e-08
+    1.166648349917915e-07
+    4.325740051639246e-07
+    3.553458333139457e-08
+    6.308142878301549e-08
+    1.803198180536365e-07
+    4.417242879684916e-07
+ 4.77e+10    
+    4.419239049604446e-07
+    1.800294996191603e-07
+    4.331253077450818e-07
+    6.311134047448625e-08
+    1.167212714144759e-07
+    4.326715647636032e-07
+    3.552006859487281e-08
+    6.309903628886362e-08
+     1.80406190078742e-07
+    4.418507130556077e-07
+ 4.78e+10    
+    4.420501016246846e-07
+     1.80116206898028e-07
+    4.332227806634244e-07
+    6.312901833363697e-08
+     1.16777702384986e-07
+    4.327692505809145e-07
+    3.550536919978344e-08
+    6.311651281614349e-08
+    1.804926201355785e-07
+    4.419773393987609e-07
+ 4.79e+10    
+    4.421764978905515e-07
+    1.802029725827511e-07
+    4.333203800604297e-07
+    6.314656460393351e-08
+     1.16834127828588e-07
+    4.328670625580652e-07
+    3.549048528911567e-08
+    6.313385821176179e-08
+    1.805791079060877e-07
+    4.421041669740476e-07
+ 4.8e+10     
+    4.423030937338064e-07
+    1.802897963561113e-07
+    4.334181058808207e-07
+    6.316397913278861e-08
+    1.168905476709173e-07
+    4.329650006374615e-07
+    3.547541700981013e-08
+    6.315107232468659e-08
+    1.806656530718226e-07
+    4.422311957582093e-07
+ 4.81e+10    
+    4.424298891308523e-07
+    1.803766779005204e-07
+    4.335159580694975e-07
+    6.318126176973338e-08
+    1.169469618379876e-07
+    4.330630647617223e-07
+    3.546016451279623e-08
+    6.316815500597267e-08
+    1.807522553139759e-07
+    4.423584257286497e-07
+ 4.82e+10    
+    4.425568840587475e-07
+    1.804636168980477e-07
+    4.336139365715484e-07
+    6.319841236644189e-08
+    1.170033702562001e-07
+    4.331612548736897e-07
+    3.544472795302913e-08
+    6.318510610878608e-08
+     1.80838914313407e-07
+     4.42485856863443e-07
+ 4.83e+10    
+    4.426840784952156e-07
+    1.805506130304476e-07
+    4.337120413322637e-07
+    6.321543077675599e-08
+    1.170597728523536e-07
+    4.332595709164409e-07
+    3.542910748952636e-08
+    6.320192548842881e-08
+    1.809256297506697e-07
+    4.426134891413486e-07
+ 4.84e+10    
+    4.428114724186607e-07
+    1.806376659791873e-07
+    4.338102722971478e-07
+    6.323231685670936e-08
+    1.171161695536531e-07
+    4.333580128333031e-07
+     3.54133032854037e-08
+    6.321861300236309e-08
+    1.810124013060403e-07
+    4.427413225418223e-07
+ 4.85e+10    
+     4.42939065808176e-07
+    1.807247754254722e-07
+    4.339086294119277e-07
+    6.324907046455153e-08
+    1.171725602877191e-07
+    4.334565805678618e-07
+    3.539731550791062e-08
+    6.323516851023523e-08
+    1.810992286595438e-07
+    4.428693570450284e-07
+ 4.86e+10    
+    4.430668586435595e-07
+    1.808119410502757e-07
+     4.34007112622572e-07
+    6.326569146077165e-08
+    1.172289449825968e-07
+    4.335552740639739e-07
+    3.538114432846526e-08
+     6.32515918738994e-08
+    1.811861114909818e-07
+    4.429975926318516e-07
+ 4.87e+10    
+    4.431948509053201e-07
+    1.808991625343624e-07
+    4.341057218752948e-07
+     6.32821797081215e-08
+    1.172853235667649e-07
+    4.336540932657799e-07
+    3.536478992268871e-08
+    6.326788295744084e-08
+    1.812730494799589e-07
+     4.43126029283908e-07
+ 4.88e+10    
+    4.433230425746955e-07
+    1.809864395583175e-07
+    4.342044571165724e-07
+    6.329853507163904e-08
+    1.173416959691444e-07
+    4.337530381177134e-07
+    3.534825247043898e-08
+    6.328404162719917e-08
+    1.813600423059098e-07
+    4.432546669835565e-07
+ 4.89e+10    
+    4.434514336336585e-07
+    1.810737718025715e-07
+    4.343033182931515e-07
+    6.331475741867084e-08
+    1.173980621191077e-07
+    4.338521085645151e-07
+     3.53315321558443e-08
+    6.330006775179113e-08
+    1.814470896481258e-07
+    4.433835057139122e-07
+ 4.9e+10     
+     4.43580024064928e-07
+    1.811611589474272e-07
+    4.344023053520635e-07
+    6.333084661889461e-08
+    1.174544219464865e-07
+    4.339513045512413e-07
+     3.53146291673357e-08
+    6.331596120213289e-08
+    1.815341911857807e-07
+    4.435125454588522e-07
+ 4.91e+10    
+    4.437088138519838e-07
+    1.812486006730851e-07
+    4.345014182406338e-07
+    6.334680254434148e-08
+    1.175107753815811e-07
+    4.340506260232758e-07
+    3.529754369767947e-08
+     6.33317218514625e-08
+    1.816213465979576e-07
+    4.436417862030325e-07
+ 4.92e+10    
+    4.438378029790722e-07
+      1.8133609665967e-07
+    4.346006569064915e-07
+    6.336262506941787e-08
+    1.175671223551684e-07
+    4.341500729263419e-07
+     3.52802759440087e-08
+    6.334734957536173e-08
+    1.817085555636748e-07
+    4.437712279318935e-07
+ 4.93e+10    
+    4.439669914312204e-07
+     1.81423646587256e-07
+     4.34700021297584e-07
+    6.337831407092689e-08
+    1.176234627985103e-07
+    4.342496452065103e-07
+    3.526282610785435e-08
+    6.336284425177764e-08
+    1.817958177619113e-07
+    4.439008706316733e-07
+ 4.94e+10    
+    4.440963791942446e-07
+    1.815112501358925e-07
+    4.347995113621845e-07
+    6.339386942808995e-08
+    1.176797966433624e-07
+    4.343493428102133e-07
+    3.524519439517587e-08
+    6.337820576104407e-08
+    1.818831328716332e-07
+    4.440307142894182e-07
+ 4.95e+10    
+    4.442259662547597e-07
+    1.815989069856286e-07
+    4.348991270489038e-07
+     6.34092910225675e-08
+    1.177361238219813e-07
+    4.344491656842529e-07
+     3.52273810163911e-08
+    6.339343398590241e-08
+    1.819705005718183e-07
+    4.441607588929899e-07
+ 4.96e+10    
+    4.443557526001909e-07
+    1.816866168165395e-07
+    4.349988683067002e-07
+     6.34245787384798e-08
+    1.177924442671332e-07
+    4.345491137758105e-07
+    3.520938618640576e-08
+     6.34085288115226e-08
+     1.82057920541482e-07
+    4.442910044310779e-07
+ 4.97e+10    
+    4.444857382187827e-07
+    1.817743793087506e-07
+    4.350987350848923e-07
+    6.343973246242727e-08
+    1.178487579121022e-07
+    4.346491870324595e-07
+    3.519121012464222e-08
+    6.342349012552348e-08
+    1.821453924597024e-07
+    4.444214508932082e-07
+ 4.98e+10    
+    4.446159230996072e-07
+    1.818621941424622e-07
+    4.351987273331641e-07
+    6.345475208351072e-08
+    1.179050646906971e-07
+    4.347493854021747e-07
+    3.517285305506778e-08
+    6.343831781799293e-08
+    1.822329160056451e-07
+    4.445520982697539e-07
+ 4.99e+10    
+    4.447463072325755e-07
+    1.819500609979748e-07
+    4.352988450015816e-07
+    6.346963749335094e-08
+    1.179613645372603e-07
+    4.348497088333394e-07
+     3.51543152062223e-08
+    6.345301178150764e-08
+    1.823204908585877e-07
+    4.446829465519417e-07
+ 5e+10       
+     4.44876890608445e-07
+    1.820379795557125e-07
+     4.35399088040597e-07
+    6.348438858610845e-08
+    1.180176573866747e-07
+    4.349501572747602e-07
+    3.513559681124543e-08
+    6.346757191115292e-08
+    1.824081166979453e-07
+    4.448139957318654e-07
+ 5.01e+10    
+    4.450076732188301e-07
+    1.821259494962483e-07
+    4.354994564010626e-07
+    6.349900525850236e-08
+    1.180739431743716e-07
+     4.35050730675672e-07
+    3.511669810790292e-08
+    6.348199810454162e-08
+    1.824957932032937e-07
+     4.44945245802491e-07
+ 5.02e+10    
+     4.45138655056209e-07
+    1.822139705003268e-07
+    4.355999500342376e-07
+    6.351348740982953e-08
+    1.181302218363382e-07
+    4.351514289857502e-07
+     3.50976193386127e-08
+    6.349629026183344e-08
+    1.825835200543945e-07
+    4.450766967576674e-07
+ 5.03e+10    
+    4.452698361139354e-07
+    1.823020422488894e-07
+    4.357005688918008e-07
+    6.352783494198315e-08
+     1.18186493309125e-07
+    4.352522521551212e-07
+    3.507836075047008e-08
+    6.351044828575333e-08
+    1.826712969312189e-07
+    4.452083485921349e-07
+ 5.04e+10    
+    4.454012163862435e-07
+     1.82390164423097e-07
+    4.358013129258565e-07
+    6.354204775947078e-08
+    1.182427575298527e-07
+    4.353532001343673e-07
+    3.505892259527255e-08
+    6.352447208160989e-08
+    1.827591235139708e-07
+    4.453402013015333e-07
+ 5.05e+10    
+    4.455327958682588e-07
+    1.824783367043536e-07
+    4.359021820889467e-07
+    6.355612576943255e-08
+    1.182990144362197e-07
+    4.354542728745409e-07
+    3.503930512954386e-08
+    6.353836155731357e-08
+    1.828469994831118e-07
+    4.454722548824108e-07
+ 5.06e+10    
+    4.456645745560058e-07
+    1.825665587743304e-07
+    4.360031763340601e-07
+    6.357006888165898e-08
+    1.183552639665098e-07
+    4.355554703271708e-07
+    3.501950861455762e-08
+    6.355211662339443e-08
+    1.829349245193835e-07
+    4.456045093322316e-07
+ 5.07e+10    
+    4.457965524464157e-07
+    1.826548303149874e-07
+    4.361042956146388e-07
+    6.358387700860787e-08
+    1.184115060595981e-07
+    4.356567924442719e-07
+    3.499953331636002e-08
+    6.356573719301934e-08
+    1.830228983038313e-07
+     4.45736964649385e-07
+ 5.08e+10    
+    4.459287295373341e-07
+    1.827431510085973e-07
+    4.362055398845907e-07
+    6.359755006542189e-08
+    1.184677406549586e-07
+    4.357582391783544e-07
+    3.497937950579232e-08
+    6.357922318200949e-08
+    1.831109205178272e-07
+    4.458696208331918e-07
+ 5.09e+10    
+    4.460611058275305e-07
+    1.828315205377682e-07
+    4.363069090982957e-07
+    6.361108796994504e-08
+    1.185239676926708e-07
+    4.358598104824322e-07
+    3.495904745851246e-08
+    6.359257450885701e-08
+    1.831989908430929e-07
+    4.460024778839121e-07
+ 5.1e+10     
+     4.46193681316702e-07
+    1.829199385854655e-07
+    4.364084032106165e-07
+    6.362449064273921e-08
+    1.185801871134267e-07
+    4.359615063100305e-07
+    3.493853745501612e-08
+    6.360579109474172e-08
+    1.832871089617222e-07
+    4.461355358027551e-07
+ 5.11e+10    
+    4.463264560054854e-07
+    1.830084048350346e-07
+    4.365100221769055e-07
+     6.36377580071004e-08
+    1.186363988585372e-07
+    4.360633266151973e-07
+     3.49178497806572e-08
+    6.361887286354727e-08
+    1.833752745562039e-07
+    4.462687945918845e-07
+ 5.12e+10    
+    4.464594298954618e-07
+    1.830969189702232e-07
+    4.366117659530148e-07
+    6.365088998907444e-08
+    1.186926028699387e-07
+    4.361652713525086e-07
+    3.489698472566758e-08
+    6.363181974187706e-08
+    1.834634873094434e-07
+    4.464022542544255e-07
+ 5.13e+10    
+    4.465926029891635e-07
+    1.831854806752023e-07
+    4.367136344953035e-07
+    6.366388651747271e-08
+    1.187487990901998e-07
+     4.36267340477079e-07
+    3.487594258517645e-08
+    6.364463165907013e-08
+    1.835517469047854e-07
+    4.465359147944732e-07
+ 5.14e+10    
+    4.467259752900825e-07
+     1.83274089634589e-07
+    4.368156277606471e-07
+    6.367674752388723e-08
+    1.188049874625271e-07
+    4.363695339445681e-07
+    3.485472365922871e-08
+    6.365730854721614e-08
+    1.836400530260353e-07
+    4.466697762170985e-07
+ 5.15e+10    
+    4.468595468026767e-07
+    1.833627455334674e-07
+    4.369177457064459e-07
+    6.368947294270578e-08
+    1.188611679307725e-07
+    4.364718517111906e-07
+    3.483332825280314e-08
+    6.366985034117091e-08
+    1.837284053574817e-07
+    4.468038385283567e-07
+ 5.16e+10    
+    4.469933175323758e-07
+    1.834514480574101e-07
+    4.370199882906308e-07
+    6.370206271112628e-08
+     1.18917340439438e-07
+    4.365742937337218e-07
+    3.481175667582951e-08
+    6.368225697857071e-08
+    1.838168035839165e-07
+    4.469381017352919e-07
+ 5.17e+10    
+    4.471272874855886e-07
+    1.835401968924989e-07
+    4.371223554716743e-07
+    6.371451676917142e-08
+    1.189735049336832e-07
+    4.366768599695087e-07
+    3.479000924320534e-08
+    6.369452839984707e-08
+    1.839052473906576e-07
+    4.470725658459446e-07
+ 5.18e+10    
+    4.472614566697108e-07
+    1.836289917253464e-07
+     4.37224847208597e-07
+    6.372683505970242e-08
+    1.190296613593305e-07
+    4.367795503764743e-07
+    3.476808627481198e-08
+    6.370666454824061e-08
+    1.839937364635687e-07
+    4.472072308693578e-07
+ 5.19e+10    
+     4.47395825093128e-07
+    1.837178322431159e-07
+     4.37327463460975e-07
+    6.373901752843304e-08
+    1.190858096628713e-07
+    4.368823649131276e-07
+    3.474598809553001e-08
+     6.37186653698153e-08
+    1.840822704890818e-07
+    4.473420968155853e-07
+ 5.2e+10     
+     4.47530392765224e-07
+    1.838067181335425e-07
+    4.374302041889481e-07
+    6.375106412394257e-08
+    1.191419497914716e-07
+    4.369853035385709e-07
+    3.472371503525389e-08
+    6.373053081347154e-08
+    1.841708491542157e-07
+    4.474771636956943e-07
+ 5.21e+10    
+    4.476651596963874e-07
+    1.838956490849535e-07
+    4.375330693532279e-07
+    6.376297479768949e-08
+     1.19198081692978e-07
+    4.370883662125062e-07
+    3.470126742890625e-08
+     6.37422608309597e-08
+    1.842594721465985e-07
+    4.476124315217733e-07
+ 5.22e+10    
+     4.47800125898016e-07
+    1.839846247862877e-07
+    4.376360589151047e-07
+     6.37747495040238e-08
+    1.192542053159236e-07
+    4.371915528952434e-07
+    3.467864561645123e-08
+    6.375385537689298e-08
+    1.843481391544864e-07
+    4.477479003069386e-07
+ 5.23e+10    
+    4.479352913825231e-07
+    1.840736449271162e-07
+    4.377391728364542e-07
+    6.378638820019977e-08
+    1.193103206095329e-07
+    4.372948635477073e-07
+     3.46558499429074e-08
+    6.376531440876008e-08
+    1.844368498667849e-07
+    4.478835700653387e-07
+ 5.24e+10    
+    4.480706561633429e-07
+    1.841627091976613e-07
+     4.37842411079746e-07
+    6.379789084638798e-08
+    1.193664275237278e-07
+    4.373982981314445e-07
+     3.46328807583599e-08
+    6.377663788693747e-08
+    1.845256039730673e-07
+    4.480194408121608e-07
+ 5.25e+10    
+    4.482062202549365e-07
+    1.842518172888168e-07
+    4.379457736080509e-07
+    6.380925740568741e-08
+     1.19422526009133e-07
+    4.375018566086316e-07
+    3.460973841797195e-08
+    6.378782577470147e-08
+    1.846144011635961e-07
+    4.481555125636353e-07
+ 5.26e+10    
+    4.483419836727964e-07
+    1.843409688921663e-07
+    4.380492603850462e-07
+    6.382048784413677e-08
+    1.194786160170811e-07
+    4.376055389420804e-07
+    3.458642328199577e-08
+    6.379887803823992e-08
+    1.847032411293404e-07
+    4.482917853370417e-07
+ 5.27e+10    
+    4.484779464334519e-07
+    1.844301637000029e-07
+    4.381528713750246e-07
+    6.383158213072599e-08
+    1.195346974996179e-07
+    4.377093450952459e-07
+    3.456293571578278e-08
+    6.380979464666363e-08
+    1.847921235619969e-07
+    4.484282591507144e-07
+ 5.28e+10    
+    4.486141085544756e-07
+    1.845194014053483e-07
+    4.382566065428994e-07
+    6.384254023740711e-08
+    1.195907704095077e-07
+    4.378132750322331e-07
+    3.453927608979321e-08
+    6.382057557201758e-08
+    1.848810481540079e-07
+    4.485649340240458e-07
+ 5.29e+10    
+    4.487504700544857e-07
+    1.846086817019706e-07
+    4.383604658542139e-07
+    6.385336213910482e-08
+    1.196468347002381e-07
+    4.379173287178023e-07
+    3.451544477960491e-08
+     6.38312207892916e-08
+    1.849700145985803e-07
+    4.487018099774938e-07
+ 5.3e+10     
+    4.488870309531527e-07
+    1.846980042844036e-07
+    4.384644492751442e-07
+    6.386404781372701e-08
+    1.197028903260253e-07
+    4.380215061173777e-07
+    3.449144216592175e-08
+    6.384173027643097e-08
+    1.850590225897045e-07
+    4.488388870325844e-07
+ 5.31e+10    
+    4.490237912712042e-07
+    1.847873688479646e-07
+     4.38568556772509e-07
+     6.38745972421747e-08
+    1.197589372418184e-07
+    4.381258071970516e-07
+    3.446726863458112e-08
+    6.385210401434657e-08
+     1.85148071822172e-07
+    4.489761652119178e-07
+ 5.32e+10    
+    4.491607510304277e-07
+    1.848767750887719e-07
+    4.386727883137741e-07
+    6.388501040835189e-08
+    1.198149754033052e-07
+    4.382302319235933e-07
+    3.444292457656085e-08
+    6.386234198692491e-08
+    1.852371619915949e-07
+     4.49113644539172e-07
+ 5.33e+10    
+    4.492979102536772e-07
+     1.84966222703764e-07
+    4.387771438670611e-07
+    6.389528729917475e-08
+    1.198710047669156e-07
+    4.383347802644521e-07
+    3.441841038798558e-08
+    6.387244418103753e-08
+    1.853262927944223e-07
+    4.492513250391074e-07
+ 5.34e+10    
+    4.494352689648762e-07
+    1.850557113907161e-07
+    4.388816234011508e-07
+    6.390542790458112e-08
+    1.199270252898275e-07
+    4.384394521877668e-07
+     3.43937264701323e-08
+    6.388241058655055e-08
+    1.854154639279594e-07
+    4.493892067375722e-07
+ 5.35e+10    
+    4.495728271890209e-07
+    1.851452408482574e-07
+    4.389862268854905e-07
+     6.39154322175391e-08
+    1.199830369299706e-07
+    4.385442476623698e-07
+     3.43688732294353e-08
+    6.389224119633346e-08
+    1.855046750903841e-07
+    4.495272896615045e-07
+ 5.36e+10    
+    4.497105849521884e-07
+    1.852348107758894e-07
+    4.390909542902014e-07
+     6.39253002340556e-08
+    1.200390396460311e-07
+    4.386491666577932e-07
+    3.434385107749053e-08
+    6.390193600626796e-08
+    1.855939259807648e-07
+    4.496655738389383e-07
+ 5.37e+10    
+    4.498485422815341e-07
+    1.853244208740015e-07
+    4.391958055860824e-07
+    6.393503195318452e-08
+    1.200950333974558e-07
+    4.387542091442743e-07
+    3.431866043105913e-08
+    6.391149501525617e-08
+    1.856832162990773e-07
+    4.498040592990057e-07
+ 5.38e+10    
+    4.499866992053021e-07
+    1.854140708438887e-07
+    4.393007807446182e-07
+     6.39446273770349e-08
+    1.201510181444569e-07
+    4.388593750927633e-07
+    3.429330171207043e-08
+    6.392091822522897e-08
+    1.857725457462219e-07
+    4.499427460719426e-07
+ 5.39e+10    
+    4.501250557528241e-07
+    1.855037603877678e-07
+    4.394058797379826e-07
+    6.395408651077818e-08
+    1.202069938480158e-07
+    4.389646644749266e-07
+    3.426777534762428e-08
+    6.393020564115367e-08
+    1.858619140240399e-07
+    4.500816341890911e-07
+ 5.4e+10     
+    4.502636119545262e-07
+     1.85593489208794e-07
+    4.395111025390468e-07
+    6.396340936265582e-08
+    1.202629604698874e-07
+    4.390700772631542e-07
+    3.424208176999261e-08
+    6.393935727104144e-08
+    1.859513208353301e-07
+    4.502207236829029e-07
+ 5.41e+10    
+    4.504023678419298e-07
+    1.856832570110766e-07
+    4.396164491213822e-07
+    6.397259594398612e-08
+    1.203189179726039e-07
+    4.391756134305635e-07
+    3.421622141662044e-08
+    6.394837312595455e-08
+    1.860407658838651e-07
+    4.503600145869434e-07
+ 5.42e+10    
+    4.505413234476563e-07
+     1.85773063499695e-07
+    4.397219194592685e-07
+    6.398164626917097e-08
+    1.203748663194792e-07
+    4.392812729510055e-07
+    3.419019473012619e-08
+    6.395725322001339e-08
+    1.861302488744075e-07
+    4.504995069358959e-07
+ 5.43e+10    
+    4.506804788054312e-07
+     1.85862908380715e-07
+    4.398275135276978e-07
+    6.399056035570235e-08
+    1.204308054746124e-07
+    4.393870557990715e-07
+    3.416400215830121e-08
+    6.396599757040278e-08
+    1.862197695127253e-07
+    4.506392007655618e-07
+ 5.44e+10    
+    4.508198339500854e-07
+    1.859527913612037e-07
+    4.399332313023806e-07
+    6.399933822416817e-08
+    1.204867354028919e-07
+    4.394929619500952e-07
+     3.41376441541089e-08
+    6.397460619737854e-08
+     1.86309327505608e-07
+     4.50779096112867e-07
+ 5.45e+10    
+     4.50959388917558e-07
+    1.860427121492446e-07
+    4.400390727597491e-07
+    6.400797989825835e-08
+    1.205426560699984e-07
+    4.395989913801605e-07
+    3.411112117568286e-08
+    6.398307912427332e-08
+    1.863989225608816e-07
+    4.509191930158631e-07
+ 5.46e+10    
+    4.510991437449022e-07
+    1.861326704539534e-07
+    4.401450378769652e-07
+    6.401648540477021e-08
+    1.205985674424097e-07
+    4.397051440661058e-07
+    3.408443368632464e-08
+    6.399141637750233e-08
+    1.864885543874242e-07
+    4.510594915137316e-07
+ 5.47e+10    
+     4.51239098470285e-07
+    1.862226659854923e-07
+    4.402511266319236e-07
+    6.402485477361355e-08
+    1.206544694874032e-07
+    4.398114199855273e-07
+    3.405758215450059e-08
+     6.39996179865687e-08
+    1.865782226951805e-07
+    4.511999916467843e-07
+ 5.48e+10    
+    4.513792531329904e-07
+    1.863126984550844e-07
+     4.40357339003257e-07
+    6.403308803781576e-08
+      1.2071036217306e-07
+    4.399178191167874e-07
+    3.403056705383827e-08
+    6.400768398406869e-08
+    1.866679271951769e-07
+    4.513406934564688e-07
+ 5.49e+10    
+    4.515196077734239e-07
+    1.864027675750297e-07
+    4.404636749703424e-07
+    6.404118523352628e-08
+    1.207662454682678e-07
+    4.400243414390151e-07
+    3.400338886312203e-08
+    6.401561440569637e-08
+    1.867576675995361e-07
+     4.51481596985369e-07
+ 5.5e+10     
+    4.516601624331115e-07
+    1.864928730587167e-07
+    4.405701345133028e-07
+    6.404914640002075e-08
+    1.208221193427245e-07
+     4.40130986932114e-07
+    3.397604806628796e-08
+    6.402340929024803e-08
+     1.86847443621491e-07
+    4.516227022772083e-07
+ 5.51e+10    
+    4.518009171547061e-07
+     1.86583014620639e-07
+    4.406767176130157e-07
+    6.405697157970536e-08
+    1.208779837669414e-07
+    4.402377555767654e-07
+    3.394854515241825e-08
+     6.40310686796267e-08
+     1.86937254975399e-07
+    4.517640093768523e-07
+ 5.52e+10    
+    4.519418719819863e-07
+    1.866731919764071e-07
+    4.407834242511149e-07
+    6.406466081812032e-08
+    1.209338387122464e-07
+    4.403446473544328e-07
+    3.392088061573484e-08
+    6.403859261884582e-08
+    1.870271013767568e-07
+    4.519055183303106e-07
+ 5.53e+10    
+    4.520830269598609e-07
+    1.867634048427637e-07
+    4.408902544099964e-07
+    6.407221416394329e-08
+    1.209896841507869e-07
+    4.404516622473677e-07
+     3.38930549555923e-08
+    6.404598115603276e-08
+    1.871169825422121e-07
+    4.520472291847384e-07
+ 5.54e+10    
+    4.522243821343697e-07
+    1.868536529375953e-07
+    4.409972080728214e-07
+    6.407963166899243e-08
+    1.210455200555326e-07
+    4.405588002386111e-07
+    3.386506867647028e-08
+    6.405323434243237e-08
+     1.87206898189579e-07
+    4.521891419884397e-07
+ 5.55e+10    
+    4.523659375526849e-07
+    1.869439359799472e-07
+    4.411042852235229e-07
+    6.408691338822936e-08
+     1.21101346400279e-07
+    4.406660613120003e-07
+    3.383692228796509e-08
+    6.406035223240996e-08
+    1.872968480378503e-07
+    4.523312567908682e-07
+ 5.56e+10    
+     4.52507693263115e-07
+    1.870342536900346e-07
+    4.412114858468068e-07
+    6.409405937976155e-08
+    1.211571631596496e-07
+    4.407734454521729e-07
+    3.380861630478075e-08
+    6.406733488345384e-08
+    1.873868318072109e-07
+    4.524735736426298e-07
+ 5.57e+10    
+    4.526496493151048e-07
+    1.871246057892573e-07
+     4.41318809928161e-07
+    6.410106970484454e-08
+    1.212129703090988e-07
+    4.408809526445679e-07
+    3.378015124671932e-08
+    6.407418235617804e-08
+    1.874768492190503e-07
+    4.526160925954844e-07
+ 5.58e+10    
+    4.527918057592377e-07
+    1.872149920002101e-07
+    4.414262574538527e-07
+    6.410794442788398e-08
+    1.212687678249148e-07
+    4.409885828754338e-07
+     3.37515276386705e-08
+    6.408089471432413e-08
+    1.875668999959752e-07
+    4.527588137023457e-07
+ 5.59e+10    
+    4.529341626472355e-07
+    1.873054120466971e-07
+    4.415338284109387e-07
+    6.411468361643712e-08
+     1.21324555684222e-07
+    4.410963361318296e-07
+    3.372274601060084e-08
+    6.408747202476341e-08
+    1.876569838618226e-07
+    4.529017370172859e-07
+ 5.6e+10     
+     4.53076720031964e-07
+    1.873958656537425e-07
+    4.416415227872656e-07
+     6.41212873412143e-08
+    1.213803338649835e-07
+    4.412042124016305e-07
+    3.369380689754194e-08
+    6.409391435749818e-08
+     1.87747100541671e-07
+    4.530448625955342e-07
+ 5.61e+10    
+    4.532194779674291e-07
+    1.874863525476027e-07
+    4.417493405714751e-07
+    6.412775567607973e-08
+    1.214361023460033e-07
+    4.413122116735287e-07
+    3.366471083957829e-08
+    6.410022178566319e-08
+    1.878372497618533e-07
+    4.531881904934804e-07
+ 5.62e+10    
+    4.533624365087822e-07
+    1.875768724557787e-07
+    4.418572817530072e-07
+    6.413408869805265e-08
+    1.214918611069293e-07
+    4.414203339370412e-07
+    3.363545838183432e-08
+    6.410639438552663e-08
+    1.879274312499677e-07
+    4.533317207686735e-07
+ 5.63e+10    
+    4.535055957123199e-07
+    1.876674251070269e-07
+    4.419653463221042e-07
+    6.414028648730745e-08
+    1.215476101282548e-07
+    4.415285791825094e-07
+    3.360605007446079e-08
+    6.411243223649064e-08
+      1.8801764473489e-07
+    4.534754534798256e-07
+ 5.64e+10    
+    4.536489556354831e-07
+    1.877580102313704e-07
+    4.420735342698134e-07
+    6.414634912717397e-08
+     1.21603349391321e-07
+     4.41636947401105e-07
+    3.357648647262061e-08
+    6.411833542109192e-08
+    1.881078899467846e-07
+    4.536193886868114e-07
+ 5.65e+10    
+    4.537925163368614e-07
+      1.8784862756011e-07
+    4.421818455879927e-07
+    6.415227670413744e-08
+    1.216590788783192e-07
+    4.417454385848331e-07
+    3.354676813647396e-08
+    6.412410402500185e-08
+    1.881981666171156e-07
+    4.537635264506697e-07
+ 5.66e+10    
+    4.539362778761917e-07
+    1.879392768258362e-07
+     4.42290280269312e-07
+    6.415806930783809e-08
+    1.217147985722929e-07
+    4.418540527265341e-07
+    3.351689563116279e-08
+    6.412973813702612e-08
+    1.882884744786576e-07
+    4.539078668336028e-07
+ 5.67e+10    
+    4.540802403143603e-07
+    1.880299577624378e-07
+    4.423988383072563e-07
+    6.416372703107035e-08
+    1.217705084571392e-07
+     4.41962789819888e-07
+    3.348686952679467e-08
+    6.413523784910446e-08
+    1.883788132655069e-07
+    4.540524098989804e-07
+ 5.68e+10    
+    4.542244037134013e-07
+    1.881206701051138e-07
+    4.425075196961311e-07
+    6.416924996978191e-08
+    1.218262085176116e-07
+    4.420716498594179e-07
+    3.345669039842595e-08
+    6.414060325630986e-08
+    1.884691827130914e-07
+    4.541971557113363e-07
+ 5.69e+10    
+    4.543687681365004e-07
+    1.882114135903836e-07
+    4.426163244310638e-07
+    6.417463822307269e-08
+    1.218818987393208e-07
+     4.42180632840493e-07
+     3.34263588260445e-08
+    6.414583445684765e-08
+    1.885595825581817e-07
+    4.543421043363728e-07
+ 5.7e+10     
+    4.545133336479918e-07
+    1.883021879560962e-07
+    4.427252525080067e-07
+    6.417989189319292e-08
+    1.219375791087371e-07
+    4.422897387593293e-07
+    3.339587539455142e-08
+    6.415093155205389e-08
+    1.886500125388998e-07
+    4.544872558409575e-07
+ 5.71e+10    
+    4.546581003133626e-07
+    1.883929929414409e-07
+    4.428343039237419e-07
+    6.418501108554173e-08
+    1.219932496131918e-07
+     4.42398967612997e-07
+    3.336524069374258e-08
+    6.415589464639428e-08
+    1.887404723947308e-07
+    4.546326102931276e-07
+ 5.72e+10    
+    4.548030681992496e-07
+    1.884838282869563e-07
+    4.429434786758822e-07
+     6.41899959086648e-08
+    1.220489102408789e-07
+    4.425083193994185e-07
+    3.333445531828914e-08
+    6.416072384746181e-08
+    1.888309618665309e-07
+    4.547781677620862e-07
+ 5.73e+10    
+    4.549482373734419e-07
+    1.885746937345399e-07
+    4.430527767628746e-07
+    6.419484647425198e-08
+    1.221045609808562e-07
+    4.426177941173745e-07
+    3.330351986771772e-08
+    6.416541926597499e-08
+    1.889214806965379e-07
+    4.549239283182065e-07
+ 5.74e+10    
+    4.550936079048795e-07
+    1.886655890274574e-07
+    4.431621981840035e-07
+    6.419956289713475e-08
+    1.221602018230473e-07
+    4.427273917665049e-07
+    3.327243494638971e-08
+    6.416998101577519e-08
+      1.8901202862838e-07
+    4.550698920330279e-07
+ 5.75e+10    
+    4.552391798636542e-07
+    1.887565139103516e-07
+    4.432717429393933e-07
+    6.420414529528334e-08
+    1.222158327582426e-07
+    4.428371123473124e-07
+    3.324120116348028e-08
+    6.417440921382421e-08
+     1.89102605407085e-07
+      4.5521605897926e-07
+ 5.76e+10    
+    4.553849533210094e-07
+    1.888474681292514e-07
+    4.433814110300107e-07
+    6.420859378980333e-08
+    1.222714537781006e-07
+    4.429469558611652e-07
+     3.32098191329564e-08
+    6.417870398020102e-08
+    1.891932107790894e-07
+    4.553624292307798e-07
+ 5.77e+10    
+    4.555309283493402e-07
+    1.889384514315799e-07
+    4.434912024576672e-07
+    6.421290850493228e-08
+    1.223270648751491e-07
+    4.430569223102973e-07
+     3.31782894735545e-08
+     6.41828654380987e-08
+    1.892838444922462e-07
+    4.555090028626327e-07
+ 5.78e+10    
+    4.556771050221925e-07
+    1.890294635661633e-07
+    4.436011172250223e-07
+    6.421708956803598e-08
+    1.223826660427863e-07
+    4.431670116978143e-07
+    3.314661280875745e-08
+    6.418689371382095e-08
+    1.893745062958341e-07
+    4.556557799510316e-07
+ 5.79e+10    
+    4.558234834142641e-07
+     1.89120504283239e-07
+     4.43711155335585e-07
+    6.422113710960439e-08
+    1.224382572752817e-07
+    4.432772240276912e-07
+    3.311478976677096e-08
+    6.419078893677821e-08
+    1.894651959405658e-07
+    4.558027605733583e-07
+ 5.8e+10     
+    4.559700636014029e-07
+    1.892115733344632e-07
+    4.438213167937161e-07
+    6.422505126324747e-08
+    1.224938385677777e-07
+    4.433875593047812e-07
+    3.308282098049924e-08
+    6.419455123948369e-08
+    1.895559131785954e-07
+    4.559499448081612e-07
+ 5.81e+10    
+    4.561168456606066e-07
+    1.893026704729191e-07
+    4.439316016046326e-07
+    6.422883216569031e-08
+    1.225494099162899e-07
+    4.434980175348103e-07
+    3.305070708752029e-08
+    6.419818075754897e-08
+    1.896466577635268e-07
+    4.560973327351557e-07
+ 5.82e+10    
+    4.562638296700252e-07
+    1.893937954531251e-07
+    4.440420097744072e-07
+    6.423247995676872e-08
+    1.226049713177078e-07
+    4.436085987243848e-07
+    3.301844873006043e-08
+     6.42016776296795e-08
+    1.897374294504209e-07
+    4.562449244352236e-07
+ 5.83e+10    
+    4.564110157089547e-07
+    1.894849480310402e-07
+    4.441525413099699e-07
+    6.423599477942372e-08
+    1.226605227697961e-07
+     4.43719302880991e-07
+     3.29860465549682e-08
+    6.420504199766963e-08
+    1.898282279958033e-07
+    4.563927199904133e-07
+ 5.84e+10    
+    4.565584038578409e-07
+    1.895761279640733e-07
+    4.442631962191143e-07
+    6.423937677969635e-08
+    1.227160642711949e-07
+    4.438301300129976e-07
+    3.295350121368786e-08
+    6.420827400639764e-08
+    1.899190531576714e-07
+    4.565407194839379e-07
+ 5.85e+10    
+    4.567059941982792e-07
+    1.896673350110897e-07
+    4.443739745104955e-07
+    6.424262610672218e-08
+    1.227715958214208e-07
+    4.439410801296578e-07
+    3.292081336223212e-08
+    6.421137380382023e-08
+    1.900099046955018e-07
+    4.566889230001753e-07
+ 5.86e+10    
+    4.568537868130103e-07
+    1.897585689324168e-07
+    4.444848761936331e-07
+    6.424574291272523e-08
+    1.228271174208669e-07
+    4.440521532411102e-07
+    3.288798366115442e-08
+    6.421434154096703e-08
+    1.901007823702564e-07
+    4.568373306246671e-07
+ 5.87e+10    
+     4.57001781785922e-07
+    1.898498294898523e-07
+    4.445959012789134e-07
+    6.424872735301171e-08
+    1.228826290708037e-07
+    4.441633493583822e-07
+     3.28550127755205e-08
+    6.421717737193438e-08
+    1.901916859443897e-07
+    4.569859424441181e-07
+ 5.88e+10    
+    4.571499792020464e-07
+    1.899411164466693e-07
+    4.447070497775917e-07
+    6.425157958596395e-08
+     1.22938130773379e-07
+    4.442746684933903e-07
+     3.28219013748795e-08
+    6.421988145387954e-08
+    1.902826151818548e-07
+    4.571347585463942e-07
+ 5.89e+10    
+    4.572983791475616e-07
+    1.900324295676233e-07
+    4.448183217017922e-07
+    6.425429977303337e-08
+     1.22993622531619e-07
+    4.443861106589402e-07
+    3.278865013323452e-08
+    6.422245394701409e-08
+    1.903735698481102e-07
+    4.572837790205234e-07
+ 5.9e+10     
+    4.574469817097876e-07
+    1.901237686189581e-07
+    4.449297170645113e-07
+    6.425688807873388e-08
+    1.230491043494278e-07
+     4.44497675868734e-07
+    3.275525972901248e-08
+    6.422489501459725e-08
+    1.904645497101253e-07
+    4.574330039566934e-07
+ 5.91e+10    
+    4.575957869771874e-07
+    1.902151333684118e-07
+    4.450412358796196e-07
+    6.425934467063439e-08
+    1.231045762315877e-07
+    4.446093641373631e-07
+    3.272173084503351e-08
+     6.42272048229289e-08
+    1.905555545363862e-07
+    4.575824334462497e-07
+ 5.92e+10    
+    4.577447950393644e-07
+    1.903065235852219e-07
+    4.451528781618606e-07
+    6.426166971935156e-08
+      1.2316003818376e-07
+    4.447211754803179e-07
+     3.26880641684798e-08
+    6.422938354134253e-08
+    1.906465840969019e-07
+     4.57732067581696e-07
+ 5.93e+10    
+    4.578940059870623e-07
+    1.903979390401311e-07
+    4.452646439268548e-07
+    6.426386339854202e-08
+     1.23215490212484e-07
+    4.448331099139832e-07
+    3.265426039086389e-08
+    6.423143134219769e-08
+    1.907376381632096e-07
+    4.578819064566923e-07
+ 5.94e+10    
+    4.580434199121631e-07
+    1.904893795053933e-07
+    4.453765331910995e-07
+    6.426592588489455e-08
+    1.232709323251779e-07
+    4.449451674556428e-07
+    3.262032020799632e-08
+    6.423334840087239e-08
+    1.908287165083797e-07
+    4.580319501660545e-07
+ 5.95e+10    
+    4.581930369076846e-07
+    1.905808447547771e-07
+    4.454885459719722e-07
+    6.426785735812169e-08
+    1.233263645301382e-07
+    4.450573481234787e-07
+    3.258624431995289e-08
+    6.423513489575508e-08
+    1.909198189070211e-07
+    4.581821988057496e-07
+ 5.96e+10    
+    4.583428570677824e-07
+    1.906723345635723e-07
+    4.456006822877287e-07
+    6.426965800095152e-08
+    1.233817868365394e-07
+    4.451696519365734e-07
+     3.25520334310412e-08
+    6.423679100823646e-08
+    1.910109451352864e-07
+    4.583326524728985e-07
+ 5.97e+10    
+     4.58492880487744e-07
+    1.907638487085939e-07
+    4.457129421575065e-07
+    6.427132799911891e-08
+    1.234371992544344e-07
+    4.452820789149109e-07
+    3.251768824976694e-08
+    6.423831692270117e-08
+    1.911020949708759e-07
+    4.584833112657733e-07
+ 5.98e+10    
+    4.586431072639914e-07
+    1.908553869681865e-07
+    4.458253256013256e-07
+    6.427286754135647e-08
+    1.234926017947536e-07
+    4.453946290793766e-07
+    3.248320948879929e-08
+    6.423971282651905e-08
+    1.911932681930428e-07
+    4.586341752837928e-07
+ 5.99e+10    
+    4.587935374940745e-07
+    1.909469491222292e-07
+    4.459378326400885e-07
+    6.427427681938553e-08
+    1.235479944693048e-07
+    4.455073024517593e-07
+    3.244859786493609e-08
+    6.424097891003616e-08
+    1.912844645825976e-07
+    4.587852446275248e-07
+ 6e+10       
+    4.589441712766752e-07
+    1.910385349521393e-07
+    4.460504632955824e-07
+    6.427555602790668e-08
+    1.236033772907728e-07
+    4.456200990547512e-07
+    3.241385409906838e-08
+    6.424211536656568e-08
+    1.913756839219115e-07
+     4.58936519398682e-07
+ 6.01e+10    
+    4.590950087116014e-07
+    1.911301442408766e-07
+    4.461632175904793e-07
+    6.427670536459014e-08
+    1.236587502727188e-07
+    4.457330189119497e-07
+    3.237897891614441e-08
+    6.424312239237864e-08
+    1.914669259949213e-07
+    4.590879997001218e-07
+ 6.02e+10    
+    4.592460498997863e-07
+    1.912217767729471e-07
+    4.462760955483364e-07
+    6.427772503006592e-08
+    1.237141134295798e-07
+    4.458460620478569e-07
+    3.234397304513318e-08
+    6.424400018669414e-08
+    1.915581905871328e-07
+    4.592396856358429e-07
+ 6.03e+10    
+    4.593972949432887e-07
+     1.91313432334407e-07
+    4.463890971935996e-07
+     6.42786152279136e-08
+    1.237694667766681e-07
+    4.459592284878818e-07
+     3.23088372189875e-08
+    6.424474895166947e-08
+    1.916494774856242e-07
+    4.593915773109841e-07
+ 6.04e+10    
+    4.595487439452863e-07
+    1.914051107128652e-07
+    4.465022225515991e-07
+    6.427937616465208e-08
+    1.238248103301708e-07
+    4.460725182583394e-07
+    3.227357217460643e-08
+    6.424536889239013e-08
+    1.917407864790501e-07
+    4.595436748318225e-07
+ 6.05e+10    
+    4.597003970100787e-07
+    1.914968116974881e-07
+    4.466154716485552e-07
+    6.428000804972891e-08
+     1.23880144107148e-07
+    4.461859313864515e-07
+     3.22381786527975e-08
+    6.424586021685945e-08
+    1.918321173576446e-07
+    4.596959783057721e-07
+ 6.06e+10    
+    4.598522542430829e-07
+    1.915885350790014e-07
+    4.467288445115768e-07
+    6.428051109550963e-08
+     1.23935468125534e-07
+    4.462994679003478e-07
+    3.220265739823809e-08
+    6.424622313598809e-08
+    1.919234699132238e-07
+    4.598484878413805e-07
+ 6.07e+10    
+    4.600043157508318e-07
+     1.91680280649694e-07
+    4.468423411686602e-07
+    6.428088551726665e-08
+     1.23990782404134e-07
+    4.464131278290659e-07
+    3.216700915943659e-08
+    6.424645786358312e-08
+    1.920148439391898e-07
+    4.600012035483274e-07
+ 6.08e+10    
+    4.601565816409702e-07
+    1.917720482034197e-07
+    4.469559616486934e-07
+    6.428113153316782e-08
+    1.240460869626251e-07
+    4.465269112025525e-07
+    3.213123468869307e-08
+    6.424656461633716e-08
+    1.921062392305325e-07
+    4.601541255374229e-07
+ 6.09e+10    
+    4.603090520222575e-07
+    1.918638375356013e-07
+    4.470697059814524e-07
+     6.42812493642654e-08
+    1.241013818215543e-07
+    4.466408180516614e-07
+    3.209533474205934e-08
+    6.424654361381712e-08
+    1.921976555838329e-07
+    4.603072539206047e-07
+ 6.1e+10     
+    4.604617270045595e-07
+    1.919556484432318e-07
+    4.471835741976045e-07
+    6.428123923448384e-08
+    1.241566670023375e-07
+     4.46754848408157e-07
+    3.205931007929863e-08
+    6.424639507845272e-08
+     1.92289092797265e-07
+    4.604605888109362e-07
+ 6.11e+10    
+    4.606146066988503e-07
+    1.920474807248771e-07
+    4.472975663287066e-07
+    6.428110137060822e-08
+    1.242119425272584e-07
+    4.468690023047098e-07
+    3.202316146384491e-08
+    6.424611923552472e-08
+    1.923805506705984e-07
+    4.606141303226038e-07
+ 6.12e+10    
+    4.607676912172084e-07
+    1.921393341806786e-07
+    4.474116824072084e-07
+    6.428083600227193e-08
+    1.242672084194681e-07
+    4.469832797749033e-07
+    3.198688966276157e-08
+    6.424571631315333e-08
+       1.924720290052e-07
+    4.607678785709158e-07
+ 6.13e+10    
+    4.609209806728151e-07
+    1.922312086123541e-07
+    4.475259224664482e-07
+    6.428044336194449e-08
+    1.243224647029823e-07
+    4.470976808532275e-07
+    3.195049544669984e-08
+    6.424518654228582e-08
+    1.925635276040365e-07
+    4.609218336722978e-07
+ 6.14e+10    
+    4.610744751799497e-07
+    1.923231038232006e-07
+    4.476402865406561e-07
+    6.427992368491871e-08
+    1.243777114026813e-07
+    4.472122055750817e-07
+    3.191397958985659e-08
+    6.424453015668419e-08
+    1.926550462716751e-07
+    4.610759957442922e-07
+ 6.15e+10    
+    4.612281748539917e-07
+    1.924150196180958e-07
+    4.477547746649547e-07
+     6.42792772092982e-08
+     1.24432948544308e-07
+    4.473268539767758e-07
+    3.187734286993198e-08
+    6.424374739291299e-08
+    1.927465848142868e-07
+     4.61230364905556e-07
+ 6.16e+10    
+    4.613820798114141e-07
+    1.925069558034987e-07
+    4.478693868753556e-07
+    6.427850417598428e-08
+    1.244881761544668e-07
+    4.474416260955273e-07
+    3.184058606808634e-08
+    6.424283849032617e-08
+    1.928381430396462e-07
+    4.613849412758562e-07
+ 6.17e+10    
+     4.61536190169782e-07
+     1.92598912187452e-07
+    4.479841232087631e-07
+    6.427760482866266e-08
+    1.245433942606215e-07
+    4.475565219694629e-07
+    3.180370996889683e-08
+    6.424180369105445e-08
+    1.929297207571332e-07
+    4.615397249760693e-07
+ 6.18e+10    
+    4.616905060477511e-07
+    1.926908885795825e-07
+    4.480989837029714e-07
+    6.427657941379024e-08
+    1.245986028910945e-07
+     4.47671541637618e-07
+    3.176671536031377e-08
+    6.424064323999188e-08
+    1.930213177777346e-07
+    4.616947161281779e-07
+ 6.19e+10    
+     4.61845027565064e-07
+    1.927828847911027e-07
+    4.482139683966654e-07
+    6.427542818058147e-08
+    1.246538020750646e-07
+    4.477866851399366e-07
+    3.172960303361636e-08
+    6.423935738478283e-08
+    1.931129339140448e-07
+    4.618499148552674e-07
+ 6.2e+10     
+    4.619997548425483e-07
+     1.92874900634811e-07
+    4.483290773294215e-07
+    6.427415138099442e-08
+    1.247089918425656e-07
+    4.479019525172698e-07
+    3.169237378336812e-08
+    6.423794637580807e-08
+     1.93204568980266e-07
+    4.620053212815245e-07
+ 6.21e+10    
+    4.621546880021135e-07
+    1.929669359250932e-07
+    4.484443105417054e-07
+     6.42727492697169e-08
+    1.247641722244845e-07
+     4.48017343811377e-07
+    3.165502840737193e-08
+    6.423641046617136e-08
+    1.932962227922098e-07
+    4.621609355322349e-07
+ 6.22e+10    
+    4.623098271667479e-07
+    1.930589904779217e-07
+    4.485596680748735e-07
+    6.427122210415229e-08
+    1.248193432525597e-07
+    4.481328590649247e-07
+    3.161756770662473e-08
+     6.42347499116853e-08
+    1.933878951672972e-07
+    4.623167577337786e-07
+ 6.23e+10    
+    4.624651724605169e-07
+    1.931510641108581e-07
+    4.486751499711715e-07
+    6.426957014440508e-08
+    1.248745049593791e-07
+    4.482484983214862e-07
+    3.157999248527168e-08
+    6.423296497085719e-08
+    1.934795859245587e-07
+    4.624727880136292e-07
+ 6.24e+10    
+    4.626207240085594e-07
+    1.932431566430508e-07
+     4.48790756273734e-07
+     6.42677936532664e-08
+    1.249296573783783e-07
+    4.483642616255403e-07
+    3.154230355056017e-08
+    6.423105590487482e-08
+     1.93571294884635e-07
+    4.626290265003488e-07
+ 6.25e+10    
+    4.627764819370851e-07
+    1.933352678952373e-07
+    4.489064870265843e-07
+    6.426589289619905e-08
+    1.249848005438386e-07
+    4.484801490224721e-07
+     3.15045017127933e-08
+    6.422902297759179e-08
+    1.936630218697764e-07
+    4.627854733235881e-07
+ 6.26e+10    
+    4.629324463733714e-07
+    1.934273976897426e-07
+    4.490223422746343e-07
+    6.426386814132268e-08
+    1.250399344908846e-07
+    4.485961605585698e-07
+    3.146658778528306e-08
+    6.422686645551296e-08
+    1.937547667038431e-07
+    4.629421286140813e-07
+ 6.27e+10    
+    4.630886174457629e-07
+    1.935195458504803e-07
+    4.491383220636829e-07
+    6.426171965939895e-08
+    1.250950592554831e-07
+    4.487122962810295e-07
+    3.142856258430321e-08
+    6.422458660777937e-08
+    1.938465292123052e-07
+    4.630989925036437e-07
+ 6.28e+10    
+    4.632449952836632e-07
+     1.93611712202951e-07
+    4.492544264404162e-07
+    6.425944772381551e-08
+      1.2515017487444e-07
+    4.488285562379467e-07
+     3.13904269290417e-08
+    6.422218370615343e-08
+    1.939383092222419e-07
+    4.632560651251698e-07
+ 6.29e+10    
+    4.634015800175381e-07
+    1.937038965742429e-07
+    4.493706554524069e-07
+    6.425705261057117e-08
+    1.252052813853982e-07
+    4.489449404783217e-07
+    3.135218164155294e-08
+    6.421965802500337e-08
+    1.940301065623406e-07
+    4.634133466126288e-07
+ 6.3e+10     
+    4.635583717789077e-07
+    1.937960987930305e-07
+    4.494870091481117e-07
+    6.425453459825987e-08
+    1.252603788268362e-07
+    4.490614490520565e-07
+    3.131382754670944e-08
+    6.421700984128787e-08
+    1.941219210628968e-07
+    4.635708371010622e-07
+ 6.31e+10    
+    4.637153707003479e-07
+    1.938883186895741e-07
+    4.496034875768744e-07
+    6.425189396805496e-08
+    1.253154672380647e-07
+    4.491780820099536e-07
+    3.127536547215357e-08
+    6.421423943454073e-08
+    1.942137525558134e-07
+     4.63728536726582e-07
+ 6.32e+10    
+    4.638725769154826e-07
+    1.939805560957193e-07
+    4.497200907889207e-07
+    6.424913100369315e-08
+    1.253705466592252e-07
+    4.492948394037153e-07
+    3.123679624824853e-08
+    6.421134708685462e-08
+    1.943056008745989e-07
+    4.638864456263654e-07
+ 6.33e+10    
+    4.640299905589848e-07
+    1.940728108448947e-07
+    4.498368188353607e-07
+    6.424624599145823e-08
+    1.254256171312868e-07
+    4.494117212859432e-07
+    3.119812070802935e-08
+    6.420833308286542e-08
+    1.943974658543671e-07
+    4.640445639386535e-07
+ 6.34e+10    
+    4.641876117665707e-07
+    1.941650827721122e-07
+    4.499536717681858e-07
+    6.424323922016491e-08
+    1.254806786960446e-07
+    4.495287277101374e-07
+     3.11593396871535e-08
+     6.42051977097361e-08
+    1.944893473318354e-07
+    4.642028918027482e-07
+ 6.35e+10    
+    4.643454406749978e-07
+     1.94257371713965e-07
+    4.500706496402687e-07
+    6.424011098114214e-08
+    1.255357313961164e-07
+    4.496458587306947e-07
+    3.112045402385113e-08
+    6.420194125714034e-08
+    1.945812451453237e-07
+    4.643614293590075e-07
+ 6.36e+10    
+    4.645034774220627e-07
+    1.943496775086259e-07
+     4.50187752505362e-07
+    6.423686156821632e-08
+    1.255907752749405e-07
+    4.497631144029067e-07
+    3.108146455887508e-08
+    6.419856401724595e-08
+    1.946731591347526e-07
+    4.645201767488445e-07
+ 6.37e+10    
+    4.646617221465955e-07
+    1.944419999958469e-07
+    4.503049804180991e-07
+    6.423349127769479e-08
+    1.256458103767734e-07
+    4.498804947829607e-07
+    3.104237213545071e-08
+    6.419506628469852e-08
+    1.947650891416421e-07
+    4.646791341147222e-07
+ 6.38e+10    
+    4.648201749884601e-07
+    1.945343390169559e-07
+    4.504223334339891e-07
+    6.423000040834842e-08
+    1.257008367466862e-07
+    4.499979999279367e-07
+    3.100317759922529e-08
+    6.419144835660434e-08
+    1.948570350091091e-07
+    4.648383016001519e-07
+ 6.39e+10    
+    4.649788360885463e-07
+     1.94626694414856e-07
+    4.505398116094191e-07
+    6.422638926139477e-08
+    1.257558544305634e-07
+    4.501156298958083e-07
+    3.096388179821727e-08
+    6.418771053251384e-08
+    1.949489965818669e-07
+    4.649976793496901e-07
+ 6.4e+10     
+    4.651377055887725e-07
+    1.947190660340236e-07
+    4.506574150016522e-07
+     6.42226581404806e-08
+    1.258108634750987e-07
+    4.502333847454379e-07
+    3.092448558276515e-08
+      6.4183853114404e-08
+    1.950409737062214e-07
+    4.651572675089328e-07
+ 6.41e+10    
+    4.652967836320767e-07
+    1.948114537205054e-07
+    4.507751436688254e-07
+    6.421880735166434e-08
+    1.258658639277929e-07
+    4.503512645365792e-07
+    3.088498980547633e-08
+    6.417987640666157e-08
+    1.951329662300706e-07
+    4.653170662245164e-07
+ 6.42e+10    
+    4.654560703624175e-07
+    1.949038573219173e-07
+    4.508929976699494e-07
+    6.421483720339871e-08
+     1.25920855836951e-07
+    4.504692693298734e-07
+    3.084539532117547e-08
+    6.417578071606549e-08
+    1.952249740029013e-07
+    4.654770756441106e-07
+ 6.43e+10    
+    4.656155659247693e-07
+    1.949962766874418e-07
+    4.510109770649061e-07
+    6.421074800651279e-08
+    1.259758392516794e-07
+    4.505873991868482e-07
+     3.08057029868528e-08
+    6.417156635176912e-08
+    1.953169968757867e-07
+     4.65637295916417e-07
+ 6.44e+10    
+     4.65775270465118e-07
+     1.95088711667825e-07
+    4.511290819144492e-07
+    6.420654007419401e-08
+    1.260308142218824e-07
+    4.507056541699167e-07
+    3.076591366161206e-08
+    6.416723362528294e-08
+    1.954090347013844e-07
+    4.657977271911656e-07
+ 6.45e+10    
+    4.659351841304604e-07
+    1.951811621153747e-07
+       4.512473122802e-07
+    6.420221372197045e-08
+    1.260857807982603e-07
+    4.508240343423771e-07
+    3.072602820661851e-08
+    6.416278285045653e-08
+    1.955010873339339e-07
+    4.659583696191119e-07
+ 6.46e+10    
+    4.660953070687974e-07
+    1.952736278839574e-07
+    4.513656682246489e-07
+    6.419776926769218e-08
+     1.26140739032305e-07
+     4.50942539768408e-07
+    3.068604748504628e-08
+    6.415821434346056e-08
+     1.95593154629253e-07
+    4.661192233520336e-07
+ 6.47e+10    
+    4.662556394291347e-07
+    1.953661088289963e-07
+     4.51484149811152e-07
+    6.419320703151337e-08
+    1.261956889762981e-07
+    4.510611705130691e-07
+    3.064597236202591e-08
+    6.415352842276873e-08
+    1.956852364447354e-07
+    4.662802885427252e-07
+ 6.48e+10    
+    4.664161813614759e-07
+    1.954586048074669e-07
+      4.5160275710393e-07
+    6.418852733587358e-08
+     1.26250630683307e-07
+    4.511799266423005e-07
+    3.060580370459159e-08
+    6.414872540913957e-08
+    1.957773326393482e-07
+    4.664415653449979e-07
+ 6.49e+10    
+    4.665769330168223e-07
+    1.955511156778957e-07
+    4.517214901680669e-07
+    6.418373050547927e-08
+    1.263055642071823e-07
+    4.512988082229185e-07
+    3.056554238162813e-08
+    6.414380562559794e-08
+    1.958694430736278e-07
+     4.66603053913674e-07
+ 6.5e+10     
+    4.667378945471664e-07
+    1.956436413003559e-07
+    4.518403490695094e-07
+    6.417881686728495e-08
+    1.263604896025542e-07
+    4.514178153226152e-07
+    3.052518926381785e-08
+    6.413876939741667e-08
+    1.959615676096778e-07
+    4.667647544045846e-07
+ 6.51e+10    
+    4.668990661054904e-07
+    1.957361815364648e-07
+    4.519593338750625e-07
+    6.417378675047463e-08
+    1.264154069248294e-07
+    4.515369480099572e-07
+    3.048474522358718e-08
+    6.413361705209788e-08
+    1.960537061111647e-07
+    4.669266669745657e-07
+ 6.52e+10    
+    4.670604478457644e-07
+    1.958287362493804e-07
+    4.520784446523909e-07
+    6.416864048644249e-08
+    1.264703162301878e-07
+    4.516562063543836e-07
+    3.044421113505334e-08
+    6.412834891935401e-08
+    1.961458584433151e-07
+    4.670887917814551e-07
+ 6.53e+10    
+    4.672220399229398e-07
+    1.959213053037981e-07
+     4.52197681470016e-07
+    6.416337840877404e-08
+    1.265252175755791e-07
+    4.517755904262027e-07
+    3.040358787397065e-08
+    6.412296533108947e-08
+    1.962380244729122e-07
+    4.672511289840895e-07
+ 6.54e+10    
+    4.673838424929475e-07
+    1.960138885659465e-07
+    4.523170443973133e-07
+    6.415800085322687e-08
+    1.265801110187195e-07
+     4.51895100296593e-07
+    3.036287631767667e-08
+    6.411746662138092e-08
+    1.963302040682918e-07
+    4.674136787423005e-07
+ 6.55e+10    
+    4.675458557126962e-07
+    1.961064859035848e-07
+    4.524365335045121e-07
+    6.415250815771124e-08
+    1.266349966180882e-07
+    4.520147360375986e-07
+     3.03220773450385e-08
+    6.411185312645878e-08
+    1.964223970993386e-07
+    4.675764412169109e-07
+ 6.56e+10    
+    4.677080797400649e-07
+    1.961990971859984e-07
+    4.525561488626929e-07
+    6.414690066227081e-08
+    1.266898744329241e-07
+    4.521344977221291e-07
+    3.028119183639853e-08
+    6.410612518468761e-08
+     1.96514603437483e-07
+    4.677394165697323e-07
+ 6.57e+10    
+    4.678705147339042e-07
+    1.962917222839953e-07
+     4.52675890543786e-07
+    6.414117870906285e-08
+    1.267447445232221e-07
+    4.522543854239568e-07
+    3.024022067352045e-08
+    6.410028313654693e-08
+    1.966068229556963e-07
+    4.679026049635613e-07
+ 6.58e+10    
+    4.680331608540298e-07
+    1.963843610699021e-07
+    4.527957586205696e-07
+    6.413534264233884e-08
+    1.267996069497298e-07
+    4.523743992177155e-07
+    3.019916473953497e-08
+     6.40943273246118e-08
+    1.966990555284873e-07
+    4.680660065621765e-07
+ 6.59e+10    
+    4.681960182612207e-07
+    1.964770134175602e-07
+    4.529157531666672e-07
+    6.412939280842459e-08
+    1.268544617739435e-07
+    4.524945391788965e-07
+    3.015802491888535e-08
+    6.408825809353297e-08
+    1.967913010318977e-07
+    4.682296215303327e-07
+ 6.6e+10     
+    4.683590871172141e-07
+    1.965696792023216e-07
+    4.530358742565474e-07
+    6.412332955570037e-08
+    1.269093090581051e-07
+    4.526148053838502e-07
+    3.011680209727314e-08
+    6.408207579001773e-08
+    1.968835593434987e-07
+    4.683934500337625e-07
+ 6.61e+10    
+    4.685223675847062e-07
+     1.96662358301045e-07
+    4.531561219655193e-07
+      6.4117153234581e-08
+     1.26964148865198e-07
+    4.527351979097795e-07
+    3.007549716160344e-08
+    6.407578076280956e-08
+    1.969758303423856e-07
+    4.685574922391676e-07
+ 6.62e+10    
+    4.686858598273419e-07
+    1.967550505920905e-07
+    4.532764963697325e-07
+     6.41108641974957e-08
+    1.270189812589438e-07
+    4.528557168347424e-07
+    3.003411099993031e-08
+    6.406937336266862e-08
+    1.970681139091741e-07
+    4.687217483142185e-07
+ 6.63e+10    
+     4.68849564009718e-07
+    1.968477559553162e-07
+    4.533969975461747e-07
+    6.410446279886802e-08
+    1.270738063037982e-07
+    4.529763622376455e-07
+    2.999264450140227e-08
+    6.406285394235175e-08
+     1.97160409925996e-07
+    4.688862184275507e-07
+ 6.64e+10    
+    4.690134802973767e-07
+    1.969404742720741e-07
+    4.535176255726703e-07
+    6.409794939509572e-08
+    1.271286240649477e-07
+    4.530971341982458e-07
+    2.995109855620725e-08
+    6.405622285659236e-08
+    1.972527182764939e-07
+    4.690509027487603e-07
+ 6.65e+10    
+    4.691776088568032e-07
+    1.970332054252045e-07
+    4.536383805278762e-07
+    6.409132434453004e-08
+    1.271834346083053e-07
+     4.53218032797145e-07
+    2.990947405551806e-08
+    6.404948046208028e-08
+    1.973450388458172e-07
+    4.692158014484029e-07
+ 6.66e+10    
+    4.693419498554216e-07
+    1.971259492990317e-07
+    4.537592624912815e-07
+    6.408458800745573e-08
+    1.272382380005067e-07
+    4.533390581157896e-07
+    2.986777189143725e-08
+    6.404262711744129e-08
+    1.974373715206168e-07
+    4.693809146979861e-07
+ 6.67e+10    
+     4.69506503461592e-07
+    1.972187057793601e-07
+    4.538802715432053e-07
+    6.407774074607023e-08
+     1.27293034308907e-07
+    4.534602102364685e-07
+    2.982599295694248e-08
+     6.40356631832174e-08
+    1.975297161890409e-07
+    4.695462426699713e-07
+ 6.68e+10    
+    4.696712698446068e-07
+     1.97311474753468e-07
+    4.540014077647939e-07
+     6.40707829244632e-08
+    1.273478236015762e-07
+    4.535814892423098e-07
+    2.978413814583137e-08
+    6.402858902184571e-08
+    1.976220727407295e-07
+    4.697117855377651e-07
+ 6.69e+10    
+    4.698362491746881e-07
+     1.97404256110104e-07
+    4.541226712380186e-07
+    6.406371490859588e-08
+    1.274026059472955e-07
+    4.537028952172778e-07
+    2.974220835266672e-08
+     6.40214049976385e-08
+      1.9771444106681e-07
+    4.698775434757217e-07
+ 6.7e+10     
+    4.700014416229844e-07
+    1.974970497394817e-07
+    4.542440620456743e-07
+    6.405653706628027e-08
+    1.274573814155532e-07
+    4.538244282461738e-07
+    2.970020447272143e-08
+    6.401411147676222e-08
+    1.978068210598914e-07
+    4.700435166591337e-07
+ 6.71e+10    
+    4.701668473615664e-07
+    1.975898555332741e-07
+    4.543655802713757e-07
+    6.404924976715833e-08
+    1.275121500765409e-07
+    4.539460884146303e-07
+    2.965812740192356e-08
+    6.400670882721714e-08
+    1.978992126140598e-07
+    4.702097052642329e-07
+ 6.72e+10    
+    4.703324665634237e-07
+    1.976826733846092e-07
+    4.544872259995575e-07
+    6.404185338268112e-08
+    1.275669120011494e-07
+    4.540678758091109e-07
+    2.961597803680132e-08
+    6.399919741881653e-08
+     1.97991615624873e-07
+     4.70376109468185e-07
+ 6.73e+10    
+    4.704982994024627e-07
+     1.97775503188065e-07
+    4.546089993154694e-07
+    6.403434828608782e-08
+    1.276216672609645e-07
+    4.541897905169068e-07
+    2.957375727442823e-08
+    6.399157762316581e-08
+     1.98084029989355e-07
+    4.705427294490874e-07
+ 6.74e+10    
+     4.70664346053503e-07
+    1.978683448396633e-07
+    4.547309003051755e-07
+    6.402673485238471e-08
+    1.276764159282629e-07
+    4.543118326261342e-07
+    2.953146601236803e-08
+    6.398384981364183e-08
+    1.981764556059908e-07
+    4.707095653859649e-07
+ 6.75e+10    
+    4.708306066922718e-07
+     1.97961198236865e-07
+    4.548529290555517e-07
+    6.401901345832394e-08
+    1.277311580760085e-07
+    4.544340022257327e-07
+    2.948910514861978e-08
+    6.397601436537171e-08
+    1.982688923747212e-07
+     4.70876617458767e-07
+ 6.76e+10    
+    4.709970814954055e-07
+    1.980540632785657e-07
+    4.549750856542817e-07
+    6.401118448238272e-08
+    1.277858937778475e-07
+    4.545562994054632e-07
+    2.944667558156304e-08
+    6.396807165521208e-08
+    1.983613401969366e-07
+    4.710438858483639e-07
+ 6.77e+10    
+    4.711637706404406e-07
+    1.981469398650876e-07
+    4.550973701898581e-07
+    6.400324830474176e-08
+     1.27840623108105e-07
+    4.546787242559036e-07
+    2.940417820990298e-08
+    6.396002206172791e-08
+    1.984537989754725e-07
+    4.712113707365451e-07
+ 6.78e+10    
+    4.713306743058149e-07
+    1.982398278981772e-07
+     4.55219782751577e-07
+    6.399520530726403e-08
+    1.278953461417799e-07
+    4.548012768684472e-07
+    2.936161393261548e-08
+    6.395186596517136e-08
+    1.985462686146023e-07
+     4.71379072306013e-07
+ 6.79e+10    
+    4.714977926708626e-07
+    1.983327272809973e-07
+    4.553423234295363e-07
+    6.398705587347379e-08
+    1.279500629545418e-07
+     4.54923957335302e-07
+    2.931898364889261e-08
+    6.394360374746081e-08
+    1.986387490200337e-07
+    4.715469907403827e-07
+ 6.8e+10     
+    4.716651259158113e-07
+    1.984256379181227e-07
+     4.55464992314633e-07
+    6.397880038853476e-08
+    1.280047736227256e-07
+    4.550467657494846e-07
+    2.927628825808771e-08
+    6.393523579215939e-08
+     1.98731240098901e-07
+     4.71715126224178e-07
+ 6.81e+10    
+    4.718326742217786e-07
+    1.985185597155343e-07
+    4.555877894985629e-07
+      6.3970439239229e-08
+     1.28059478223328e-07
+    4.551697022048201e-07
+    2.923352865966089e-08
+     6.39267624844539e-08
+    1.988237417597602e-07
+    4.718834789428256e-07
+ 6.82e+10    
+    4.720004377707682e-07
+    1.986114925806122e-07
+    4.557107150738137e-07
+    6.396197281393523e-08
+    1.281141768340024e-07
+    4.552927667959388e-07
+    2.919070575312447e-08
+    6.391818421113328e-08
+    1.989162539125829e-07
+    4.720520490826558e-07
+ 6.83e+10    
+    4.721684167456691e-07
+    1.987044364221319e-07
+    4.558337691336675e-07
+     6.39534015026076e-08
+    1.281688695330558e-07
+     4.55415959618275e-07
+    2.914782043798862e-08
+     6.39095013605676e-08
+     1.99008776468751e-07
+    4.722208368308975e-07
+ 6.84e+10    
+    4.723366113302503e-07
+    1.987973911502566e-07
+    4.559569517721941e-07
+    6.394472569675383e-08
+    1.282235563994429e-07
+    4.555392807680608e-07
+     2.91048736137068e-08
+    6.390071432268615e-08
+     1.99101309341049e-07
+    4.723898423756732e-07
+ 6.85e+10    
+    4.725050217091581e-07
+    1.988903566765327e-07
+    4.560802630842513e-07
+    6.393594578941383e-08
+    1.282782375127627e-07
+    4.556627303423274e-07
+    2.906186617962178e-08
+    6.389182348895655e-08
+    1.991938524436603e-07
+    4.725590659059999e-07
+ 6.86e+10    
+    4.726736480679128e-07
+    1.989833329138825e-07
+    4.562037031654816e-07
+    6.392706217513796e-08
+    1.283329129532541e-07
+    4.557863084388999e-07
+    2.901879903491119e-08
+    6.388282925236278e-08
+     1.99286405692159e-07
+    4.727285076117824e-07
+ 6.87e+10    
+    4.728424905929073e-07
+    1.990763197765995e-07
+    4.563272721123085e-07
+    6.391807524996548e-08
+    1.283875828017908e-07
+    4.559100151563962e-07
+    2.897567307853381e-08
+      6.3873732007384e-08
+    1.993789690035049e-07
+    4.728981676838112e-07
+ 6.88e+10    
+     4.73011549471402e-07
+    1.991693171803411e-07
+     4.56450970021934e-07
+    6.390898541140261e-08
+    1.284422471398771e-07
+    4.560338505942215e-07
+    2.893248920917546e-08
+    6.386453214997276e-08
+    1.994715422960368e-07
+    4.730680463137607e-07
+ 6.89e+10    
+    4.731808248915212e-07
+    1.992623250421234e-07
+    4.565747969923385e-07
+    6.389979305840121e-08
+    1.284969060496439e-07
+    4.561578148525709e-07
+    2.888924832519523e-08
+    6.385523007753356e-08
+    1.995641254894669e-07
+    4.732381436941846e-07
+ 6.9e+10     
+    4.733503170422533e-07
+    1.993553432803147e-07
+    4.566987531222743e-07
+    6.389049859133668e-08
+    1.285515596138436e-07
+    4.562819080324204e-07
+    2.884595132457198e-08
+    6.384582618890112e-08
+    1.996567185048731e-07
+    4.734084600185121e-07
+ 6.91e+10    
+    4.735200261134452e-07
+     1.99448371814629e-07
+    4.568228385112664e-07
+    6.388110241198632e-08
+    1.286062079158457e-07
+     4.56406130235528e-07
+     2.88025991048508e-08
+    6.383632088431895e-08
+    1.997493212646944e-07
+    4.735789954810485e-07
+ 6.92e+10    
+    4.736899522957987e-07
+    1.995414105661201e-07
+    4.569470532596077e-07
+    6.387160492350758e-08
+    1.286608510396323e-07
+    4.565304815644313e-07
+    2.875919256308956e-08
+    6.382671456541739e-08
+    1.998419336927233e-07
+    4.737497502769675e-07
+ 6.93e+10    
+    4.738600957808707e-07
+    1.996344594571754e-07
+    4.570713974683563e-07
+    6.386200653041615e-08
+    1.287154890697936e-07
+    4.566549621224414e-07
+    2.871573259580596e-08
+    6.381700763519216e-08
+    1.999345557140995e-07
+    4.739207246023117e-07
+ 6.94e+10    
+    4.740304567610664e-07
+     1.99727518411509e-07
+    4.571958712393348e-07
+    6.385230763856427e-08
+    1.287701220915229e-07
+     4.56779572013643e-07
+    2.867222009892435e-08
+    6.380720049798256e-08
+    2.000271872553038e-07
+    4.740919186539873e-07
+ 6.95e+10    
+    4.742010354296396e-07
+    1.998205873541559e-07
+    4.573204746751251e-07
+    6.384250865511877e-08
+    1.288247501906129e-07
+    4.569043113428917e-07
+    2.862865596772297e-08
+    6.379729355944978e-08
+    2.001198282441514e-07
+    4.742633326297631e-07
+ 6.96e+10    
+    4.743718319806868e-07
+    1.999136662114652e-07
+    4.574452078790679e-07
+    6.383260998853925e-08
+    1.288793734534498e-07
+    4.570291802158085e-07
+    2.858504109678129e-08
+     6.37872872265551e-08
+     2.00212478609785e-07
+     4.74434966728266e-07
+ 6.97e+10    
+    4.745428466091473e-07
+    2.000067549110934e-07
+    4.575700709552569e-07
+     6.38226120485562e-08
+    1.289339919670093e-07
+    4.571541787387794e-07
+     2.85413763799276e-08
+    6.377718190753831e-08
+    2.003051382826687e-07
+    4.746068211489791e-07
+ 6.98e+10    
+    4.747140795107993e-07
+     2.00099853381999e-07
+    4.576950640085405e-07
+    6.381251524614933e-08
+    1.289886058188527e-07
+    4.572793070189519e-07
+    2.849766271018673e-08
+    6.376697801189573e-08
+     2.00397807194581e-07
+    4.747788960922377e-07
+ 6.99e+10    
+    4.748855308822547e-07
+    2.001929615544345e-07
+     4.57820187144514e-07
+    6.380231999352531e-08
+    1.290432150971206e-07
+    4.574045651642326e-07
+    2.845390097972792e-08
+    6.375667595035865e-08
+    2.004904852786084e-07
+    4.749511917592278e-07
+ 7e+10       
+    4.750572009209595e-07
+    2.002860793599409e-07
+    4.579454404695213e-07
+     6.37920267040962e-08
+    1.290978198905292e-07
+    4.575299532832819e-07
+    2.841009207981307e-08
+    6.374627613487148e-08
+    2.005831724691381e-07
+    4.751237083519819e-07
* NOTE: Solution at 1e+08 Hz used as DC point.

.model g_m4lines_port_1 sp N=4 SPACING=nonuniform VALTYPE=real
+ INTERPOLATION=spline
+ DATA = 700
+ 0           
+    0.0008625639485742468
+   -0.0001648424890465852
+    0.0008704502393055881
+   -1.131980998041023e-06
+   -6.997825681320198e-05
+    0.0008682078926154774
+    1.891793655724844e-07
+   -1.163263054663917e-06
+   -0.0001645904670047619
+    0.0008643958326090265
+ 2e+08       
+     0.001801008666589373
+   -0.0003566931862677911
+     0.001822473152308518
+   -1.670221319520845e-06
+   -0.0001516255535572703
+     0.001819149675254844
+     -1.2969556981752e-06
+   -1.760025138819056e-06
+   -0.0003571097875232234
+     0.001805155202781535
+ 3e+08       
+     0.002627997480741298
+   -0.0005074027002600783
+     0.002655532659538103
+   -4.194723723644677e-06
+   -0.0002146107953591286
+     0.002649856934038569
+   -6.903757770653383e-07
+   -4.338498924753106e-06
+   -0.0005069597962626945
+     0.002633700275531452
+ 4e+08       
+     0.003457615432385194
+   -0.0006609611433716831
+     0.003490530213143012
+   -5.180834650121862e-06
+   -0.0002799811309286256
+     0.003482149117782107
+    3.387341055123298e-07
+   -5.333188021696124e-06
+   -0.0006600053310387597
+     0.003464963535880437
+ 5e+08       
+      0.00430876955691653
+   -0.0008225518201561701
+     0.004348023426139348
+    -5.56033188530456e-06
+   -0.0003488583298650385
+     0.004336984583073532
+    1.136913136464673e-06
+   -5.721515821264115e-06
+   -0.0008212911779741628
+      0.00431788384733446
+ 6e+08       
+     0.005169468381852566
+   -0.0009870862010409008
+     0.005215953319131178
+   -6.091774527363477e-06
+   -0.0004187217817258212
+     0.005202466791705683
+    1.687323632629368e-06
+   -6.274545545065477e-06
+   -0.0009855705745006639
+     0.005180395420935325
+ 7e+08       
+     0.006029617880561672
+    -0.001151040518544732
+     0.006083790414804052
+   -6.928907318293624e-06
+   -0.0004881365076699089
+     0.006068074580208911
+    2.135648685128547e-06
+   -7.141894124602379e-06
+    -0.001149272963428848
+     0.006042359428637471
+ 8e+08       
+     0.006886436684547718
+    -0.001313707205208065
+      0.00694834311478585
+   -7.889852065127529e-06
+   -0.0005569186892929223
+     0.006930516217613721
+     2.61437516279021e-06
+   -8.135153067935811e-06
+    -0.001311685579149925
+     0.006900981640998201
+ 9e+08       
+     0.007742587427504242
+    -0.001476170061089323
+      0.00781207358847117
+   -8.691893157829463e-06
+    -0.000625591028468161
+     0.007792102391996755
+    3.207615935813026e-06
+   -8.967245715929751e-06
+    -0.001473895010356015
+     0.007758932929820467
+ 1e+09       
+     0.008603508045135577
+    -0.001640273141283548
+     0.008680516422904273
+    -9.07049029467961e-06
+   -0.0006949498722108631
+     0.008658211981492503
+    3.961235314617779e-06
+   -9.371710753998017e-06
+    -0.001637747578022007
+     0.008621671946039621
+ 1.1e+09     
+     0.009480532818627027
+    -0.001779227543447545
+     0.009557094230670686
+   -6.706790096732237e-06
+   -0.0007592169281512265
+     0.009530130392426079
+    1.126095676817585e-05
+   -7.282032989474761e-06
+    -0.001775336372251179
+     0.009500043498760978
+ 1.2e+09     
+      0.01035907632026234
+    -0.001926116476009326
+      0.01043628468847772
+   -4.454623462753174e-06
+     -0.00082534896200912
+      0.01040479443499359
+    1.921364507436414e-05
+   -5.277557964244127e-06
+    -0.001921077936742385
+       0.0103800260962127
+ 1.3e+09     
+      0.01123608236746707
+    -0.002079101535379419
+      0.01131496348381693
+   -2.470801701311174e-06
+   -0.0008926891335817984
+       0.0112791400931016
+    2.738365151365605e-05
+   -3.509264497018481e-06
+    -0.002073105757821298
+      0.01125854537337876
+ 1.4e+09     
+      0.01210980750098187
+    -0.002236622408230177
+      0.01219131817178826
+   -8.353881069625576e-07
+   -0.0009607413080937018
+      0.01215140001305758
+    3.535755530369706e-05
+   -2.053795289962319e-06
+    -0.002229833859586287
+      0.01213384456051502
+ 1.5e+09     
+      0.01297939817860109
+    -0.002397390043041374
+      0.01306442734671108
+    4.330995886264087e-07
+    -0.001029141737540308
+      0.01302068386536439
+     4.27749110997294e-05
+    -9.28430167782717e-07
+    -0.002389950807866811
+      0.01300506059042255
+ 1.6e+09     
+      0.01384458247641268
+    -0.002560361878653058
+       0.0139339531241501
+    1.360070690018008e-06
+    -0.001097630960209699
+      0.01388667260804305
+     4.93487393271428e-05
+   -1.083238840202095e-07
+    -0.002552394951018313
+      0.01387191474059615
+ 1.7e+09     
+      0.01470545304702728
+    -0.002724710072272164
+      0.01479992465541726
+    1.998405339924511e-06
+      -0.0011660292764528
+      0.01474940404676393
+     5.48763190393621e-05
+     4.57472948908104e-07
+      -0.0027163223040195
+        0.014734494721126
+ 1.8e+09     
+      0.01556231844234982
+    -0.002889788816776836
+      0.01566259004973839
+    2.414900117036727e-06
+    -0.001234216794129836
+        0.015609126807248
+    5.924145701525769e-05
+    8.328826306679702e-07
+    -0.002881073412828281
+      0.01559310535125761
+ 1.9e+09     
+      0.01641560359083812
+     -0.00305510378289559
+      0.01652231743402621
+    2.680152614436498e-06
+    -0.001302117850969518
+       0.0164662032689749
+     6.24097993838822e-05
+    1.085057327731003e-06
+    -0.003046142348783525
+      0.01644816858913071
+ 2e+09       
+      0.01726578462608229
+    -0.003220284956208591
+      0.01737953019374584
+     2.86172226178153e-06
+    -0.001369689145009689
+      0.01732104639593543
+    6.441896491471904e-05
+    1.277843973667586e-06
+    -0.003211149144762524
+      0.01730015806517255
+ 2.1e+09     
+      0.01811334723746977
+    -0.003385063191456276
+      0.01823466543591309
+    3.020054801621298e-06
+    -0.001436910802279866
+       0.0181740794576215
+    6.536532529297605e-05
+    1.467941149538407e-06
+    -0.003375816002733222
+      0.01814955724332239
+ 2.2e+09     
+      0.01895876088304134
+    -0.003549250339126737
+      0.01908814794969781
+    3.206533127815985e-06
+    -0.001503779678417697
+      0.01902571091273412
+    6.538915025427528e-05
+    1.703115629475213e-06
+    -0.003539947121471145
+        0.018996833512055
+ 2.3e+09     
+      0.01980246356560969
+    -0.003712722596733472
+      0.01994037436738258
+    3.463026969567805e-06
+     -0.00157030431751671
+      0.01987631918638065
+     6.46596012971054e-05
+    2.021860282440499e-06
+    -0.003703411787974499
+      0.01984242287869131
+ 2.4e+09     
+      0.02064485355994174
+    -0.003875406673054916
+      0.02079170396590697
+    3.822395905122547e-06
+    -0.001636501124006274
+      0.02072624382860512
+     6.33607382175862e-05
+    2.453958574867945e-06
+    -0.003866130313873489
+      0.02068672163680088
+ 2.5e+09     
+      0.02148628565240467
+    -0.004037268357433601
+      0.02164245375444146
+    4.309513039335423e-06
+    -0.001702391419844939
+      0.02157578075811474
+    6.167934638973697e-05
+    3.021533728820225e-06
+    -0.004028062405229738
+      0.02153008255763151
+ 2.6e+09     
+      0.02232707025779117
+    -0.004198303120508525
+      0.02249289631179186
+    4.942493930910246e-06
+    -0.001767999153322573
+      0.02242518011777445
+    5.979504541675295e-05
+    3.740276947249762e-06
+    -0.004189197591524588
+      0.02237281396520047
+ 2.7e+09     
+      0.02316747432280739
+    -0.004358528418274802
+      0.02334325938516166
+    5.733921332166586e-06
+     -0.00183334909775157
+      0.02327464581587868
+    5.787283702892983e-05
+    4.620653812864952e-06
+    -0.004349547387528147
+      0.02321518060299571
+ 2.8e+09     
+      0.02400772329356373
+    -0.004517977418682166
+      0.02419372662482678
+     6.69194312894943e-06
+    -0.001898465431298164
+      0.02412433618657647
+    5.605801323706861e-05
+    5.668973395100757e-06
+    -0.004509138910507378
+      0.02405740557022595
+ 2.9e+09     
+      0.02484800367259772
+    -0.004676693914659491
+      0.02504443906806244
+    7.821186139688778e-06
+    -0.001963370626776094
+      0.02497436543539881
+    5.447318199057591e-05
+    6.888268504245672e-06
+    -0.004668009720454518
+      0.02489967285485561
+ 3e+09       
+      0.02568846585858171
+     -0.00483472822755026
+      0.02589549714133881
+    9.123473309914347e-06
+    -0.002028084605791906
+      0.02582480568322027
+    5.321707287241724e-05
+    8.278979136746851e-06
+    -0.004826203690845614
+      0.02574213015868184
+ 3.1e+09     
+      0.02652922707522661
+    -0.004992133939750981
+      0.02674696304969195
+    1.059835947180003e-05
+    -0.002092624128083329
+      0.02667568951179786
+    5.236474838142069e-05
+     9.83945763042616e-06
+    -0.004983767751265933
+       0.0265848918229863
+ 3.2e+09     
+      0.02737037427252287
+    -0.005148965324750708
+       0.0275988634841637
+    1.224351516941235e-05
+    -0.002157002396566876
+       0.0275270129643975
+    5.196885253757542e-05
+    1.156632733275559e-05
+    -0.005140749371063153
+       0.0274280417395156
+ 3.3e+09     
+      0.02821196693501919
+    -0.005305275366971863
+      0.02845119261395479
+     1.40549929886305e-05
+    -0.002221228863345719
+      0.02837873897792626
+    5.206156320586812e-05
+    1.345473057947787e-05
+    -0.005297194675335884
+      0.02827163618249131
+ 3.4e+09     
+      0.02905403976610703
+    -0.005461114283180158
+      0.02930391534714077
+    1.602740976828299e-05
+    -0.002285309223147406
+      0.02923080122660399
+    5.265696486315502e-05
+    1.549849987129189e-05
+    -0.005453147101552036
+      0.02911570653087334
+ 3.5e+09     
+      0.02989660523946937
+    -0.005616528472244812
+      0.03015697084773015
+    1.815407367070875e-05
+    -0.002349245579473903
+      0.03008310834747821
+     5.37536145704088e-05
+    1.769028098837016e-05
+    -0.005608646517583413
+      0.02996026187148531
+ 3.6e+09     
+      0.03073965602251604
+    -0.005771559831246746
+      0.03101027629133919
+    2.042707926893713e-05
+    -0.002413036766035733
+      0.03093554849971743
+    5.533712871127366e-05
+    2.002163031926288e-05
+    -0.005763728730710969
+      0.03080529148646229
+ 3.7e+09     
+      0.03158316728421795
+    -0.005926245383966139
+      0.03186373082987392
+    2.283738781451425e-05
+    -0.002476678802533954
+      0.03178799418666487
+    5.738266735553241e-05
+    2.248310216873626e-05
+    -0.005918425323044612
+      0.03165076723530565
+ 3.8e+09     
+      0.03242709890300541
+    -0.006080617173280831
+      0.03271721971998978
+     2.53749044106405e-05
+    -0.002540165460166677
+      0.03264030724575349
+    5.985723477072626e-05
+    2.506433599367103e-05
+    -0.006072763752695461
+      0.03249664584441379
+ 3.9e+09     
+      0.03327139759056971
+    -0.006234702372633317
+       0.0335706185531375
+    2.802855927521683e-05
+    -0.002603488908903385
+      0.03349234388988545
+    6.272174802945593e-05
+    2.775414876074597e-05
+    -0.006226767662801572
+      0.03334287111661111
+ 4e+09       
+      0.03411599894545334
+    -0.006388523574125542
+      0.03442379750891657
+    3.078639673336904e-05
+    -0.002666640416043245
+      0.03434395966761686
+    6.593285121831588e-05
+    3.054063403102225e-05
+    -0.006380457342934225
+      0.03418937607089469
+ 4.1e+09     
+      0.03496082944695344
+    -0.006542099212576703
+      0.03527662554021611
+    3.363567297608402e-05
+     -0.00272961106421142
+      0.03519501420069983
+    6.944447137013931e-05
+     3.34112669023107e-05
+    -0.006533850290169002
+      0.03503608501912146
+ 4.2e+09     
+      0.03580580839567603
+    -0.006695444086558072
+      0.03612897438987588
+    3.656296183456465e-05
+    -0.002792392456997393
+      0.03604537555765153
+    7.320912507300683e-05
+    3.635301244018108e-05
+    -0.006686961820685225
+       0.0358829155822354
+ 4.3e+09     
+      0.03665084980252024
+    -0.006848569939422866
+      0.03698072233555204
+    3.955426669688899e-05
+    -0.002854977382017159
+      0.03689492413154377
+    7.717899294475724e-05
+    3.935243452320375e-05
+    -0.006839805687447251
+      0.03672978064434857
+ 4.4e+09     
+      0.03749586422332053
+    -0.007001486065976019
+      0.03783175756278768
+    4.259513608731693e-05
+    -0.002917360404262016
+      0.03774355590866908
+    8.130678389481154e-05
+     4.23958019287133e-05
+    -0.006992394665390049
+      0.03757659023887165
+ 4.5e+09     
+      0.03834076053212017
+    -0.007154199913835871
+      0.03868198107602774
+    4.567078020919647e-05
+    -0.002979538367015485
+      0.03859118504075786
+    8.554641326671505e-05
+    4.546918881322723e-05
+    -0.007144741072450314
+      0.03842325335721034
+ 4.6e+09     
+      0.03918544762233347
+    -0.007306717652749573
+      0.03953130907294251
+    4.876618581310042e-05
+    -0.003041510783090116
+      0.03943774566488924
+    8.985351933256424e-05
+    4.855856733690335e-05
+    -0.007296857202452599
+      0.03926967966747733
+ 4.7e+09     
+      0.04002983602204022
+     -0.00745904469002693
+      0.04037967472784747
+    5.186622700721779e-05
+    -0.003103280105280513
+      0.04028319294957792
+    9.418584179476692e-05
+    5.164989090961406e-05
+    -0.007448755653870917
+      0.04011578112835181
+ 4.8e+09     
+      0.04087383940748322
+    -0.007611186115649668
+         0.04122702935372
+    5.495577000990979e-05
+    -0.003164851871319208
+      0.04112750337998975
+    9.850348439326443e-05
+    5.472916729017466e-05
+    -0.007600449546379409
+      0.04096147348172663
+ 4.9e+09     
+      0.04171737599756296
+     -0.00776314706621489
+      0.04207334293755006
+    5.801977030135371e-05
+    -0.003226234724828259
+      0.04197067432725547
+    0.0001027690817457942
+     5.77825214702263e-05
+     -0.00775195262443862
+      0.04180667760715864
+ 5e+09       
+      0.04256036981179542
+    -0.007914933002381361
+      0.04291860406868784
+    6.104336111909672e-05
+    -0.003287440319387159
+      0.04281272297423135
+    0.0001069478883945693
+    6.079624886643408e-05
+    -0.007903279253557754
+      0.04265132072139453
+ 5.1e+09     
+      0.04340275177479329
+    -0.008066549899605131
+      0.04376281930275383
+    6.401193272600342e-05
+     -0.00334848311757138
+       0.0436536846912442
+     0.000111007805849637
+    6.375685979917944e-05
+     -0.00805444432006064
+      0.04349533740736158
+ 5.2e+09     
+      0.04424446065181276
+    -0.008218004356422389
+      0.04460601202311378
+    6.691120232954129e-05
+    -0.003409380100435861
+      0.04449361096947355
+    0.0001149193613059901
+    6.665111654283423e-05
+    -0.008205463049014984
+      0.04433867045894931
+ 5.3e+09     
+       0.0450854438022014
+     -0.00836930362817153
+      0.04544822087686279
+    6.972727492617417e-05
+    -0.003470150405316033
+      0.04533256702651163
+    0.0001186556497278862
+    6.946606439758515e-05
+    -0.008356350757443436
+      0.04518127153058906
+ 5.4e+09     
+      0.04592565774057179
+    -0.008520455596729617
+      0.04628949787211756
+    7.244669566730999e-05
+    -0.003530814910992285
+      0.04617062919875067
+    0.0001221922491721046
+    7.218905827276537e-05
+    -0.008507122561108901
+      0.04602310158397087
+ 5.5e+09     
+      0.04676506849908989
+    -0.008671468688540436
+      0.04712990622806122
+    7.505649458394915e-05
+    -0.003591395789301947
+       0.0470078822295061
+    0.0001255071175762732
+    7.480778621053968e-05
+    -0.008657793053227928
+      0.04686413112809002
+ 5.6e+09     
+      0.04760365178824642
+    -0.008822351753974184
+      0.04796951806891326
+    7.754422466228463e-05
+    -0.003651916041346464
+      0.04784441655144032
+    0.0001285804777717567
+    7.731029114310889e-05
+    -0.008808375972637127
+      0.04770434025304156
+ 5.7e+09     
+      0.04844139295770732
+    -0.008973113920983794
+      0.04880841204842325
+    7.989799433461009e-05
+    -0.003712399034735756
+      0.04868032564828552
+    0.0001313946961882846
+    7.968499199255863e-05
+    -0.008958883877461899
+      0.04854371846240663
+ 5.8e+09     
+      0.04927828676313987
+    -0.009123764435253335
+      0.04964667098345484
+    8.210649544635324e-05
+    -0.003772868056062488
+      0.04951570356543961
+    0.0001339341595912935
+    8.192070501376251e-05
+    -0.009109327838446181
+      0.04938226431351707
+ 5.9e+09     
+      0.05011433694910116
+    -0.009274312497733453
+       0.0504843795646988
+     8.41590276927266e-05
+    -0.003833345890229313
+      0.05035064262297415
+    0.0001361851532214028
+    8.400666606651766e-05
+    -0.009259717164002954
+      0.05021998487915001
+ 6e+09       
+      0.05094955566199282
+     -0.00942476710879863
+      0.05132162220050674
+    8.604552040104504e-05
+    -0.003893854435565086
+      0.05118523136897462
+    0.0001381357428769919
+    8.593255429828646e-05
+    -0.009410059166902652
+      0.05105689504811666
+ 6.1e+09     
+      0.05178396271055886
+    -0.009575136926395935
+      0.05215848103717519
+    8.775655238273897e-05
+    -0.003954414361032758
+      0.05201955279671276
+    0.0001397756627824016
+    8.768851753347576e-05
+     -0.00956035898044643
+      0.05189301668559271
+ 6.2e+09     
+      0.05261758469431723
+     -0.00972543014362743
+      0.05299503418652313
+    8.928337040744637e-05
+    -0.004015044809383988
+      0.05285368283646277
+    0.0001410962105033856
+     8.92651995046366e-05
+    -0.009710619430050776
+      0.05272837767676446
+ 6.3e+09     
+      0.05345045402255359
+    -0.009875654389328319
+      0.05383135417990526
+    9.061790667389143e-05
+    -0.004075763147947097
+      0.05368768912211262
+    0.0001420901496955492
+    9.065376892797858e-05
+    -0.009860840964432245
+      0.05356301087932205
+ 6.4e+09     
+      0.05428260784800526
+     -0.01002581665345605
+      0.05466750665734953
+     9.17527954807426e-05
+    -0.004136584766900034
+      0.05452163002418008
+    0.0001427516210883288
+    9.184595031927869e-05
+     -0.01001102164903137
+      0.05439695301145837
+ 6.5e+09     
+      0.05511408694009716
+     -0.01017592323754994
+      0.05550354929156394
+    9.268138914450601e-05
+     -0.00419752292340149
+       0.0553555539343721
+    0.0001430760618050207
+    9.283405636473729e-05
+     -0.01016115722294097
+      0.05523024350231648
+ 6.6e+09     
+      0.05594493452256165
+     -0.01032597972919345
+      0.05633953093926952
+    9.339777307750517e-05
+    -0.004258588628827396
+      0.05618949878224534
+     0.000143060132887304
+    9.361102160056894e-05
+     -0.01031124121937114
+      0.05606292333127545
+ 6.7e+09     
+      0.05677519509952472
+     -0.01047599099832333
+      0.05717549100667678
+    9.389677983162738e-05
+    -0.004319790575563773
+      0.05702349176161067
+    0.0001427016547202757
+     9.41704371119601e-05
+     -0.01046126514856872
+      0.05689503388115722
+ 6.8e+09     
+      0.05760491329274827
+     -0.01062596121239106
+       0.0580114590118555
+    9.417400183446317e-05
+    -0.004381135099303794
+      0.05785754924279026
+    0.0001419995499316185
+    9.450658593125778e-05
+     -0.01061121874107062
+      0.05772661582844182
+ 6.9e+09     
+       0.0584341327107728
+     -0.01077589386677342
+      0.05884745432409028
+    9.422580249421195e-05
+    -0.004442626172544119
+      0.05869167684641707
+    0.0001409537932573648
+    9.461447879412525e-05
+     -0.01076109024819234
+      0.05855770809103683
+ 7e+09       
+      0.05926289486832896
+     -0.01092579182644631
+       0.0596834860588849
+    9.404932532610332e-05
+    -0.004504265424927186
+      0.05952586965489744
+    0.0001395653678189863
+    9.448988989680307e-05
+     -0.01091086679570962
+      0.05938834685117132
+ 7.1e+09     
+      0.06009123817169325
+     -0.01107565737474825
+      0.06051955310686425
+    9.364250075419658e-05
+    -0.004566052186186356
+      0.06036011253869311
+    0.0001378362272352262
+    9.412939228511073e-05
+     -0.01106053478577529
+      0.06021856466772605
+ 7.2e+09     
+      0.06091919698278943
+     -0.01122549226505545
+        0.061355644275215
+    9.300405026421216e-05
+    -0.004627983547679276
+      0.06119438057603235
+    0.0001357692629911438
+      9.3530392494249e-05
+     -0.01121008034122382
+      0.06104838968890255
+ 7.3e+09     
+       0.0617468007718923
+     -0.01137529777133782
+      0.06219173852131748
+    9.213348762199703e-05
+     -0.00469005443880356
+      0.06202863954635108
+     0.000133368276501064
+    9.269116404658512e-05
+     -0.01135948978555635
+      0.06187784497270955
+ 7.4e+09     
+      0.06257407336589035
+     -0.01152507473384632
+      0.06302780525966341
+    9.103111692423835e-05
+    -0.004752257714947182
+      0.06286284647957276
+    0.0001306379553272763
+    9.161087940160514e-05
+     -0.01150875015108274
+      0.06270694791941238
+ 7.5e+09     
+      0.06340103229630099
+     -0.01167482359657153
+      0.06386380472488752
+    8.969802730919346e-05
+    -0.004814584254008773
+      0.06369695024515729
+    0.0001275838530486856
+     9.02896399382039e-05
+     -0.01165784970694057
+      0.06353570981696294
+ 7.6e+09     
+      0.06422768824868148
+     -0.01182454443358777
+      0.06469968837563267
+    8.813608422188093e-05
+    -0.004877023058909243
+      0.06453089216662096
+    0.0001242123723105637
+    8.872850353485416e-05
+     -0.01180677849803403
+      0.06436413549757115
+ 7.7e+09     
+      0.06505404461279853
+      -0.0119742369619335
+      0.06553539932591342
+    8.634791719677786e-05
+    -0.004939561363892483
+      0.06536460664890374
+    0.0001205307506257827
+    8.692950929919735e-05
+     -0.01195552888536049
+      0.06519222310106113
+ 7.8e+09     
+      0.06588009713095319
+     -0.01212390053925746
+       0.0663708727925746
+    8.433690418910403e-05
+    -0.005002184742766934
+      0.06619802180751098
+    0.0001165470485379155
+    8.489569898649692e-05
+     -0.01210409607774243
+      0.06601996393851331
+ 7.9e+09     
+      0.06670583364021566
+     -0.01227353414505631
+      0.06720603654928703
+    8.210715255051231e-05
+    -0.005064877217566616
+      0.06703106008978131
+    0.0001122701397961838
+    8.263113463785783e-05
+     -0.01225247864468041
+      0.06684734244794924
+ 8e+09       
+       0.0675312339030192
+     -0.01242313634492459
+      0.06804081137925037
+    7.966347680441062e-05
+    -0.005127621366403709
+      0.06786363887992299
+    0.0001077097032308857
+    8.014091196639371e-05
+     -0.01240067899990838
+      0.06767433623247232
+ 8.1e+09     
+      0.06835626951958443
+     -0.01257270523781602
+       0.0688751115203534
+     7.70113734291712e-05
+    -0.005190398429544963
+      0.06869567108063353
+    0.0001028762160550565
+    7.743116902387583e-05
+     -0.01254870384528831
+      0.06850091617033457
+ 8.2e+09     
+      0.06918090391496651
+     -0.01272223838685479
+      0.06970884509795902
+    7.415699290247196e-05
+    -0.005253188412970329
+      0.06952706566518449
+    9.778094835390951e-05
+    7.450908969455425e-05
+     -0.01269656456493838
+      0.06932704658582221
+ 8.3e+09     
+      0.07000509239312018
+     -0.01287173273472731
+      0.07054191454172884
+    7.110710929696844e-05
+    -0.005315970188865098
+      0.07035772819482933
+    9.243595855777209e-05
+    7.138290158770211e-05
+     -0.01284427755996316
+      0.07015268546963299
+ 8.4e+09     
+      0.07082878225021899
+     -0.01302118450511427
+      0.07137421698398204
+    6.786908774559261e-05
+    -0.005378721592659837
+       0.0711875612972962
+    8.685408972744415e-05
+    6.806186793778361e-05
+     -0.01299186451484984
+      0.07097778473750722
+ 8.5e+09     
+       0.0716519129395158
+     -0.01317058909198417
+      0.07220564463800318
+    6.445085011451022e-05
+    -0.005441419516366846
+      0.07201646510297539
+    8.104896651289664e-05
+    6.455627317191685e-05
+     -0.01313935258751236
+       0.0718022905162419
+ 8.6e+09     
+       0.0724744162802476
+     -0.01331994093885259
+      0.07303608515547258
+    6.086083923307424e-05
+    -0.005504039998070833
+      0.07284433763621793
+    7.503499267778792e-05
+      6.0877401868636e-05
+     -0.01328677451610055
+      0.07262614344682135
+ 8.7e+09     
+      0.07329621670343878
+      -0.0134692334103204
+      0.07386542196282045
+    5.710798203405497e-05
+    -0.005566558307519101
+      0.07367107515993294
+    6.882734911317526e-05
+    5.703751091035419e-05
+      -0.0134341686370301
+      0.07344927899520329
+ 8.8e+09     
+      0.07411723152790456
+     -0.01361845865833168
+      0.07469353457679968
+    5.320165195394169e-05
+    -0.005628949027823733
+      0.07449657247242743
+    6.244199229454178e-05
+    5.304979472256673e-05
+     -0.01358157881021177
+      0.07427162776225685
+ 8.9e+09     
+      0.07493737126027349
+     -0.01376760748564718
+      0.07552029889995071
+    4.915163093384563e-05
+    -0.005691186133339442
+      0.07532072315615984
+    5.589565316675184e-05
+    4.892834359559442e-05
+      -0.0137290542491357
+      0.07509311578542752
+ 9e+09       
+      0.07575653991340277
+     -0.01391666920901233
+       0.0763455874969137
+    4.496807134679901e-05
+    -0.005753243063817869
+      0.07614341977879678
+    4.920583647170904e-05
+    4.468809519642125e-05
+     -0.01387664925526657
+      0.07591366482586612
+ 9.1e+09     
+      0.07657463533813538
+     -0.01406563152441932
+      0.07716926985273591
+    4.066145815804345e-05
+    -0.005815092794963951
+      0.07696455404765538
+    4.239082056337875e-05
+    4.034477949690571e-05
+      -0.0140244228580829
+      0.07673319263595989
+ 9.2e+09     
+      0.07739154956392139
+     -0.01421448037672841
+      0.07799121261444369
+    3.624257160264572e-05
+    -0.005876707905536344
+      0.07778401691928002
+    3.546965778383543e-05
+    3.591485746679175e-05
+     -0.01417243836400535
+      0.07755161320342632
+ 9.3e+09     
+      0.07820716914438323
+     -0.01436319983573125
+      0.07881127981720636
+    3.172245063911926e-05
+    -0.005938060641141218
+      0.07860169866653659
+    2.846217550217132e-05
+    3.141545400257807e-05
+     -0.01432076281935163
+      0.07836883696932254
+ 9.4e+09     
+      0.07902137550443433
+     -0.01451177198052163
+      0.07962933309642976
+    2.711235741136324e-05
+    -0.005999122974871283
+      0.07941748890619507
+    2.138897794459011e-05
+    2.686428568173969e-05
+     -0.01446946639427731
+      0.07918477101848265
+ 9.5e+09     
+      0.07983404528605746
+     -0.01466017679379354
+      0.08044523188708774
+     2.24237429226593e-05
+    -0.006059866664939037
+       0.0802312765905026
+    1.427144896857971e-05
+    2.227958404303967e-05
+     -0.01461862169635952
+      0.07999931924196832
+ 9.6e+09     
+      0.08064505069030541
+     -0.01480839206742351
+      0.08125883361154027
+    1.766821409723927e-05
+    -0.006120263309447717
+      0.08104294996671631
+    7.131755956143451e-06
+    1.768001519318651e-05
+     -0.01476830302400291
+      0.08081238247211306
+ 9.7e+09     
+      0.08145425981349917
+     -0.01495639332042238
+      0.08206999385700689
+    1.285750237647816e-05
+    -0.006180284398435059
+      0.08185239650894725
+   -7.144979921516054e-09
+     1.30845966248563e-05
+     -0.01491858557114548
+       0.0816238585916092
+ 9.8e+09     
+      0.08226153697596922
+     -0.01510415373006828
+      0.08287856654376589
+     8.00343396874226e-06
+    -0.006239901363315764
+      0.08265950282696702
+   -7.121502267158977e-06
+    8.512612197570431e-06
+     -0.01506954459577989
+      0.08243364261884172
+ 9.9e+09     
+      0.08306674304201439
+     -0.01525164407676748
+      0.08368440408504954
+    3.117901845009225e-06
+    -0.006299085623838944
+      0.08346415455683109
+   -1.418676040072136e-05
+    3.983526278727566e-06
+     -0.01522125456554506
+      0.08324162677228382
+ 1e+10       
+      0.08386973573003725
+     -0.01539883270293341
+      0.08448735753949155
+   -1.787160453532569e-06
+    -0.006357808632666265
+       0.0842662362382663
+   -2.117754949797017e-05
+   -4.831019343514917e-07
+     -0.01537378829406591
+      0.08404770051724203
+ 1.01e+10    
+      0.08470798959986381
+     -0.01554062362857664
+      0.08531877221044902
+   -7.092743096723687e-06
+    -0.006420083217346269
+      0.08509580812300417
+   -2.877728909897632e-05
+   -5.754620057981698e-06
+     -0.01551517727946193
+      0.08488743761393766
+ 1.02e+10    
+      0.08554521292379391
+     -0.01568269276821771
+      0.08614941562485755
+   -1.252800812870586e-05
+    -0.006482347279154904
+      0.08592460188826651
+   -3.656826092712372e-05
+   -1.115544117769474e-05
+     -0.01565685313063418
+      0.08572615588763692
+ 1.03e+10    
+      0.08638135859459609
+     -0.01582502605194324
+       0.0869792566041778
+   -1.809533108593231e-05
+    -0.006544594789863485
+      0.08675258532725286
+   -4.455220467378183e-05
+   -1.668804655895802e-05
+     -0.01579880135751934
+      0.08656380802533689
+ 1.04e+10    
+      0.08721638279236538
+     -0.01596760972918152
+       0.0878082668422738
+   -2.379697732289338e-05
+    -0.006606820007287356
+      0.08757972917964224
+   -5.273071411300242e-05
+   -2.235480330147963e-05
+     -0.01594100779964833
+       0.0874003499879429
+ 1.05e+10    
+      0.08805024489620507
+     -0.01611043036912044
+      0.08863642079586531
+   -2.963510118669885e-05
+    -0.006669017474259986
+      0.08840600702225253
+    -6.11052364041971e-05
+   -2.815796339834201e-05
+     -0.01608345862691457
+      0.08823574092188576
+ 1.06e+10    
+      0.08888290739672187
+     -0.01625347486100498
+      0.08946369557655572
+   -3.561174549382201e-05
+    -0.006731182017258544
+      0.08923139516103623
+   -6.967707165516984e-05
+   -3.409966311157184e-05
+     -0.01622614034016565
+      0.08906994307158331
+ 1.07e+10    
+      0.08971433580939131
+     -0.01639673041430468
+      0.09029007084449495
+   -4.172884129796228e-05
+    -0.006793308744684631
+      0.09005587252448553
+   -7.844737273726048e-05
+   -4.018192265296469e-05
+     -0.01636903977161127
+      0.08990292169280353
+ 1.08e+10    
+      0.09054449858884253
+      -0.0165401845587435
+      0.09111552870373595
+   -4.798820793661942e-05
+    -0.006855393044805916
+      0.09087942055851085
+   -8.741714534369347e-05
+   -4.640664615754948e-05
+     -0.01651214408504104
+      0.09073464496697807
+ 1.09e+10    
+      0.09137336704410277
+     -0.01668382514418265
+      0.09194005359933467
+   -5.439155334467866e-05
+    -0.006917430583365272
+      0.09170202312285547
+   -9.658724828204247e-05
+   -5.277562193745566e-05
+     -0.01665544077584646
+      0.09156508391650732
+ 1.1e+10     
+      0.09220091525483623
+     -0.01682764034034906
+      0.09276363221623714
+   -6.094047462234663e-05
+    -0.006979417300864494
+      0.09252366638909633
+   -0.0001059583939922266
+   -5.929052300309269e-05
+     -0.01679891767084096
+      0.09239421232109292
+ 1.11e+10    
+      0.09302711998860402
+       -0.016971618636402
+      0.09358625337999317
+   -6.763645884463822e-05
+    -0.007041349409531336
+      0.09334433874028381
+   -0.0001155311492801029
+   -6.595290783921242e-05
+     -0.01694256292787333
+      0.09322200663512469
+ 1.12e+10    
+      0.09385196061917021
+     -0.01711574884033038
+      0.09440790795932857
+   -7.448088410008712e-05
+    -0.007103223389978685
+       0.0941640306722603
+   -0.0001253059362580503
+   -7.276422142204857e-05
+     -0.01708636503522967
+      0.09404844590614557
+ 1.13e+10    
+      0.09467541904586643
+     -0.01726002007817483
+      0.09522858877060665
+   -8.147502074521806e-05
+     -0.00716503598756589
+      0.09498273469669737
+   -0.0001352830334828952
+    -7.97257964647571e-05
+      -0.0172303128108198
+      0.09487351169441219
+ 1.14e+10    
+      0.09549747961403095
+     -0.01740442179306818
+      0.09604829048420375
+   -8.862003286245188e-05
+    -0.007226784208473439
+      0.09580044524588872
+   -0.0001454625772818671
+   -8.683885487764231e-05
+     -0.01737439540114485
+       0.0956971879935607
+ 1.15e+10    
+      0.09631812903652624
+     -0.01754894374408871
+      0.09686700953281559
+   -9.591697990797229e-05
+    -0.007288465315501499
+      0.09661715857932608
+   -0.0001558445632572889
+   -9.410450942986355e-05
+     -0.01751860228004259
+      0.09651946115238884
+ 1.16e+10    
+      0.09713735631633851
+     -0.01769357600492182
+      0.09768474402171796
+   -0.0001033668185373598
+    -0.007350076823604935
+      0.09743287269208625
+   -0.0001664288479606775
+   -0.0001015237655995404
+     -0.01766292324720811
+      0.09734031979775347
+ 1.17e+10    
+      0.09795515267025946
+     -0.01783830896232539
+      0.09850149364099002
+   -0.0001109704045953043
+    -0.007411616495177372
+      0.09824758722505515
+   -0.0001772151507270247
+   -0.0001090975235986157
+     -0.01780734842648841
+      0.09815975475858578
+ 1.18e+10    
+      0.09877151145364399
+     -0.01798313331439494
+      0.09931725957971145
+    -0.000118728495257953
+    -0.007473082335096649
+      0.09906130337700618
+   -0.0001882030556598336
+   -0.0001168265805600354
+     -0.01795186826394895
+       0.0989777589910186
+ 1.19e+10    
+      0.09958642808623715
+     -0.01812804006862593
+        0.100132044442146
+   -0.0001266417513143117
+    -0.007534472585546072
+      0.09987402381855336
+   -0.0001993920137580347
+   -0.0001247116328739039
+     -0.01809647352571144
+       0.0997943275046172
+ 1.2e+10     
+       0.1003998999790599
+     -0.01827302053976987
+       0.1009458521659099
+   -0.0001347107395750117
+    -0.007595785720624415
+       0.1006857526079935
+   -0.0002107813451756885
+   -0.0001327532786598272
+     -0.01824115529556336
+       0.1006094572897066
+ 1.21e+10    
+        0.101211926462341
+     -0.01841806634748302
+       0.1017586879421342
+   -0.0001429359353965514
+    -0.007657020440759527
+       0.1014964951090505
+    -0.000222370241605362
+   -0.0001409520203635283
+     -0.01838590497233843
+       0.1014231472457779
+ 1.22e+10    
+       0.1020225087144798
+     -0.01856316941376555
+       0.1025705581376175
+    -0.000151317725308462
+    -0.007718175666939469
+       0.1023062579105325
+   -0.0002341577687765524
+   -0.0001493082674645946
+     -0.01853071426706969
+       0.1022353981109627
+ 1.23e+10    
+       0.1028316496920232
+      -0.0187083219601909
+       0.1033814702189722
+   -0.0001598564097329959
+    -0.007779250534776103
+       0.1031150487479112
+   -0.0002461428690606043
+   -0.0001578223392843863
+     -0.01867557519991676
+       0.1030462123925571
+ 1.24e+10    
+         0.10363935406064
+     -0.01885351650492463
+       0.1041914326787581
+   -0.0001685522057851206
+    -0.007840244388415702
+       0.1039228764268285
+   -0.0002583243641732483
+   -0.0001664944678816324
+     -0.01882048009686842
+       0.1038555942985765
+ 1.25e+10    
+       0.1044456281270713
+     -0.01899874585953357
+       0.1050004549636002
+   -0.0001774052501423806
+    -0.007901156774311711
+       0.1047297507485387
+   -0.0002707009579669332
+    -0.000175324801024718
+     -0.01896542158622376
+       0.1046635496703216
+ 1.26e+10    
+       0.1052504797720383
+     -0.01914400312558562
+       0.1058085474042867
+    -0.000186415601974211
+    -0.007961987434874416
+       0.1055356824372869
+     -0.00028327123930421
+   -0.0001843134052296729
+      -0.0191103925948549
+       0.1054700859159366
+ 1.27e+10    
+       0.1060539183840866
+     -0.01928928169104219
+       0.1066157211478376
+   -0.0001955832459200835
+    -0.008022736302012468
+       0.1063406830696269
+   -0.0002960336850046826
+    -0.000193460268853092
+     -0.01925538634425426
+       0.1062752119449353
+ 1.28e+10    
+       0.1068559547943442
+     -0.01943457522644513
+       0.1074219880915367
+    -0.000204908095107356
+    -0.008083403490581108
+       0.1071447650056795
+   -0.0003089866628574046
+   -0.0002027653052297726
+     -0.01940039634637108
+       0.1070789381036754
+ 1.29e+10    
+       0.1076566012121754
+     -0.01957987768090085
+       0.1082273608189189
+   -0.0002143899941982431
+    -0.008143989291752338
+       0.1079479413223314
+   -0.0003221284346913624
+   -0.0002122283558449066
+      -0.0195454163992415
+       0.1078812761117585
+ 1.3e+10     
+       0.1084558711617043
+      -0.0197251832778643
+       0.1090318525376999
+   -0.0002240287224580507
+    -0.008204494166321004
+       0.1087502257483702
+   -0.0003354571594963982
+   -0.0002218491935317701
+     -0.01969044058241687
+       0.1086822389993318
+ 1.31e+10    
+       0.1092537794191917
+     -0.01987048651072724
+        0.109835477019638
+   -0.0002338239968351258
+    -0.008264918737961948
+       0.1095516326015552
+   -0.0003489708965875539
+   -0.0002316275256852495
+     -0.01983546325219611
+        0.109481841045272
+ 1.32e+10    
+       0.1100503419512423
+     -0.02001578213821474
+       0.1106382485423187
+   -0.0002437754750446872
+    -0.008325263786452212
+       0.1103521767276197
+   -0.0003626676088060469
+   -0.0002415629974827568
+     -0.01998047903666824
+       0.1102800977162276
+ 1.33e+10    
+       0.1108455758538236
+     -0.02016106517959396
+       0.1114401818328422
+   -0.0002538827586484778
+    -0.008385530240872243
+       0.1111518734411968
+   -0.0003765451657495615
+     -0.00025165519510422
+     -0.02012548283057046
+       0.1110770256065001
+ 1.34e+10    
+       0.1116394992920762
+     -0.02030633090970124
+       0.1122412920134069
+   -0.0002641453961225824
+    -0.008445719172800348
+       0.1119507384686664
+   -0.0003906013470260229
+   -0.0002619036489430052
+     -0.02027046978996993
+       0.1118726423787423
+ 1.35e+10    
+          0.1124321314409
+     -0.02045157485379341
+       0.1130415945487713
+   -0.0002745628859067795
+    -0.008505831789513252
+       0.1127487878929135
+   -0.0004048338455241809
+   -0.0002723078368004226
+     -0.02041543532677478
+       0.1126669667054551
+ 1.36e+10    
+       0.1132234924262988
+     -0.02059679278222798
+       0.1138411051955763
+   -0.0002851346794283381
+    -0.008565869427206368
+       0.1135460380999894
+   -0.0004192402706949465
+   -0.0002828671870566575
+     -0.02056037510308334
+       0.1134600182112648
+ 1.37e+10    
+       0.1140136032674657
+     -0.02074198070498037
+        0.114639839953518
+   -0.0002958601840941517
+    -0.008625833544246075
+       0.1143425057276685
+   -0.0004338181518377181
+   -0.0002935810818115265
+     -0.02070528502537813
+       0.1142518174159625
+ 1.38e+10    
+       0.1148024858196005
+     -0.02088713486600488
+       0.1154378150183481
+   -0.0003067387662450511
+    -0.008685725714466895
+       0.1151382076158885
+   -0.0004485649413862617
+   -0.0003044488599883979
+     -0.02085016123857405
+       0.1150423856782914
+ 1.39e+10    
+        0.115590162717443
+     -0.02103225173744616
+       0.1162350467366878
+   -0.0003177697540675967
+     -0.00874554762052481
+       0.1159331607590633
+    -0.000463478018188549
+   -0.0003154698203959479
+     -0.02099500011992828
+       0.1158317451404663
+ 1.4e+10     
+       0.1163766573195132
+     -0.02117732801370967
+       0.1170315515626367
+   -0.0003289524404569159
+    -0.008805301047318725
+       0.1167273822602566
+   -0.0004785546907756146
+   -0.0003266432247416651
+     -0.02113979827282106
+       0.1166199186734134
+ 1.41e+10    
+       0.1171619936530499
+      -0.0213223606053994
+        0.117827346016157
+   -0.0003402860858272676
+    -0.008864987875490693
+       0.1175208892872017
+   -0.0004937922006144541
+   -0.0003379683005925241
+     -0.02128455252041676
+       0.1174069298227197
+ 1.42e+10    
+       0.1179461963596422
+     -0.02146734663313137
+       0.1186224466432146
+   -0.0003517699208651162
+    -0.008924610075015677
+        0.118313699030157
+   -0.0005091877253404911
+   -0.0003494442442776502
+     -0.02142925989921429
+       0.1181928027552816
+ 1.43e+10    
+       0.1187292906415474
+     -0.02161228342123171
+       0.1194168699776557
+   -0.0003634031492207595
+    -0.008984169698890709
+       0.1191058286615754
+   -0.0005247383819650575
+   -0.0003610702237289831
+     -0.02157391765249659
+       0.1189775622066473
+ 1.44e+10    
+       0.1195113022086934
+     -0.02175716849132903
+       0.1202106325048006
+   -0.0003751849501355731
+    -0.009043668876932707
+       0.1198972952975768
+   -0.0005404412300538414
+   -0.0003728453812558933
+     -0.02171852322368888
+       0.1197612334290453
+ 1.45e+10    
+       0.1202922572263666
+      -0.0219019995558505
+       0.1210037506267296
+   -0.0003871144810005903
+    -0.009103109809694433
+       0.1206881159612058
+    -0.000556293274872454
+    -0.000384768836249879
+     -0.02186307424963612
+       0.1205438421400972
+ 1.46e+10    
+        0.121072182263585
+     -0.02204677451143154
+       0.1217962406292437
+   -0.0003991908798445991
+    -0.009162494762506378
+       0.1214783075474525
+   -0.0005722914704952347
+   -0.0003968396878166374
+      -0.0220075685538098
+        0.121325414472214
+ 1.47e+10    
+       0.1218511042421623
+      -0.0221914914322497
+       0.1225881186504724
+   -0.0004114132677482214
+    -0.009221826059652825
+       0.1222678867900211
+   -0.0005884327228741801
+   -0.0004090570173320204
+     -0.02215200413945428
+        0.122105976922674
+ 1.48e+10    
+       0.1226290503864668
+     -0.02233614856329302
+       0.1233794006511103
+   -0.0004237807511822325
+    -0.009281106078689412
+       0.1230568702298246
+   -0.0006047138928644761
+   -0.0004214198909197999
+     -0.02229637918268392
+       0.1228855563043883
+ 1.49e+10    
+       0.1234060481738855
+       -0.022480744313573
+       0.1241701023862531
+   -0.0004362924242682124
+    -0.009340337244908292
+       0.1238452741851822
+   -0.0006211317992040333
+   -0.0004339273618487174
+     -0.02244069202554077
+       0.1236641796973561
+ 1.5e+10     
+       0.1241821252860032
+     -0.02262527724929495
+       0.1249602393788144
+   -0.0004489473709594723
+    -0.009399522025958335
+       0.1246331147237013
+   -0.0006376832214438489
+   -0.0004465784728471056
+     -0.02258494116902506
+       0.1244418744008191
+ 1.51e+10    
+       0.1249573095605085
+     -0.02276974608699444
+       0.1257498268944921
+   -0.0004617446671414085
+    -0.009458662926624301
+       0.1254204076358147
+   -0.0006543649028272732
+   -0.0004593722583332007
+     -0.02272912526610806
+       0.1252186678861221
+ 1.52e+10    
+       0.1257316289438411
+     -0.02291414968665321
+       0.1265388799182636
+   -0.0004746833826498363
+    -0.009517762483771626
+       0.1262071684099549
+   -0.0006711735531153133
+   -0.0004723077465602485
+     -0.02287324311473955
+       0.1259945877502924
+ 1.53e+10    
+       0.1265051114445989
+     -0.02305848704480504
+       0.1273274131323792
+   -0.0004877625832066838
+    -0.009576823261460182
+       0.1269934122093331
+   -0.0006881058513563323
+   -0.0004853839616749773
+      -0.0230172936508603
+       0.1267696616703506
+ 1.54e+10    
+       0.1272777850877218
+     -0.02320275728764333
+       0.1281154408958288
+   -0.0005009813322725801
+    -0.009635847846231489
+       0.1277791538503042
+    -0.000705158448598215
+   -0.0004985999256889887
+     -0.02316127594143111
+        0.127543917358367
+ 1.55e+10    
+        0.128049677869473
+     -0.02334695966414237
+       0.1289029772252538
+   -0.0005143386928157143
+    -0.009694838842572488
+        0.128564407782282
+   -0.0007223279705412832
+   -0.0005119546603623952
+     -0.02330518917748947
+       0.1283173825172831
+ 1.56e+10    
+       0.1288208177132417
+     -0.02349109353920367
+       0.1296900357772742
+   -0.0005278337289974613
+    -0.009753798868559002
+       0.1293491880691822
+   -0.0007396110201306019
+   -0.0005254471889994984
+     -0.02344903266724515
+       0.1290900847975149
+ 1.57e+10    
+       0.1295912324261879
+     -0.02363515838683982
+       0.1304766298322051
+   -0.0005414655077741695
+    -0.009812730551680898
+       0.1301335083723612
+   -0.0007570041800867024
+   -0.0005390765381567113
+     -0.02359280582922601
+       0.1298620517543589
+ 1.58e+10    
+       0.1303609496567603
+     -0.02377915378340689
+       0.1312627722791282
+   -0.0005552331004166208
+     -0.00987163652485059
+       0.1309173819350196
+   -0.0007745040153731135
+   -0.0005528417392627093
+     -0.02373650818548451
+       0.1306333108062235
+ 1.59e+10    
+       0.1311299968531075
+       -0.023923079400898
+       0.1320484756022924
+    -0.000569135583946304
+    -0.009930519422596817
+       0.1317008215680423
+   -0.0007921070756007832
+   -0.0005667418301512836
+     -0.02388013935487745
+       0.1314038891937115
+ 1.6e+10     
+        0.131898401222419
+     -0.02406693500030968
+       0.1328337518688111
+    -0.000583172042490735
+    -0.009989381877443547
+       0.1324838396372376
+   -0.0008098098973678544
+   -0.0005807758565077792
+     -0.02402369904642792
+       0.1321738139395741
+ 1.61e+10    
+       0.1326661896912186
+     -0.02421072042509232
+       0.1336186127176232
+   -0.0005973415685575974
+     -0.01004822651647508
+       0.1332664480519484
+   -0.0008276090065350754
+   -0.0005949428732297292
+     -0.02416718705278256
+        0.132943111809569
+ 1.62e+10    
+        0.133433388866645
+     -0.02435443559469717
+         0.13440306934969
+   -0.0006116432642296292
+     -0.01010705595808645
+       0.1340486582549969
+   -0.0008455009204361066
+   -0.0006092419457029482
+     -0.02431060324377297
+       0.1337118092742459
+ 1.63e+10    
+       0.1342000249987511
+     -0.02449808049823055
+       0.1351871325193905
+   -0.0006260762422809715
+     -0.01016587280891922
+       0.1348304812139306
+   -0.0008634821500230097
+   -0.0006236721509938221
+     -0.02445394756009324
+       0.1344799324716906
+ 1.64e+10    
+       0.1349661239438522
+     -0.02464165518822752
+       0.1359708125270873
+   -0.0006406396272168887
+     -0.01022467966098074
+       0.1356119274135339
+   -0.0008815492019466284
+   -0.0006382325789599085
+     -0.02459722000710316
+       0.1352475071712564
+ 1.65e+10    
+       0.1357317111289586
+     -0.02478515977455571
+       0.1367541192128272
+   -0.0006553325562379873
+     -0.01028347908894598
+        0.136393006849569
+   -0.0008996985805723896
+   -0.0006529223332796853
+     -0.02474042064876784
+       0.1360145587383138
+ 1.66e+10    
+       0.1364968115173251
+     -0.02492859441845996
+       0.1375370619511421
+   -0.0006701541801306684
+        -0.01034227364764
+       0.1371737290237094
+   -0.0009179267899318273
+   -0.0006677405324032647
+     -0.02488354960174346
+       0.1367811121000496
+ 1.67e+10    
+       0.1372614495751483
+     -0.02507195932675932
+       0.1383196496469193
+   -0.0006851036640860242
+     -0.01040106586969807
+       0.1379541029396303
+   -0.0009362303356101726
+   -0.0006826863104261467
+     -0.02502660702961904
+       0.1375471917123459
+ 1.68e+10    
+        0.138025649239452
+     -0.02521525474620654
+       0.1391018907323053
+    -0.000700180188448459
+     -0.01045985826340177
+        0.138734137100215
+   -0.0009546057265709508
+   -0.0006977588178875005
+     -0.02516959313732365
+       0.1383128215277735
+ 1.69e+10    
+       0.1387894338871851
+     -0.02535848095801945
+       0.1398837931646076
+    -0.000715382949396235
+     -0.01051865331068732
+       0.1395138395058445
+   -0.0009730494769181592
+   -0.0007129572224951978
+     -0.02531250816570779
+       0.1390780249647264
+ 1.7e+10     
+       0.1395528263055723
+     -0.02550163827259522
+       0.1406653644251606
+   -0.0007307111595562276
+     -0.01057745346532301
+       0.1402932176537253
+   -0.0009915581075970567
+    -0.000728280709779424
+     -0.02545535238630862
+       0.1398428248777344
+ 1.71e+10    
+       0.1403158486637462
+     -0.02564472702441588
+       0.1414466115191234
+   -0.0007461640485546773
+     -0.01063626115125223
+       0.1410722785382227
+    -0.001010128148034435
+   -0.0007437284836775962
+     -0.02559812609630668
+       0.1406072435289822
+ 1.72e+10    
+        0.141078522485693
+     -0.02578774756715467
+       0.1422275409761678
+   -0.0007617408635061113
+     -0.01069507876109809
+       0.1418510286521557
+    -0.001028756137719688
+   -0.0007592997670518358
+     -0.02574082961368243
+       0.1413713025610655
+ 1.73e+10    
+        0.141840868624543
+     -0.02593070026899151
+       0.1430081588520302
+   -0.0007774408694429544
+     -0.01075390865482543
+        0.142629473989018
+    -0.001047438627727666
+   -0.0007749938021424773
+     -0.02588346327258047
+       0.1421350229710155
+ 1.74e+10    
+       0.1426029072382345
+     -0.02607358550814559
+       0.1437884707308829
+   -0.0007932633496877749
+     -0.01081275315855589
+        0.143407620046083
+    -0.001066172182184706
+   -0.0007908098509589144
+      -0.0260260274188884
+         0.14289842508562
+ 1.75e+10    
+       0.1433646577665783
+     -0.02621640366863282
+       0.1445684817284963
+   -0.0008092076061706342
+     -0.01087161456353113
+       0.1441854718283534
+    -0.001084953379679366
+   -0.0008067471956107776
+     -0.02616852240603681
+       0.1436615285380696
+ 1.76e+10    
+        0.144126138909752
+     -0.02635915513625521
+       0.1453481964961553
+   -0.0008252729596936431
+     -0.01093049512522018
+       0.1449630338533184
+    -0.001103778814618904
+   -0.0008228051385817019
+     -0.02631094859102781
+       0.1444243522459557
+ 1.77e+10    
+       0.1448873686082446
+      -0.0265018402948283
+       0.1461276192252906
+   -0.0008414587501454683
+     -0.01098939706256473
+       0.1457403101564761
+    -0.001122645098533384
+   -0.0008389830029480114
+     -0.02645330633069631
+       0.1451869143906455
+ 1.78e+10    
+       0.1456483640242772
+     -0.02664445952265281
+       0.1469067536527967
+   -0.0008577643366674212
+     -0.01104832255735826
+       0.1465173042975826
+    -0.001141548861328781
+    -0.000855280132545112
+     -0.02659559597821056
+       0.1459492323980574
+ 1.79e+10    
+       0.1464091415247185
+      -0.0267870131892358
+       0.1476856030669952
+   -0.0008741890977743059
+     -0.01110727375375338
+       0.1472940193675882
+    -0.001160486752490643
+   -0.0008716958920833079
+     -0.02673781787981578
+       0.1467113229208593
+ 1.8e+10     
+       0.1471697166655137
+     -0.02692950165226574
+       0.1484641703142122
+   -0.0008907324314315207
+     -0.01116625275789161
+       0.1480704579962238
+    -0.001179455442240021
+   -0.0008882296672166508
+     -0.02687997237182595
+       0.1474732018221094
+ 1.81e+10    
+       0.1479301041776425
+     -0.02707192525484581
+       0.1492424578059363
+   -0.0009073937550913445
+       -0.011225261637651
+       0.1488466223601948
+    -0.001198451622643204
+   -0.0009048808645661863
+       -0.027022059777866
+       0.1482348841603562
+ 1.82e+10    
+       0.1486903179546199
+     -0.02721428432298863
+       0.1500204675265184
+   -0.0009241725056901435
+     -0.01128430242250507
+       0.1496225141919476
+    -0.001217472008677024
+   -0.0009216489117006149
+     -0.02716408040636899
+       0.1489963841762161
+ 1.83e+10    
+       0.1494503710415481
+     -0.02735657916337451
+       0.1507982010413847
+   -0.0009410681396092476
+     -0.01134337710348846
+       0.1503981347889689
+    -0.001236513339251298
+   -0.0009385332570766656
+     -0.02730603454832894
+       0.1497577152804369
+ 1.84e+10    
+       0.1502102756257291
+     -0.02749881006137659
+       0.1515756595057254
+    -0.000958080132601345
+     -0.01140248763326264
+       0.1511734850235793
+    -0.001255572378190189
+   -0.0009555333699414279
+     -0.02744792247531223
+        0.150518890043462
+ 1.85e+10    
+       0.1509700430288411
+     -0.02764097727935199
+       0.1523528436736274
+   -0.0009752079796845341
+     -0.01146163592627704
+       0.1519485653531877
+    -0.001274645915174033
+   -0.0009726487401992947
+     -0.02758974443772838
+       0.1512799201865014
+ 1.86e+10    
+       0.1517296837006814
+     -0.02778308105520179
+       0.1531297539076214
+   -0.0009924511950063883
+     -0.01152082385901943
+       0.1527233758309642
+    -0.001293730766643305
+    -0.000989878878245332
+     -0.02773150066335984
+       0.1520408165741129
+ 1.87e+10    
+       0.1524892072144717
+     -0.02792512160119759
+       0.1539063901886031
+    -0.001009809311680006
+     -0.01158005327034966
+       0.1534979161169015
+    -0.001312823776666468
+    -0.001007223314767947
+      -0.0278731913561517
+       0.1528015892082974
+ 1.88e+10    
+       0.1532486222637234
+     -0.02806709910307505
+       0.1546827521261072
+    -0.001027281881593779
+     -0.01163932596191227
+       0.1542721854892254
+    -0.001331921817773074
+    -0.001024681600522337
+     -0.02801481669525984
+       0.1535622472241076
+ 1.89e+10    
+       0.1540079366606528
+     -0.02820901371939232
+       0.1554588389688953
+    -0.001044868475197186
+      -0.0116986436986212
+       0.1550461828561212
+    -0.001351021791753911
+    -0.001042253306077572
+      -0.0281563768343558
+        0.154322798886764
+ 1.9e+10     
+       0.1547671573361356
+     -0.02835086558115047
+       0.1562346496158293
+    -0.001062568681264248
+     -0.01175800820921188
+       0.1558199067677405
+    -0.001370120630429537
+    -0.001059938021538878
+     -0.02829787190118645
+       0.1550832515902724
+ 1.91e+10    
+       0.1555262903411848
+      -0.0284926547916737
+       0.1570101826270025
+    -0.001080382106636618
+     -0.01181742118685522
+       0.1565933554284591
+    -0.001389215296388874
+    -0.001077735356247288
+     -0.02843930199738549
+       0.1558436118575326
+ 1.92e+10    
+       0.1562853408499342
+     -0.02863438142674432
+       0.1577854362350963
+    -0.001098308375947745
+     -0.01187688428982813
+       0.1573665267093493
+       -0.001408302783699
+    -0.001095644938458753
+     -0.02858066719853327
+       0.1566038853419246
+ 1.93e+10    
+       0.1570443131641066
+     -0.02877604553498971
+       0.1585604083569361
+    -0.001116347131330226
+     -0.01193639914223535
+       0.1581394181608366
+    -0.001427380118587755
+    -0.001113666415004357
+      -0.0287219675544606
+       0.1573640768303551
+ 1.94e+10    
+         0.15780321071894
+     -0.02891764713851363
+       0.1593350966052168
+    -0.001134498032107242
+     -0.01199596733477788
+       0.1589120270255106
+    -0.001446444360100424
+    -0.001131799450933515
+     -0.02886320308979192
+       0.1581241902477449
+ 1.95e+10    
+       0.1585620360905455
+     -0.02905918623376821
+       0.1601094983003715
+    -0.001152760754470538
+     -0.01205559042556232
+       0.1596843502510606
+      -0.0014654926007316
+    -0.001150043729141962
+     -0.02900437380472218
+       0.1588842286629332
+ 1.96e+10    
+       0.1593207910046648
+     -0.02920066279265874
+       0.1608836104825572
+    -0.001171134991145409
+     -0.01211526994094747
+       0.1604563845033054
+    -0.001484521967033586
+    -0.001168398949985893
+     -0.02914547967602155
+       0.1596441942959754
+ 1.97e+10    
+       0.1600794763467913
+     -0.02934207676387435
+       0.1616574299237321
+     -0.00118962045104459
+     -0.01217500737642219
+       0.1612281261792896
+    -0.001503529620202231
+    -0.001186864830884366
+       -0.029286520658261
+       0.1604040885268009
+ 1.98e+10    
+       0.1608380921736196
+     -0.02948342807443702
+       0.1624309531397979
+    -0.001208216858912204
+     -0.01223480419751129
+       0.1619995714204226
+     -0.00152251275664147
+      -0.0012054411059106
+     -0.02942749668525236
+        0.161163911905201
+ 1.99e+10    
+       0.1615966377257825
+     -0.02962471663146009
+       0.1632041764027857
+    -0.001226923954958989
+     -0.01229466184070422
+       0.1627707161256295
+    -0.001541468608507301
+    -0.001224127525374393
+     -0.02956840767169383
+       0.1619236641621126
+ 2e+10       
+       0.1623551114418309
+     -0.02976594232410801
+       0.1639770957530593
+    -0.001245741494489691
+     -0.01235458171440271
+       0.1635415559644908
+    -0.001560394444232211
+    -0.001242923855396418
+     -0.02970925351501349
+       0.1626833442221564
+ 2.01e+10    
+       0.1631135109734112
+     -0.02990710502574709
+       0.1647497070115171
+    -0.001264669247524084
+      -0.0124145651998832
+       0.1643120863903489
+    -0.001579287569030724
+    -0.001261829877475931
+     -0.02985003409740169
+       0.1634429502173918
+ 2.02e+10    
+       0.1638718332015933
+     -0.03004820459627773
+       0.1655220057917667
+    -0.001283706998411953
+     -0.01247461365227071
+       0.1650823026533554
+    -0.001598145325387003
+     -0.00128084538805264
+     -0.02999074928802398
+        0.164202479502244
+ 2.03e+10    
+        0.164630074254295
+      -0.0301892408846378
+       0.1662939875122554
+     -0.00130285454544364
+     -0.01253472840151966
+       0.1658521998134392
+    -0.001616965093524788
+    -0.001299970198064425
+     -0.03013139894540297
+       0.1649619286695562
+ 2.04e+10    
+       0.1653882295247556
+     -0.03033021373146665
+       0.1670656474083347
+    -0.001322111700456297
+     -0.01259491075339877
+       0.1666217727531717
+    -0.001635744291860691
+    -0.001319204132501185
+      -0.0302719829199606
+       0.1657212935677198
+ 2.05e+10    
+        0.166146293690996
+     -0.03047112297191733
+       0.1678369805442394
+    -0.001341478288436902
+     -0.01265516199047653
+       0.1673910161905139
+     -0.00165448037744083
+    -0.001338547029956115
+     -0.03041250105671049
+       0.1664805693188327
+ 2.06e+10    
+       0.1669042607362149
+     -0.03061196843860764
+       0.1686079818249661
+    -0.001360954147122903
+     -0.01271548337310411
+       0.1681599246914208
+    -0.001673170846361574
+    -0.001357998742175256
+     -0.03055295319808761
+       0.1672397503378302
+ 2.07e+10    
+       0.1676621239700596
+     -0.03075274996469591
+       0.1693786460080281
+    -0.001380539126600283
+     -0.01277587614039275
+       0.1689284926822895
+    -0.001691813234174645
+    -0.001377559133605708
+     -0.03069333918690713
+       0.1679988303525398
+ 2.08e+10    
+       0.1684198760507125
+     -0.03089346738707172
+       0.1701489677150785
+    -0.001400233088900654
+     -0.01283634151118288
+       0.1696967144622328
+    -0.001710405116276623
+     -0.00139722808094371
+      -0.0308336588694384
+       0.1687578024245971
+ 2.09e+10    
+        0.169177509007731
+     -0.03103412054964724
+       0.1709189414433769
+    -0.001420035907596972
+     -0.01289688068500226
+       0.1704645842151601
+    -0.001728944108283268
+    -0.001417005472682547
+     -0.03097391209858368
+       0.1695166589711693
+ 2.1e+10     
+       0.1699350142655808
+     -0.03117470930673906
+       0.1716885615770937
+    -0.001439947467398565
+      -0.0129574948430111
+       0.1712320960216551
+    -0.001747427866388723
+    -0.001436891208661302
+     -0.03111409873715033
+       0.1702753917874282
+ 2.11e+10    
+       0.1706923826677962
+       -0.031315233526526
+       0.1724578223984304
+    -0.001459967663745972
+     -0.01301818514893127
+        0.171999243870632
+    -0.001765854087709579
+    -0.001456885199614785
+     -0.03125421866120374
+       0.1710339920697115
+ 2.12e+10    
+       0.1714496045017081
+     -0.03145569309457157
+       0.1732267180985491
+    -0.001480096402405524
+     -0.01307895274995841
+       0.1727660216707613
+    -0.001784220510613688
+    -0.001476987366724759
+     -0.03139427176348889
+       0.1717924504393087
+ 2.13e+10    
+       0.1722066695236724
+     -0.03159608791739817
+       0.1739952427882959
+    -0.001500333599064321
+     -0.01313979877765393
+       0.1735324232616482
+    -0.001802524915033951
+    -0.001497197641173275
+      -0.0315342579569096
+        0.172550756966817
+ 2.14e+10    
+        0.172963566984736
+     -0.03173641792610092
+       0.1747633905087073
+     -0.00152067917892535
+     -0.01320072434881656
+       0.1742984424247588
+    -0.001820765122766624
+    -0.001517515963697948
+     -0.03167417717805233
+       0.1733089011969994
+ 2.15e+10    
+       0.1737202856566757
+     -0.03187668307998763
+       0.1755311552412898
+    -0.001541133076303191
+     -0.01326173056633036
+       0.1750640728940788
+    -0.001838938997754094
+    -0.001537942284149585
+     -0.03181402939074304
+       0.1740668721740851
+ 2.16e+10    
+       0.1744768138583488
+     -0.03201688337023389
+       0.1762985309180631
+     -0.00156169523422031
+     -0.01332281851998917
+       0.1758293083664969
+    -0.001857044446351913
+    -0.001558476561052496
+     -0.03195381458962483
+       0.1748246584674506
+ 2.17e+10    
+       0.1752331394822871
+     -0.03215701882354031
+       0.1770655114313577
+    -0.001582365604003888
+     -0.01338398928729539
+       0.1765941425119067
+    -0.001875079417579739
+    -0.001579118761167067
+     -0.03209353280374486
+       0.1755822481976183
+ 2.18e+10    
+       0.1759892500214758
+     -0.03229708950577934
+       0.1778320906433581
+    -0.001603144144883525
+     -0.01344524393423208
+       0.1773585689830181
+     -0.00189304190335588
+    -0.001599868859055416
+      -0.0322331841001389
+       0.1763396290625107
+ 2.19e+10    
+       0.1767451325962548
+     -0.03243709552562171
+       0.1785982623953868
+    -0.001624030823589351
+     -0.01350658351600801
+       0.1781225814248701
+    -0.001910929938715109
+    -0.001620726836649659
+      -0.0323727685874014
+       0.1770967883639013
+ 2.2e+10     
+        0.177500773981279
+     -0.03257703703812902
+       0.1793640205169199
+     -0.00164502561395095
+     -0.01356800907777391
+       0.1788861734840416
+    -0.001928741602009367
+    -0.001641692682822686
+     -0.03251228641922997
+       0.1778537130339987
+ 2.21e+10    
+       0.1782561606324817
+     -0.03271691424830218
+         0.18012935883433
+    -0.001666128496496693
+     -0.01362952165531033
+       0.1796493388175563
+    -0.001946475015090879
+    -0.001662766392961978
+     -0.03265173779793436
+       0.1786103896621049
+ 2.22e+10    
+       0.1790112787139801
+     -0.03285672741457515
+       0.1808942711793509
+    -0.001687339458053641
+     -0.01369112227568549
+       0.1804120711014719
+    -0.001964128343477259
+    -0.001683947968545815
+     -0.03279112297789659
+       0.1793668045212929
+ 2.23e+10    
+       0.1797661141248652
+     -0.03299647685224232
+       0.1816587513972603
+    -0.001708658491347924
+      -0.0137528119578834
+       0.1811743640391578
+    -0.001981699796498296
+    -0.001705237416722162
+     -0.03293044226897505
+       0.1801229435950399
+ 2.24e+10    
+       0.1805206525258271
+      -0.0331361629368109
+       0.1824227933547763
+    -0.001730085594605063
+     -0.01381459171340187
+       0.1819362113692528
+     -0.00199918762742371
+    -0.001726634749889829
+     -0.03306969603983939
+       0.1808787926037674
+ 2.25e+10    
+       0.1812748793655539
+     -0.03327578610726689
+       0.1831863909476649
+    -0.001751620771150847
+     -0.01387646254681973
+       0.1826976068733037
+     -0.00201659013357153
+    -0.001748139985282188
+      -0.0332088847212286
+       0.1816343370312265
+ 2.26e+10    
+       0.1820287799068597
+     -0.03341534686924701
+       0.1839495381080554
+     -0.00177326402901192
+     -0.01393842545633379
+       0.1834585443830827
+    -0.002033905656396708
+    -0.001769753144552662
+     -0.03334800880912223
+       0.1823895621506843
+ 2.27e+10    
+       0.1827823392524894
+      -0.0335548457981067
+       0.1847122288114648
+    -0.001795015380516386
+     -0.01400048143426526
+       0.1842190177875832
+    -0.002051132581559231
+    -0.001791474253362536
+     -0.03348706886781502
+       0.1831444530508507
+ 2.28e+10    
+       0.1835355423705539
+       -0.033694283541876
+       0.1854744570835248
+    -0.001816874841894052
+     -0.01406263146753539
+       0.1849790210396924
+    -0.002068269338971606
+    -0.001813303340970344
+     -0.03362606553288797
+        0.183898994661506
+ 2.29e+10    
+       0.1842883741195502
+     -0.03383366082409589
+       0.1862362170064181
+      -0.0018388424328764
+      -0.0141248765381114
+       0.1857385481625462
+    -0.002085314402824822
+    -0.001835240439822994
+     -0.03376499951406654
+       0.1846531717787758
+ 2.3e+10     
+       0.1850408192729271
+     -0.03397297844652769
+       0.1869975027250161
+     -0.00186091817629583
+     -0.01418721762342177
+         0.18649759325556
+    -0.002102266291592709
+    -0.001857285585148279
+     -0.03390387159795948
+       0.1854069690900134
+ 2.31e+10    
+       0.1857928625431501
+     -0.03411223729172778
+       0.1877583084527246
+    -0.001883102097684263
+     -0.01424965569674266
+       0.1872561505001447
+    -0.002119123568014099
+    -0.001879438814548521
+     -0.03404268265066997
+       0.1861603711982418
+ 2.32e+10    
+       0.1865444886052351
+     -0.03425143832548317
+       0.1885186284770365
+    -0.001905394224871145
+     -0.01431219172755422
+       0.1880142141651042
+    -0.002135884839052225
+    -0.001901700167595567
+     -0.03418143362027368
+       0.1869133626461214
+ 2.33e+10    
+       0.1872956821197121
+     -0.03439058259910052
+       0.1892784571647919
+     -0.00192779458758006
+     -0.01437482668186881
+       0.1887717786117207
+    -0.002152548755831199
+    -0.001924069685426371
+     -0.03432012553915743
+       0.1876659279394005
+ 2.34e+10    
+       0.1880464277549843
+     -0.03452967125154392
+       0.1900377889671492
+    -0.001950303217024689
+      -0.0144375615225308
+       0.1895288382985315
+     -0.00216911401354906
+    -0.001946547410339273
+     -0.03445875952621236
+       0.1884180515698159
+ 2.35e+10    
+       0.1887967102090595
+     -0.03466870551141752
+       0.1907966184242685
+    -0.001972920145503383
+     -0.01450039720948865
+       0.1902853877857963
+    -0.002185579351367014
+    -0.001969133385390915
+     -0.03459733678887732
+       0.1891697180374101
+ 2.36e+10    
+       0.1895465142306181
+     -0.03480768669878808
+       0.1915549401697118
+    -0.001995645405992571
+     -0.01456333470003996
+       0.1910414217396632
+    -0.002201943552274482
+    -0.001991827653993606
+     -0.03473585862502715
+       0.1899209118722322
+ 2.37e+10    
+       0.1902958246393995
+     -0.03494661622684383
+       0.1923127489345613
+    -0.002018479031738692
+     -0.01462637494905049
+       0.1917969349360387
+    -0.002218205442930016
+    -0.002014630259512375
+     -0.03487432642470352
+        0.190671617655402
+ 2.38e+10    
+       0.1910446263458822
+     -0.03508549560338785
+       0.1930700395512604
+    -0.002041421055848898
+     -0.01468951890914727
+        0.192551922264161
+    -0.002234363893477206
+    -0.002037541244862681
+      -0.0350127416716825
+       0.1914218200395008
+ 2.39e+10    
+       0.1917929043702358
+     -0.03522432643216123
+       0.1938268069571812
+    -0.002064471510880191
+     -0.01475276753088707
+       0.1933063787298886
+    -0.002250417817335929
+    -0.002060560652107536
+     -0.03515110594487827
+       0.1921715037682752
+ 2.4e+10     
+       0.1925406438605329
+      -0.0353631104139971
+       0.1945830461979236
+    -0.002087630428427087
+     -0.01481612176290077
+       0.1940602994587027
+    -0.002266366170968429
+    -0.002083688522054778
+     -0.03528942091957928
+       0.1929206536956301
+ 2.41e+10    
+       0.1932878301102012
+     -0.03550184934780087
+       0.1953387524303473
+    -0.002110897838707775
+     -0.01487958255201434
+       0.1948136796984364
+     -0.00228220795362011
+    -0.002106924893853727
+     -0.03542768836851523
+       0.1936692548038915
+ 2.42e+10    
+       0.1940344485747061
+     -0.03564054513135857
+       0.1960939209253482
+    -0.002134273770148795
+     -0.01494315084334782
+        0.195566514821729
+    -0.002297942207035056
+    -0.002130269804591613
+     -0.03556591016275377
+       0.1944172922213264
+ 2.43e+10    
+       0.1947804848874543
+     -0.03577919976197085
+       0.1968485470703757
+    -0.002157758248968108
+     -0.01500682758039225
+       0.1963188003282172
+    -0.002313568015146026
+    -0.002153723288889476
+     -0.03570408827242542
+       0.1951647512389046
+ 2.44e+10    
+       0.1955259248749104
+     -0.03591781533691377
+       0.1976026263717045
+    -0.002181351298756956
+     -0.01507061370506632
+        0.197070531846469
+    -0.002329084503738979
+    -0.002177285378497512
+     -0.03584222476727772
+       0.1959116173262935
+ 2.45e+10    
+       0.1962707545709203
+     -0.03605639405372661
+       0.1983561544564594
+    -0.002205052940060018
+     -0.01513451015775285
+       0.1978217051356626
+    -0.002344490840092148
+     -0.00220095610188994
+     -0.03598032181705601
+       0.1966578761470743
+ 2.46e+10    
+       0.1970149602302386
+     -0.03619493821032709
+        0.199109127074405
+    -0.002228863189954321
+     -0.01519851787731694
+        0.198572316087023
+    -0.002359786232589663
+    -0.002224735483858958
+     -0.03611838169171504
+       0.1974035135731782
+ 2.47e+10    
+       0.1977585283412629
+     -0.03633345020495631
+       0.1998615400995003
+    -0.002252782061627078
+     -0.01526263780110504
+       0.1993223607250167
+    -0.002374969930309705
+    -0.002248623545108691
+     -0.03625640676145825
+       0.1981485156985329
+ 2.48e+10    
+       0.1985014456379685
+     -0.03647193253595509
+       0.2006133895312313
+    -0.002276809563952108
+     -0.01532687086492822
+       0.2000718352083203
+    -0.002390041222587624
+    -0.002272620301847873
+     -0.03639439949661027
+       0.1988928688519246
+ 2.49e+10    
+       0.1992436991110559
+     -0.03661038780137232
+       0.2013646714957191
+    -0.002300945701065356
+     -0.01539121800302786
+       0.2008207358305586
+    -0.002404999438553756
+    -0.002296725765382472
+     -0.03653236246732006
+       0.1996365596090661
+ 2.5e+10     
+       0.1999852760183061
+     -0.03674881869841014
+       0.2021153822466185
+    -0.002325190471939529
+     -0.01545568014802691
+       0.2015690590208306
+    -0.002419843946646457
+    -0.002320939941707722
+     -0.03667029834310076
+       0.2003795748038835
+ 2.51e+10    
+       0.2007261638941593
+      -0.0368872280227075
+       0.2028655181658085
+    -0.002349543869957776
+     -0.01552025823086632
+       0.2023168013440228
+    -0.002434574154100487
+    -0.002345262831099516
+     -0.03680820989220633
+       0.2011219015390182
+ 2.52e+10    
+         0.20146635055852
+     -0.03702561866746476
+       0.2036150757638798
+    -0.002374005882487078
+     -0.01558495318072761
+       0.2030639595009212
+    -0.002449189506410971
+    -0.002369694427705708
+     -0.03694609998084829
+       0.2018635271955506
+ 2.53e+10    
+       0.2022058241247995
+     -0.03716399362241465
+       0.2043640516804326
+    -0.002398576490451024
+     -0.01564976592494315
+       0.2038105303281276
+    -0.002463689486773351
+    -0.002394234719136945
+     -0.03708397157225653
+        0.202604439441959
+ 2.54e+10    
+       0.2029445730072084
+     -0.03730235597264143
+       0.2051124426841834
+    -0.002423255667902358
+     -0.01571469738889401
+        0.204556510797788
+    -0.002478073615499504
+    -0.002418883686057601
+     -0.03722182772558615
+       0.2033446262423122
+ 2.55e+10    
+       0.2036825859273103
+     -0.03744070889725393
+        0.205860245672894
+    -0.002448043381595598
+     -0.01577974849589735
+       0.2053018980171419
+    -0.002492341449410634
+    -0.002443641301776524
+     -0.03735967159467619
+       0.2040840758637174
+ 2.56e+10    
+       0.2044198519198522
+     -0.03757905566791511
+       0.2066074576731243
+    -0.002472939590559714
+     -0.01584492016708291
+       0.2060466892278958
+    -0.002506492581207141
+    -0.002468507531838006
+     -0.03749750642666193
+       0.2048227768830281
+ 2.57e+10    
+       0.2051563603378834
+     -0.03771739964723365
+       0.2073540758398184
+    -0.002497944245671378
+      -0.0159102133212603
+       0.2067908818054322
+    -0.002520526638816005
+    -0.002493482333613108
+     -0.03763533556044593
+       0.2055607181928251
+ 2.58e+10    
+       0.2058921008571858
+     -0.03785574428702331
+       0.2081000974557319
+     -0.00252305728922871
+     -0.01597562887477789
+       0.2075344732578623
+    -0.002534443284716153
+    -0.002518565655891293
+     -0.03777316242503397
+       0.2062978890066911
+ 2.59e+10    
+       0.2066270634800257
+     -0.03799409312643157
+       0.2088455199307014
+    -0.002548278654526022
+     -0.01604116774137335
+       0.2082774612249224
+    -0.002548242215242329
+    -0.002543757438472863
+     -0.03791099053773678
+       0.2070342788637871
+ 2.6e+10     
+       0.2073612385382489
+     -0.03813244978994671
+       0.2095903408007716
+    -0.002573608265429646
+     -0.01610683083201736
+       0.2090198434767308
+    -0.002561923159867878
+    -0.002569057611762357
+      -0.0380488235022463
+       0.2077698776327527
+ 2.61e+10    
+       0.2080946166957367
+      -0.0382708179852851
+        0.210334557727177
+    -0.002599046035955108
+     -0.01617261905475079
+       0.2097616179124053
+    -0.002575485880467165
+    -0.002594466096362623
+     -0.03818666500658865
+       0.2085046755149426
+ 2.62e+10    
+       0.2088271889502444
+     -0.03840920150116564
+       0.2110781684951908
+    -0.002624591869846189
+     -0.01623853331451598
+       0.2105027825585511
+     -0.00258893017055803
+    -0.002619982802670623
+     -0.03832451882096039
+       0.2092386630470244
+ 2.63e+10    
+         0.20955894663464
+     -0.03854760420497709
+        0.211821171012849
+    -0.002650245660155592
+      -0.0163045745129834
+       0.2112433355676236
+    -0.002602255854525013
+    -0.002645607630474417
+     -0.03846238879545224
+       0.2099718311029475
+ 2.64e+10    
+       0.2102898814175646
+     -0.03868603004034191
+       0.2125635633095482
+    -0.002676007288828022
+     -0.01637074354837375
+       0.2119832752161803
+    -0.002615462786823936
+    -0.002671340468551957
+     -0.03860027885766752
+       0.2107041708953145
+ 2.65e+10    
+       0.2110199853035353
+     -0.03882448302458379
+       0.2133053435345326
+    -0.002701876626285746
+     -0.01643704131527613
+       0.2127225999030156
+    -0.002628550851168314
+    -0.002697181194271986
+     -0.03873819301023744
+       0.2114356739761608
+ 2.66e+10    
+        0.211749250632515
+     -0.03896296724610368
+       0.2140465099552663
+    -0.002727853531016868
+     -0.01650346870446317
+       0.2134613081471974
+    -0.002641519959698531
+    -0.002723129673196944
+     -0.03887613532824187
+       0.2121663322371786
+ 2.67e+10    
+       0.2124776700789645
+     -0.03910148686167014
+       0.2147870609557119
+    -0.002753937849166558
+     -0.01657002660270423
+       0.2141993985860071
+    -0.002654370052134196
+    -0.002749185758688313
+     -0.03901410995653994
+       0.2128961379093935
+ 2.68e+10    
+       0.2132052366504049
+      -0.0392400460936286
+       0.2155269950345025
+    -0.002780129414131745
+     -0.01663671589257596
+        0.214936869972786
+    -0.002667101094910457
+    -0.002775349291514953
+     -0.03915212110701469
+        0.213625083562322
+ 2.69e+10    
+       0.2139319436855118
+     -0.03937864922703754
+       0.2162663108030304
+    -0.002806428046159349
+     -0.01670353745227166
+       0.2156737211747001
+    -0.002679713080298991
+    -0.002801620099464131
+     -0.03929017305573968
+       0.2143531621026318
+ 2.7e+10     
+       0.2146577848517567
+     -0.03951730060673329
+       0.2170050069834456
+    -0.002832833551948367
+     -0.01677049215541007
+       0.2164099511704262
+    -0.002692206025514264
+    -0.002827997996955801
+     -0.03942827014007116
+         0.21508036677232
+ 2.71e+10    
+       0.2153827541426268
+     -0.03965600463433289
+       0.2177430824065775
+    -0.002859345724256147
+     -0.01683758087084351
+       0.2171455590477657
+    -0.002704579971805946
+     -0.00285448278466042
+     -0.03956641675567237
+       0.2158066911464413
+ 2.72e+10    
+       0.2161068458744396
+     -0.03979476576517763
+       0.2184805360097825
+    -0.002885964341509108
+     -0.01690480446246638
+       0.2178805440011913
+    -0.002716834983537913
+     -0.00288107424912051
+     -0.03970461735347439
+       0.2165321291303978
+ 2.73e+10    
+        0.216830054682776
+      -0.0399335885052244
+        0.219217366834722
+    -0.002912689167418104
+     -0.01697216378902399
+       0.2186149053293331
+    -0.002728971147254868
+    -0.002907772162376168
+     -0.03984287643658099
+       0.2172566749568202
+ 2.74e+10    
+       0.2175523755185517
+     -0.04007247740788878
+       0.2199535740250782
+    -0.002939519950598895
+     -0.01703965970392282
+       0.2193486424324119
+      -0.0027409885707371
+    -0.002934576281594806
+     -0.03998119855712053
+       0.2179803231820584
+ 2.75e+10    
+       0.2182738036437527
+     -0.04021143707084641
+       0.2206891568242122
+    -0.002966456424197679
+     -0.01710729305504182
+       0.2200817548096152
+    -0.002752887382044143
+    -0.002961486348705472
+     -0.04011958831305089
+       0.2187030686823017
+ 2.76e+10    
+       0.2189943346268484
+     -0.04035047213279656
+        0.221424114572767
+    -0.002993498305522233
+     -0.01717506468454593
+       0.2208142420564381
+    -0.002764667728548128
+    -0.002988502090037834
+     -0.04025805034492455
+       0.2194249066493558
+ 2.77e+10    
+       0.2197139643379154
+     -0.04048958727019433
+       0.2221584467062246
+    -0.003020645295678886
+     -0.01724297542870141
+       0.2215461038619757
+    -0.002776329775957457
+     -0.00301562321596623
+     -0.04039658933261594
+       0.2201458325860906
+ 2.78e+10    
+       0.2204326889434778
+     -0.04062878719395511
+       0.2228921527524185
+    -0.003047897079215233
+     -0.01731102611769427
+       0.2222773400061842
+    -0.002787873707331587
+    -0.003042849420558946
+     -0.04053520999201821
+       0.2208658423015857
+ 2.79e+10    
+       0.2211505049010949
+     -0.04076807664613642
+       0.2236252323290079
+    -0.003075253323769466
+     -0.01737921757545116
+       0.2230079503571115
+    -0.002799299722087649
+    -0.003070180381233023
+      -0.0406739170717137
+       0.2215849319059898
+ 2.8e+10     
+       0.2218674089537128
+     -0.04090746039660296
+       0.2243576851409164
+    -0.003102713679725806
+     -0.01744755061946358
+       0.2237379348680995
+    -0.002810608034999588
+    -0.003097615758414784
+     -0.04081271534962321
+       0.2223030978051189
+ 2.81e+10    
+       0.2225833981237984
+     -0.04104694323967813
+       0.2250895109777418
+    -0.003130277779876915
+      -0.0175160260606158
+       0.2244672935749682
+    -0.002821798875190546
+    -0.003125155195206258
+     -0.04095160962963832
+       0.2230203366948067
+ 2.82e+10    
+       0.2232984697072748
+     -0.04118652999078683
+         0.22582070971114
+    -0.003157945239093132
+     -0.01758464470301637
+       0.2251960265931776
+    -0.002832872485119223
+    -0.003152798317057922
+     -0.04109060473824163
+        0.223736645555034
+ 2.83e+10    
+       0.2240126212672765
+     -0.04132622548309423
+       0.2265512812921847
+    -0.003185715653998854
+     -0.01765340734383359
+       0.2259241341149807
+    -0.002843829119560855
+    -0.003180544731447757
+     -0.04122970552111953
+       0.2244520216438491
+ 2.84e+10    
+       0.2247258506277432
+     -0.04146603456414474
+       0.2272812257487122
+    -0.003213588602656241
+     -0.01772231477313554
+       0.2266516164065628
+    -0.002854669044583641
+    -0.003208394027566954
+     -0.04136891683977188
+       0.2251664624911048
+ 2.85e+10    
+       0.2254381558668679
+     -0.04160596209250402
+       0.2280105431826496
+    -0.003241563644256625
+     -0.01779136777373452
+       0.2273784738051784
+    -0.002865392536521075
+     -0.00323634577601248
+     -0.04150824356812217
+       0.2258799658920204
+ 2.86e+10    
+       0.2261495353104166
+     -0.04174601293441033
+       0.2287392337673335
+    -0.003269640318819285
+      -0.0178605671210359
+       0.2281047067162823
+    -0.002875999880941131
+    -0.003264399528486667
+     -0.04164769058913331
+        0.226592529900599
+ 2.87e+10    
+       0.2268599875249362
+     -0.04188619196043607
+       0.2294672977448187
+    -0.003297818146898622
+     -0.01792991358289196
+       0.2288303156106638
+    -0.002886491371612791
+    -0.003292554817504022
+     -0.04178726279143163
+       0.2273041528229027
+ 2.88e+10    
+       0.2275695113108656
+     -0.04202650404216602
+        0.230194735423188
+    -0.003326096629299046
+     -0.01799940791946127
+       0.2295553010215842
+    -0.002896867309470554
+    -0.003320811156105441
+     -0.04192696506594448
+        0.228014833210215
+ 2.89e+10    
+       0.2282781056955644
+      -0.0421669540488931
+       0.2309215471738546
+    -0.003354475246798197
+     -0.01806905088307242
+       0.2302796635419221
+    -0.002907128001577831
+    -0.003349168037579965
+     -0.04206680230255309
+       0.2287245698520957
+ 2.9e+10     
+        0.228985769926275
+     -0.04230754684433716
+       0.2316477334288733
+    -0.003382953459878688
+     -0.01813884321809378
+       0.2310034038213277
+    -0.002917273760089425
+    -0.003377624935194544
+     -0.04220677938676663
+       0.2294333617693534
+ 2.91e+10    
+       0.2296925034630305
+      -0.0424482872833883
+       0.2323732946782494
+    -0.003411530708468219
+     -0.01820878566080836
+       0.2317265225633931
+    -0.002927304901214242
+    -0.003406181301931259
+     -0.04234690119641865
+       0.2301412082069395
+ 2.92e+10    
+       0.2303983059715229
+     -0.04258918020887958
+       0.2330982314672642
+    -0.003440206411688392
+     -0.01827887893929434
+       0.2324490205228327
+    -0.002937221744178408
+    -0.003434836570233154
+     -0.04248717259838927
+       0.2308481086267882
+ 2.93e+10    
+       0.2311031773159436
+     -0.04273023044838944
+        0.233822544393802
+    -0.003468979967612535
+     -0.01834912377331133
+       0.2331708985026892
+    -0.002947024610189653
+     -0.00346359015175773
+     -0.04262759844535858
+       0.2315540627006073
+ 2.94e+10    
+        0.231807117551808
+     -0.04287144281107978
+       0.2345462341056956
+    -0.003497850753032111
+     -0.01841952087419202
+       0.2338921573515535
+    -0.002956713821403453
+     -0.00349244143713939
+     -0.04276818357259106
+       0.2322590703026404
+ 2.95e+10    
+       0.2325101269187752
+     -0.04301282208456916
+       0.2352693012980868
+    -0.003526818123232412
+     -0.01849007094474036
+        0.234612797960812
+    -0.002966289699891517
+    -0.003521389795759819
+     -0.04290893279475524
+        0.232963131502406
+ 2.96e+10    
+       0.2332122058334758
+     -0.04315437303184575
+        0.235991746710802
+    -0.003555881411777176
+     -0.01856077467913469
+       0.2353328212619155
+    -0.002975752566613325
+    -0.003550434575527278
+     -0.04304985090278168
+       0.2336662465574305
+ 2.97e+10    
+       0.2339133548823574
+      -0.0432961003882219
+        0.236713571125749
+    -0.003585039930302673
+      -0.0186316327628376
+       0.2360522282236796
+    -0.002985102740390945
+    -0.003579575102664526
+     -0.04319094266076088
+       0.2343684159059832
+ 2.98e+10    
+       0.2346135748145532
+     -0.04343800885833115
+       0.2374347753643352
+    -0.003614292968320806
+      -0.0187026458725111
+       0.2367710198496081
+    -0.002994340536888047
+    -0.003608810681505526
+     -0.04333221280288323
+       0.2350696401598241
+ 2.99e+10    
+        0.235312866534793
+     -0.04358010311317245
+       0.2381553602849115
+    -0.003643639793031753
+     -0.01877381467593844
+       0.2374891971752533
+    -0.003003466267593465
+    -0.003638140594301087
+     -0.04347366603042501
+       0.2357699200969789
+ 3e+10       
+       0.2360112310963537
+     -0.04372238778720063
+       0.2388753267802374
+    -0.003673079649145892
+     -0.01884513983195105
+       0.2382067612656034
+    -0.003012480238809734
+    -0.003667564101033487
+     -0.04361530700877973
+       0.2364692566545428
+ 3.01e+10    
+        0.236708669694065
+     -0.04386486747546633
+       0.2395946757749773
+    -0.003702611758715495
+     -0.01891662199036242
+       0.2389237132125077
+    -0.003021382750647269
+    -0.003697080439240157
+     -0.04375714036453929
+         0.23716765092153
+ 3.02e+10    
+       0.2374051836573769
+     -0.04400754673080787
+       0.2403134082232234
+    -0.003732235320975484
+      -0.0189882617919072
+        0.239640054132135
+     -0.00303017409602468
+    -0.003726688823846441
+     -0.04389917068262533
+       0.2378651041317727
+ 3.03e+10    
+       0.2381007744434943
+     -0.04415043006109458
+       0.2410315251060498
+    -0.003761949512194301
+     -0.01906005986818663
+       0.2403557851624695
+    -0.003038854559675516
+    -0.003756388447007692
+     -0.04404140250347265
+       0.2385616176568792
+ 3.04e+10    
+       0.2387954436305865
+     -0.04429352192652491
+       0.2417490274290976
+    -0.003791753485533893
+     -0.01913201684162002
+       0.2410709074608438
+    -0.003047424417162116
+    -0.003786178477960466
+       -0.044183840320267
+       0.2392571929992585
+ 3.05e+10    
+       0.2394891929110764
+     -0.04443682673697869
+       0.2424659162201933
+    -0.003821646370919627
+     -0.01920413332540182
+        0.241785422201513
+    -0.003055883933896917
+    -0.003816058062883014
+     -0.04432648857623758
+       0.2399518317852174
+ 3.06e+10    
+       0.2401820240850206
+     -0.04458034884942815
+       0.2431821925270017
+    -0.003851627274919726
+     -0.01927640992346484
+       0.2424993305732668
+    -0.003064233364171648
+    -0.003846026324765241
+     -0.04446935166200629
+        0.240645535758139
+ 3.07e+10    
+       0.2408739390535771
+     -0.04472409256540381
+       0.2438978574147137
+    -0.003881695280634372
+     -0.01934884723044939
+       0.2432126337770831
+    -0.003072472950194898
+    -0.003876082363287838
+     -0.04461243391299455
+       0.2413383067717443
+ 3.08e+10    
+       0.2415649398125725
+      -0.0448680621285207
+       0.2446129119637691
+    -0.003911849447594504
+     -0.01942144583167761
+       0.2439253330238249
+    -0.003080602921138423
+    -0.003906225254710937
+     -0.04475573960688953
+       0.2420301467834482
+ 3.09e+10    
+       0.2422550284461705
+     -0.04501226172206358
+       0.2453273572676197
+    -0.003942088811670088
+      -0.0194942063031345
+       0.2446374295319784
+    -0.003088623492192692
+    -0.003936454051771983
+     -0.04489927296116976
+       0.2427210578478121
+ 3.1e+10     
+       0.2429442071206465
+     -0.04515669546663262
+       0.2460411944305285
+    -0.003972412384988253
+     -0.01956712921145384
+       0.2453489245254362
+    -0.003096534863631869
+    -0.003966767783593244
+     -0.04504303813069144
+       0.2434110421100928
+ 3.11e+10    
+       0.2436324780782705
+      -0.0453013674178494
+       0.2467544245654071
+    -0.004002819155860896
+      -0.0196402151139099
+       0.2460598192313223
+    -0.003104337219888856
+    -0.003997165455598474
+     -0.04518703920533672
+       0.2441001017999054
+ 3.12e+10    
+       0.2443198436313054
+     -0.04544628156412577
+       0.2474670487916941
+     -0.00403330808872196
+     -0.01971346455841495
+       0.2467701148778642
+    -0.003112030728640626
+    -0.004027646049439084
+     -0.04533128020772361
+       0.2447882392249871
+ 3.13e+10    
+       0.2450063061561173
+      -0.0455914418244931
+        0.248179068233274
+     -0.00406387812407402
+     -0.01978687808352178
+       0.2474798126923083
+    -0.003119615539904208
+    -0.004058208522929719
+     -0.04547576509097932
+       0.2454754567650818
+ 3.14e+10    
+       0.2456918680874085
+      -0.0457368520464956
+       0.2488904840164372
+    -0.004094528178444783
+     -0.01986045621843214
+       0.2481889138988822
+    -0.003127091785143735
+    -0.004088851809993112
+      -0.0456204977365765
+       0.2461617568659352
+ 3.15e+10    
+       0.2463765319125681
+     -0.04588251600414556
+       0.2496012972678776
+    -0.004125257144352737
+     -0.01993419948300983
+       0.2488974197168021
+    -0.003134459576388846
+    -0.004119574820614301
+     -0.04576548195223339
+        0.246847142033413
+ 3.16e+10    
+       0.2470603001661484
+     -0.04602843739594244
+       0.2503115091127386
+    -0.004156063890282417
+     -0.02000810838779953
+        0.249605331358327
+    -0.003141719005364802
+    -0.004150376440804199
+     -0.04591072146987819
+       0.2475316148277384
+ 3.17e+10    
+       0.2477431754244631
+     -0.04617461984295469
+       0.2510211206726953
+    -0.004186947260668875
+      -0.0200821834340503
+       0.2503126500268578
+    -0.003148870142634614
+    -0.004181255532572332
+     -0.04605621994367761
+       0.2482151778578554
+ 3.18e+10    
+       0.2484251603003144
+     -0.04632106688696527
+        0.251730133064083
+    -0.004217906075891659
+     -0.02015642511374426
+       0.2510193769150864
+    -0.003155913036753494
+    -0.004212210933908885
+     -0.04620198094813007
+       0.2488978337759161
+ 3.19e+10    
+       0.2491062574378463
+     -0.04646778198868139
+       0.2524385473960658
+    -0.004248939132277885
+     -0.02023083390963028
+       0.2517255132031868
+    -0.003162847713436021
+    -0.004243241458775837
+     -0.04634800797622388
+       0.2495795852718982
+ 3.2e+10     
+       0.2497864695075254
+     -0.04661476852600719
+       0.2531463647688524
+    -0.004280045202114475
+     -0.02030541029526245
+       0.2524310600570587
+    -0.003169674174736095
+    -0.004274345897107285
+     -0.04649430443765974
+       0.2502604350683475
+ 3.21e+10    
+       0.2504657992012526
+      -0.0467620297923795
+       0.2538535862719487
+     -0.00431122303366979
+     -0.02038015473504242
+       0.2531360186266107
+    -0.003176392398240203
+    -0.004305523014818905
+     -0.04664087365713797
+       0.2509403859152539
+ 3.22e+10    
+       0.2511442492276027
+     -0.04690956899516881
+       0.2545602129824613
+    -0.004342471351223862
+     -0.02045506768426794
+       0.2538403900440996
+    -0.003183002336274147
+    -0.004336771553826115
+     -0.04678771887271152
+       0.2516194405850563
+ 3.23e+10    
+       0.2518218223071951
+     -0.04705738925414121
+       0.2552662459634377
+    -0.004373788855107812
+     -0.02053014958918418
+       0.2545441754225064
+    -0.003189503915123551
+    -0.004368090232071577
+     -0.04693484323420152
+       0.2522976018677785
+ 3.24e+10    
+       0.2524985211681944
+      -0.0472054935999856
+       0.2559716862622548
+    -0.004405174221752314
+     -0.02060540088704037
+       0.2552473758539673
+    -0.003195897034268291
+    -0.004399477743561246
+     -0.04708224980167938
+       0.2529748725662989
+ 3.25e+10    
+       0.2531743485419386
+     -0.04735388497290195
+       0.2566765349090472
+    -0.004436626103744444
+     -0.02068082200615037
+       0.2559499924082461
+    -0.003202181565631275
+    -0.004430932758409369
+     -0.04722994154401149
+       0.2536512554917489
+ 3.26e+10    
+       0.2538493071587007
+     -0.04750256622125328
+        0.257380792915183
+    -0.004468143129893445
+     -0.02075641336595747
+       0.2566520261312559
+    -0.003208357352841679
+    -0.004462453922892122
+     -0.04737792133746876
+       0.2543267534590457
+ 3.27e+10    
+        0.254523399743575
+     -0.04765154010027887
+       0.2580844612717784
+    -0.004499723905305134
+     -0.02083217537710295
+        0.257353478043624
+    -0.003214424210512997
+    -0.004494039859509857
+     -0.04752619196439894
+       0.2550013692825559
+ 3.28e+10    
+       0.2551966290124956
+     -0.04780080927087021
+       0.2587875409482587
+    -0.004531367011464667
+     -0.02090810844149859
+        0.258054349139306
+    -0.003220381923535905
+    -0.004525689167057987
+     -0.04767475611196291
+       0.2556751057718895
+ 3.29e+10    
+       0.2558689976683799
+     -0.04795037629840761
+        0.259490032890963
+    -0.004563071006327682
+     -0.02098421295240332
+       0.2587546403842434
+    -0.003226230246386502
+    -0.004557400420706272
+     -0.04782361637093314
+       0.2563479657278271
+ 3.3e+10     
+       0.2565405083974009
+     -0.04810024365165774
+       0.2601919380217871
+    -0.004594834424419912
+     -0.02106048929450262
+       0.2594543527150649
+    -0.003231968902449805
+     -0.00458917217208632
+     -0.04797277523455461
+       0.2570199519383721
+ 3.31e+10    
+       0.2572111638653835
+     -0.04825041370173185
+        0.260893257236875
+    -0.004626655776944837
+     -0.02113693784399241
+        0.260153487037838
+    -0.003237597583358971
+    -0.004621002949387545
+     -0.04812223509746814
+       0.2576910671749382
+ 3.32e+10    
+        0.257880966714326
+     -0.04840088872110377
+       0.2615939914053498
+    -0.004658533551899279
+     -0.02121355896866582
+         0.26085204422686
+    -0.003243115948350236
+    -0.004652891257461213
+     -0.04827199825469403
+       0.2583613141886598
+ 3.33e+10    
+       0.2585499195590467
+     -0.04855167088268737
+       0.2622941413680856
+    -0.004690466214197351
+     -0.02129035302800287
+       0.2615500251234942
+    -0.003248523623633977
+     -0.00468483557793249
+     -0.04842206690067752
+       0.2590306957068333
+ 3.34e+10    
+       0.2592180249839487
+     -0.04870276225897231
+       0.2629937079365244
+    -0.004722452205801769
+     -0.02136732037326412
+       0.2622474305350526
+    -0.003253820201781854
+    -0.004716834369320549
+     -0.04857244312839386
+       0.2596992144294817
+ 3.35e+10    
+       0.2598852855399109
+      -0.0488541648212186
+       0.2636926918915332
+    -0.004754489945863373
+     -0.02144446134758674
+       0.2629442612337194
+    -0.003259005241130452
+    -0.004748886067166306
+     -0.04872312892851315
+        0.260366873026043
+ 3.36e+10    
+       0.2605517037412903
+     -0.04900588043870796
+       0.2643910939823014
+    -0.004786577830867724
+     -0.02152177628608352
+       0.2636405179555177
+    -0.003264078265201448
+    -0.004780989084168229
+     -0.04887412618862424
+       0.2610336741321863
+ 3.37e+10    
+       0.2612172820630508
+     -0.04915791087805297
+       0.2650889149252803
+    -0.004818714234789796
+     -0.02159926551594493
+       0.2643362013993201
+    -0.003269038762138495
+    -0.004813141810325402
+     -0.04902543669251709
+       0.2616996203467439
+ 3.38e+10    
+       0.2618820229380013
+     -0.04931025780256183
+       0.2657861554031637
+    -0.004850897509255508
+     -0.02167692935654345
+       0.2650313122258991
+    -0.003273886184161053
+    -0.004845342613088433
+     -0.04917706211952222
+       0.2623647142287659
+ 3.39e+10    
+       0.2625459287541508
+     -0.04946292277165849
+       0.2664828160639068
+    -0.004883125983710835
+     -0.02175476811954076
+       0.2657258510570227
+    -0.003278619947035322
+    -0.004877589837517404
+     -0.04932900404390837
+       0.2630289582946951
+ 3.4e+10     
+       0.2632090018521734
+     -0.04961590724035838
+       0.2671788975197865
+    -0.004915397965597906
+     -0.02183278210899699
+       0.2664198184745852
+    -0.003283239429562296
+    -0.004909881806447433
+      -0.0494812639343348
+       0.2636923550156533
+ 3.41e+10    
+        0.263871244522988
+     -0.04976921255879763
+       0.2678744003465012
+    -0.004947711740538133
+     -0.02191097162148288
+       0.2671132150197856
+    -0.003287743973083402
+    -0.004942216820661196
+     -0.04963384315336076
+       0.2643549068148487
+ 3.42e+10    
+       0.2645326590054436
+     -0.04992283997181619
+       0.2685693250823068
+    -0.004980065572522178
+     -0.02198933694619301
+       0.2678060411923402
+    -0.003292132881003526
+    -0.004974593159068423
+     -0.04978674295700916
+       0.2650166160650924
+ 3.43e+10    
+       0.2651932474841111
+     -0.05007679061859329
+       0.2692636722271959
+    -0.005012457704106761
+     -0.02206787836506222
+       0.2684982974497364
+    -0.003296405418331716
+    -0.005007009078892587
+     -0.04993996449438361
+       0.2656774850864256
+ 3.44e+10    
+       0.2658530120871823
+     -0.05023106553233535
+       0.2699574422421114
+    -0.005044886356617912
+     -0.02214659615288347
+        0.269189984206528
+    -0.003300560811239859
+    -0.005039462815864097
+     -0.05009350880734011
+       0.2663375161438595
+ 3.45e+10    
+         0.26651195488447
+     -0.05038566564001427
+       0.2706506355481973
+    -0.005077349730360921
+      -0.0222254905774272
+       0.2698811018336648
+    -0.003304598246639221
+    -0.005071952584420203
+     -0.05024737683021054
+       0.2669967114452186
+ 3.46e+10    
+       0.2671700778855102
+     -0.05054059176215718
+       0.2713432525260894
+     -0.00510984600483651
+      -0.0223045618995628
+       0.2705716506578629
+    -0.003308516871775068
+    -0.005104476577911625
+     -0.05040156938957824
+       0.2676550731390931
+ 3.47e+10    
+       0.2678273830377618
+     -0.05069584461268543
+       0.2720352935152416
+    -0.005142373338963173
+     -0.02238381037338186
+        0.271261630961012
+    -0.003312315793839581
+    -0.005137032968815299
+     -0.05055608720410455
+       0.2683126033128909
+ 3.48e+10    
+       0.2684838722249049
+     -0.05085142479880201
+       0.2727267588132866
+    -0.005174929871305718
+     -0.02246323624632197
+        0.271951042979615
+    -0.003315994079603151
+    -0.005169619908953796
+      -0.0507109308844049
+        0.268969303990994
+ 3.49e+10    
+       0.2691395472652338
+     -0.05100733282092843
+       0.2734176486754353
+    -0.005207513720309812
+     -0.02254283975929326
+       0.2726398869042735
+    -0.003319550755064036
+    -0.005202235529720376
+     -0.05086610093297638
+       0.2696251771330129
+ 3.5e+10     
+       0.2697944099101417
+     -0.05116356907268769
+       0.2741079633139073
+    -0.005240122984542181
+     -0.02262262114680455
+       0.2733281628791969
+    -0.003322984805116746
+    -0.005234877942310569
+     -0.05102159774417089
+       0.2702802246321372
+ 3.51e+10    
+       0.2704484618426969
+     -0.05132013384093429
+       0.2747977028974008
+    -0.005272755742936622
+     -0.02270258063709238
+       0.2740158710017566
+    -0.003326295173239038
+    -0.005267545237959376
+     -0.05117742160421938
+        0.270934448313584
+ 3.52e+10    
+       0.2711017046763102
+     -0.05147702730583049
+       0.2754868675505913
+    -0.005305410055045599
+     -0.02278271845224931
+       0.2747030113220674
+    -0.003329480761197833
+    -0.005300235488184242
+     -0.05133357269130075
+       0.2715878499331376
+ 3.53e+10    
+       0.2717541399534847
+     -0.05163424954096744
+       0.2761754573536705
+    -0.005338083961297092
+      -0.0228630348083549
+        0.275389583842607
+    -0.003332540428773957
+    -0.005332946745033786
+     -0.05149005107565811
+         0.27224043117578
+ 3.54e+10    
+       0.2724057691446544
+     -0.05179180051352967
+       0.2768634723419107
+    -0.005370775483257007
+     -0.02294352991560588
+       0.2760755885178681
+    -0.003335472993505997
+    -0.005365677041341867
+     -0.05164685671976015
+       0.2728921936544112
+ 3.55e+10    
+       0.2730565936471049
+     -0.05194968008450514
+       0.2775509125052694
+    -0.005403482623896427
+     -0.02302420397844848
+       0.2767610252540404
+    -0.003338277230453293
+    -0.005398424390987209
+     -0.05180398947850736
+       0.2735431389086574
+ 3.56e+10    
+       0.2737066147839715
+     -0.05210788800893525
+       0.2782377777880182
+    -0.005436203367864193
+     -0.02310505719571009
+       0.2774458939087279
+    -0.003340951871978086
+    -0.005431186789158108
+     -0.05196144909948181
+       0.2741932684037623
+ 3.57e+10    
+       0.2743558338033234
+     -0.05226642393620921
+       0.2789240680884099
+    -0.005468935681764187
+     -0.02318608976073258
+       0.2781301942906974
+    -0.003343495607547097
+    -0.005463962212622256
+     -0.05211923522324026
+       0.2748425835295622
+ 3.58e+10    
+       0.2750042518773172
+     -0.05242528741039858
+       0.2796097832583734
+    -0.005501677514437291
+      -0.0232673018615052
+       0.2788139261596551
+    -0.003345907083552441
+    -0.005496748620001655
+     -0.05227734738364967
+       0.2754910855995431
+ 3.59e+10    
+       0.2756518701014307
+     -0.05258447787063197
+       0.2802949231032389
+    -0.005534426797248227
+     -0.02334869368079837
+       0.2794970892260571
+    -0.003348184903152103
+    -0.005529543952052223
+      -0.0524357850082631
+       0.2761387758499733
+ 3.6e+10     
+       0.2762986894937662
+     -0.05274399465150933
+       0.2809794873814939
+    -0.005567181444376746
+     -0.02343026539629728
+       0.2801796831509473
+    -0.003350327626129938
+    -0.005562346131948269
+     -0.05259454741873777
+       0.2767856554391181
+ 3.61e+10    
+       0.2769447109944301
+     -0.05290383698355648
+       0.2816634758045692
+    -0.005599939353112983
+     -0.02351201718073604
+       0.2808617075458245
+    -0.003352333768775475
+    -0.005595153065571318
+     -0.05275363383129168
+       0.2774317254465246
+ 3.62e+10    
+       0.2775899354649747
+     -0.05306400399371541
+       0.2823468880366515
+    -0.005632698404157387
+     -0.02359394920203166
+       0.2815431619725412
+    -0.003354201803783268
+    -0.005627962641803604
+     -0.05291304335720037
+       0.2780769868723824
+ 3.63e+10    
+       0.2782343636879146
+     -0.05322449470587409
+       0.2830297236945265
+    -0.005665456461924435
+     -0.02367606162341797
+       0.2822240459432262
+    -0.003355930160172274
+    -0.005660772732825678
+     -0.05307277500333124
+       0.2787214406369542
+ 3.64e+10    
+       0.2788779963663031
+     -0.05338530804143134
+       0.2837119823474504
+    -0.005698211374850478
+     -0.02375835460357945
+       0.2829043589202365
+    -0.003357517223224951
+    -0.005693581194418477
+     -0.05323282767271498
+       0.2793650875800766
+ 3.65e+10    
+       0.2795208341233765
+     -0.05354644281989853
+       0.2843936635170457
+    -0.005730960975705273
+     -0.02384082829678535
+       0.2835841003161383
+    -0.003358961334446471
+    -0.005726385866268967
+     -0.05339320016515539
+       0.2800079284607263
+ 3.66e+10    
+       0.2801628775022584
+     -0.05370789775953582
+       0.2850747666772267
+    -0.005763703081907334
+     -0.02392348285302254
+       0.2842632694937103
+     -0.00336026079154382
+    -0.005759184572280238
+     -0.05355389117787332
+       0.2806499639566537
+ 3.67e+10    
+       0.2808041269657256
+     -0.05386967147802303
+       0.2857552912541499
+    -0.005796435495842665
+     -0.02400631841812892
+       0.2849418657659759
+    -0.003361413848425124
+     -0.00579197512088492
+     -0.05371489930618706
+       0.2812911946640809
+ 3.68e+10    
+       0.2814445828960295
+     -0.05403176249316353
+       0.2864352366261905
+     -0.00582915600518715
+     -0.02408933513392613
+       0.2856198883962608
+    -0.003362418715218962
+    -0.005824755305362608
+     -0.05387622304422663
+       0.2819316210974579
+ 3.69e+10    
+       0.2820842455947797
+      -0.0541941692236226
+       0.2871146021239457
+    -0.005861862383231891
+     -0.02417253313835154
+       0.2862973365982724
+     -0.00336327355831403
+    -0.005857522904160528
+     -0.05403786078568157
+        0.282571243689282
+ 3.7e+10     
+        0.282723115282879
+     -0.05435688998969591
+        0.287793387030258
+    -0.005894552389212194
+     -0.02425591256558978
+       0.2869742095362073
+    -0.003363976500418942
+    -0.005890275681217739
+     -0.05419981082458257
+       0.2832100627899757
+ 3.71e+10    
+       0.2833611921005117
+     -0.05451992301411059
+       0.2884715905802699
+     -0.00592722376863898
+     -0.02433947354620389
+       0.2876505063248788
+    -0.003364525620642381
+    -0.005923011386292622
+     -0.05436207135611408
+       0.2838480786678184
+ 3.72e+10    
+        0.283998476107187
+      -0.0546832664228576
+       0.2891492119614963
+    -0.005959874253633731
+     -0.02442321620726538
+       0.2883262260298717
+    -0.003364918954593586
+     -0.00595572775529336
+     -0.05452464047745984
+       0.2844852915089366
+ 3.73e+10    
+         0.28463496728183
+     -0.05484691824605255
+       0.2898262503139226
+    -0.005992501563265632
+     -0.02450714067248374
+       0.2890013676677154
+    -0.003365154494503225
+    -0.005988422510611505
+     -0.05468751618867777
+       0.2851217014173448
+ 3.74e+10    
+       0.2852706655229232
+      -0.0550108764188276
+       0.2905027047301265
+    -0.006025103403891749
+     -0.02459124706233487
+       0.2896759302060825
+     -0.00336523018936467
+    -0.006021093361458485
+     -0.05485069639360585
+       0.2857573084150392
+ 3.75e+10    
+       0.2859055706486939
+     -0.05517513878225085
+       0.2911785742554197
+     -0.00605767746949957
+     -0.02467553549418912
+       0.2903499125640074
+    -0.003365143945095737
+     -0.00605373800420466
+     -0.05501417890079693
+       0.2863921124421412
+ 3.76e+10    
+       0.2865396823973499
+     -0.05533970308427418
+       0.2918538578880147
+    -0.006090221442052028
+     -0.02476000608243763
+       0.2910233136121265
+    -0.003364893624720861
+    -0.006086354122721283
+     -0.05517796142448245
+       0.2870261133570909
+ 3.77e+10    
+       0.2871730004273573
+     -0.05550456698070848
+       0.2925285545792087
+    -0.006122732991834498
+     -0.02484465893861821
+       0.2916961321729389
+    -0.003364477048573906
+    -0.006118939388724553
+     -0.05534204158556355
+       0.2876593109368832
+ 3.78e+10    
+       0.2878055243177615
+     -0.05566972803622521
+       0.2932026632335931
+    -0.006155209777804444
+     -0.02492949417154007
+       0.2923683670210881
+    -0.003363891994521335
+    -0.006151491462122481
+     -0.05550641691263047
+       0.2882917048773559
+ 3.79e+10    
+       0.2884372535685524
+     -0.05583518372538453
+       0.2938761827092796
+    -0.006187649447942591
+     -0.02501451188740699
+       0.2930400168836608
+    -0.003363136198206072
+    -0.006184007991363693
+     -0.05567108484300706
+       0.2889232947935165
+ 3.8e+10     
+       0.2890681876010666
+     -0.05600093143368819
+       0.2945491118181475
+    -0.006220049639606249
+     -0.02509971218993996
+       0.2937110804405105
+    -0.003362207353311826
+    -0.006216486613788366
+     -0.05583604272382266
+       0.2895540802199135
+ 3.81e+10    
+       0.2896983257584296
+     -0.05616696845865696
+       0.2952214493261121
+    -0.006252407979884353
+     -0.02518509518049809
+       0.2943815563245922
+    -0.003361103111848069
+    -0.006248924955981358
+     -0.05600128781310824
+       0.2901840606110509
+ 3.82e+10    
+       0.2903276673060377
+     -0.05633329201093359
+       0.2958931939534104
+    -0.006284722085954065
+     -0.02527066095819827
+       0.2950514431223205
+    -0.003359821084455554
+    -0.006281320634126985
+     -0.05616681728091727
+       0.2908132353418378
+ 3.83e+10    
+       0.2909562114320723
+     -0.05649989921540668
+       0.2965643443749041
+    -0.006316989565439115
+     -0.02535640962003385
+       0.2957207393739461
+    -0.003358358840732417
+    -0.006313671254365669
+     -0.05633262821047104
+       0.2914416037080825
+ 3.84e+10    
+       0.2915839572480527
+     -0.05666678711235996
+       0.2972348992204049
+    -0.006349208016769243
+     -0.02544234126099151
+       0.2963894435739455
+    -0.003356713909580842
+    -0.006345974413152163
+     -0.05649871759932613
+       0.2920691649270168
+ 3.85e+10    
+       0.2922109037894219
+     -0.05683395265864184
+       0.2979048570750135
+    -0.006381375029541226
+     -0.02552845597416699
+        0.297057554171431
+    -0.003354883779574379
+    -0.006378227697615377
+      -0.0566650823605661
+       0.2926959181378642
+ 3.86e+10    
+       0.2928370500161636
+     -0.05700139272885775
+       0.2985742164794777
+    -0.006413488184880818
+     -0.02561475385087939
+       0.2977250695705768
+    -0.003352865899345785
+    -0.006410428685919314
+     -0.05683171932401376
+       0.2933218624024349
+ 3.87e+10    
+       0.2934623948134522
+     -0.05716910411658241
+       0.2992429759305674
+    -0.006445545055806004
+      -0.0257012349807835
+       0.2983919881310586
+    -0.003350657677995343
+    -0.006442574947625785
+     -0.05699862523746527
+       0.2939469967057602
+ 3.88e+10    
+       0.2940869369923348
+     -0.05733708353559364
+       0.2999111338814659
+    -0.006477543207590915
+     -0.02578789945198149
+       0.2990583081685133
+     -0.00334825648551991
+     -0.00647466404405769
+     -0.05716579676794562
+       0.2945713199567561
+ 3.89e+10    
+        0.294710675290436
+     -0.05750532762112477
+       0.3005786887421761
+     -0.00650948019813072
+     -0.02587474735113217
+       0.2997240279550097
+    -0.003345659653262222
+    -0.006506693528663784
+     -0.05733323050298324
+       0.2951948309889181
+ 3.9e+10     
+       0.2953336083727006
+     -0.05767383293113714
+       0.3012456388799451
+    -0.006541353578307262
+     -0.02596177876355893
+       0.3003891457195346
+    -0.003342864474380993
+    -0.006538660947384129
+     -0.05750092295190491
+       0.2958175285610476
+ 3.91e+10    
+       0.2959557348321549
+     -0.05784259594761063
+       0.3019119826196995
+    -0.006573160892355108
+     -0.02604899377335625
+       0.3010536596484962
+    -0.003339868204341182
+    -0.006570563839016386
+     -0.05766887054714916
+       0.2964394113580045
+ 3.92e+10    
+       0.2965770531906987
+     -0.05801161307785281
+       0.3025777182445015
+    -0.006604899678228313
+     -0.02613639246349456
+       0.3017175678862397
+    -0.003336668061424812
+    -0.006602399735582867
+     -0.05783706964559893
+       0.2970604779914905
+ 3.93e+10    
+       0.2971975618999209
+     -0.05818088065582458
+       0.3032428439960129
+    -0.006636567467967237
+     -0.02622397491592283
+        0.302380868535573
+    -0.003333261227262292
+    -0.006634166162698156
+     -0.05800551652993005
+       0.2976807270008558
+ 3.94e+10    
+       0.2978172593419404
+     -0.05835039494348454
+       0.3039073580749788
+    -0.006668161788066039
+     -0.02631174121167017
+        0.303043559658312
+    -0.003329644847383763
+    -0.006665860639937179
+     -0.05817420740997942
+        0.298300156853935
+ 3.95e+10    
+       0.2984361438302676
+     -0.05852015213214728
+       0.3045712586417211
+    -0.006699680159839946
+     -0.02639969143094545
+        0.303705639275835
+    -0.003325816031791037
+    -0.006697480681203471
+     -0.05834313842412845
+       0.2989187659479042
+ 3.96e+10    
+       0.2990542136106924
+     -0.05869014834385966
+       0.3052345438166467
+    -0.006731120099792726
+     -0.02648782565323483
+       0.3043671053696489
+    -0.003321771855549644
+    -0.006729023795098016
+     -0.05851230564070228
+       0.2995365526101639
+ 3.97e+10    
+       0.2996714668621884
+     -0.05886037963279148
+       0.3058972116807697
+       -0.006762479119984
+       -0.026576143957398
+       0.3050279558819687
+    -0.003317509359400988
+    -0.006760487485288052
+     -0.05868170505938547
+       0.3001535150992449
+ 3.98e+10    
+       0.3002879016978422
+     -0.05903084198664051
+       0.3065592602762435
+    -0.006793754728396649
+     -0.02666464642176242
+       0.3056881887163087
+    -0.003313025550394717
+    -0.006791869250875781
+     -0.05885133261265217
+       0.3007696516057325
+ 3.99e+10    
+       0.3009035161657995
+     -0.05920153132805277
+        0.307220687606907
+    -0.006824944429303577
+     -0.02675333312421557
+       0.3063478017380848
+    -0.003308317402541101
+    -0.006823166586767217
+     -0.05902118416721081
+       0.3013849602532168
+ 4e+10       
+       0.3015183082502316
+     -0.05937244351605554
+        0.307881491638842
+    -0.006856045723634395
+     -0.02684220414229556
+       0.3070067927752278
+    -0.003303381857483309
+    -0.006854376984040884
+     -0.05919125552546282
+       0.3019994390992594
+ 4.01e+10    
+       0.3021322758723183
+     -0.05954357434750461
+       0.3085416703009428
+    -0.006887056109341267
+     -0.02693125955328014
+       0.3076651596188062
+    -0.003298215825189707
+    -0.006885497930315848
+      -0.0593615424269746
+       0.3026130861363778
+ 4.02e+10    
+       0.3027454168912486
+     -0.05971491955854254
+       0.3092012214854943
+    -0.006917973081764802
+     -0.02702049943427304
+        0.308322900023661
+    -0.003292816184665768
+    -0.006916526910119944
+     -0.05953204054996225
+        0.303225899293053
+ 4.03e+10    
+       0.3033577291052392
+     -0.05988647482607172
+        0.309860143048766
+    -0.006948794133998432
+     -0.02710992386228956
+       0.3089800117090487
+    -0.003287179784685912
+    -0.006947461405257123
+     -0.05970274551278909
+       0.3038378764347518
+ 4.04e+10    
+       0.3039692102525665
+     -0.06005823576923636
+       0.3105184328116086
+    -0.006979516757252771
+     -0.02719953291433932
+       0.3096364923592963
+    -0.003281303444544747
+    -0.006978298895174187
+     -0.05987365287547494
+       0.3044490153649631
+ 4.05e+10    
+       0.3045798580126147
+     -0.06023019795091761
+       0.3111760885600693
+    -0.007010138441218567
+     -0.02728932666750765
+       0.3102923396244613
+    -0.003275183954827986
+    -0.007009036857327094
+     -0.06004475814121585
+        0.305059313826255
+ 4.06e+10    
+       0.3051896700069374
+     -0.06040235687923894
+       0.3118331080460111
+    -0.007040656674429015
+     -0.02737930519903502
+       0.3109475511210056
+    -0.003268818078202675
+    -0.007039672767546391
+     -0.06021605675791622
+       0.3056687695013438
+ 4.07e+10    
+       0.3057986438003348
+     -0.06057470800908097
+       0.3124894889877428
+    -0.007071068944620779
+     -0.02746946858639422
+       0.3116021244324733
+    -0.003262202550226768
+    -0.007070204100401599
+      -0.0603875441197301
+       0.3062773800141784
+ 4.08e+10    
+       0.3064067769019394
+     -0.06074724674360749
+       0.3131452290706582
+    -0.007101372739093987
+     -0.02755981690736633
+       0.3122560571101816
+    -0.003255334080177872
+    -0.007100628329564842
+     -0.06055921556861289
+       0.3068851429310379
+ 4.09e+10    
+       0.3070140667663192
+      -0.0609199684357995
+       0.3138003259478859
+    -0.007131565545070931
+     -0.02765035024011413
+       0.3129093466739142
+    -0.003248209351901014
+    -0.007130942928173413
+     -0.06073106639588214
+       0.3074920557616435
+ 4.1e+10     
+        0.307620510794588
+     -0.06109286838999917
+       0.3144547772409448
+    -0.007161644850053397
+     -0.02774106866325381
+       0.3135619906126269
+    -0.003240825024675442
+    -0.007161145369190889
+     -0.06090309184378787
+       0.3080981159602808
+ 4.11e+10    
+       0.3082261063355297
+     -0.06126594186346145
+       0.3151085805404082
+    -0.007191608142178597
+     -0.02783197225592515
+       0.3142139863851582
+    -0.003233177734100055
+    -0.007191233125767372
+      -0.0610752871070903
+       0.3087033209269333
+ 4.12e+10    
+       0.3088308506867302
+      -0.0614391840679137
+       0.3157617334065776
+    -0.007221452910573561
+     -0.02792306109785909
+       0.3148653314209481
+    -0.003225264092997672
+      -0.0072212036715982
+     -0.06124764733464716
+       0.3093076680084318
+ 4.13e+10    
+       0.3094347410957221
+     -0.06161259017112408
+        0.316414233370164
+    -0.007251176645707957
+     -0.02801433526944416
+       0.3155160231207613
+    -0.003217080692337634
+    -0.007251054481281254
+     -0.06142016763100661
+       0.3099111544996062
+ 4.14e+10    
+       0.3100377747611358
+     -0.06178615529847459
+       0.3170660779329723
+    -0.007280776839745168
+     -0.02810579485179042
+       0.3161660588574203
+    -0.003208624102176968
+    -0.007280783030672727
+     -0.06159284305800942
+        0.310513777644455
+ 4.15e+10    
+       0.3106399488338598
+     -0.06195987453454353
+       0.3177172645685994
+    -0.007310250986891618
+     -0.02819743992679195
+       0.3168154359765427
+    -0.003199890872619543
+    -0.007310386797241388
+     -0.06176566863639602
+       0.3111155346373186
+ 4.16e+10    
+       0.3112412604182112
+       -0.062133742924692
+       0.3183677907231319
+    -0.007339596583744183
+     -0.02828927057718721
+        0.317464151797284
+    -0.003190877534793463
+    -0.007339863260420992
+     -0.06193863934742053
+       0.3117164226240626
+ 4.17e+10    
+       0.3118417065731103
+     -0.06230775547665737
+       0.3190176538158568
+    -0.007368811129635839
+     -0.02838128688661752
+       0.3181122036130866
+    -0.003181580601846201
+    -0.007369209901961181
+     -0.06211175013447102
+       0.3123164387032708
+ 4.18e+10    
+       0.3124412843132637
+     -0.06248190716215172
+       0.3196668512399722
+    -0.007397892126978993
+     -0.02847348893968396
+       0.3187595886924356
+    -0.003171996569957451
+    -0.007398424206276184
+     -0.06228499590469396
+       0.3129155799274426
+ 4.19e+10    
+       0.3130399906103566
+     -0.06265619291846598
+       0.3203153803633113
+    -0.007426837081607032
+     -0.02856587682200216
+       0.3194063042796161
+    -0.003162121919369626
+    -0.007427503660792079
+     -0.06245837153062533
+       0.3135138433042018
+ 4.2e+10     
+       0.3136378223942464
+     -0.06283060765007718
+       0.3209632385290613
+    -0.007455643503113523
+     -0.02865845062025496
+        0.320052347595479
+    -0.003151953115435489
+     -0.00745644575629149
+     -0.06263187185182412
+       0.3141112257975056
+ 4.21e+10    
+       0.3142347765541632
+     -0.06300514623026146
+       0.3216104230565016
+    -0.007484308905189114
+     -0.02875121042224457
+       0.3206977158382104
+    -0.003141486609683056
+      -0.0074852479872566
+     -0.06280549167651266
+       0.3147077243288667
+ 4.22e+10    
+       0.3148308499399183
+     -0.06317980350270953
+        0.322256931241732
+    -0.007512830805956235
+     -0.02884415631694084
+       0.3213424061841027
+    -0.003130718840897449
+    -0.007513907852209898
+      -0.0629792257832175
+       0.3153033357785744
+ 4.23e+10    
+       0.3154260393631148
+     -0.06335457428314693
+       0.3229027603584184
+     -0.00754120672830142
+     -0.02893728839452962
+       0.3219864157883334
+    -0.003119646236219463
+    -0.007542422854052648
+     -0.06315306892241654
+       0.3158980569869249
+ 4.24e+10    
+       0.3160203415983611
+     -0.06352945336095597
+       0.3235479076585352
+    -0.007569434200204981
+     -0.02903060674645835
+        0.322629741785746
+    -0.003108265212260612
+    -0.007570790500401093
+     -0.06332701581818723
+       0.3164918847554548
+ 4.25e+10    
+       0.3166137533844911
+     -0.06370443550080043
+       0.3241923703731159
+    -0.007597510755068423
+     -0.02912411146548017
+       0.3232723812916347
+    -0.003096572176234563
+     -0.00759900830392022
+     -0.06350106116985815
+       0.3170848158481773
+ 4.26e+10    
+       0.3172062714257871
+      -0.0638795154442546
+       0.3248361457130066
+    -0.007625433932038909
+     -0.02921780264569635
+        0.323914331402532
+    -0.003084563527104629
+     -0.00762707378265522
+     -0.06367519965366283
+       0.3176768469928256
+ 4.27e+10    
+       0.3177978923932025
+     -0.06405468791143028
+       0.3254792308696212
+    -0.007653201276331439
+     -0.02931168038259655
+       0.3245555891969997
+    -0.003072235656747146
+    -0.007654984460360333
+      -0.0638494259243943
+       0.3182679748820945
+ 4.28e+10    
+       0.3183886129255922
+     -0.06422994760260928
+       0.3261216230157054
+    -0.007680810339547921
+     -0.02940574477309826
+       0.3251961517364237
+    -0.003059584951130455
+    -0.007682737866825018
+     -0.06402373461706271
+       0.3188581961748903
+ 4.29e+10    
+       0.3189784296309402
+     -0.06440528919987452
+       0.3267633193060989
+     -0.00770825867999377
+     -0.02949999591558372
+       0.3258360160658097
+    -0.003046607791509287
+    -0.007710331538197735
+     -0.06419812034855221
+       0.3194475074975764
+ 4.3e+10     
+       0.3195673390875935
+     -0.06458070736874301
+       0.3274043168785036
+    -0.007735543862991467
+     -0.02959443390993536
+       0.3264751792145831
+    -0.003033300555634237
+    -0.007737763017306807
+     -0.06437257771928054
+       0.3200359054452293
+ 4.31e+10    
+       0.3201553378454919
+     -0.06475619675979875
+       0.3280446128542538
+    -0.007762663461191188
+     -0.02968905885757013
+       0.3271136381973898
+    -0.003019659618976296
+    -0.007765029853978575
+     -0.06454710131485662
+       0.3206233865828886
+ 4.32e+10    
+       0.3207424224274044
+     -0.06493175201032625
+       0.3286842043390881
+    -0.007789615054878529
+     -0.02978387086147152
+       0.3277513900148995
+    -0.003005681355965765
+    -0.007792129605352725
+      -0.0647216857077402
+       0.3212099474468122
+ 4.33e+10    
+       0.3213285893301646
+     -0.06510736774594368
+       0.3293230884239282
+    -0.007816396232279222
+     -0.02987887002622039
+       0.3283884316546107
+    -0.002991362141245745
+    -0.007819059836194724
+     -0.06489632545889942
+       0.3217955845457304
+ 4.34e+10    
+       0.3219138350259034
+     -0.06528303858223465
+       0.3299612621856526
+    -0.007843004589860742
+     -0.02997405645802419
+       0.3290247600916592
+    -0.002976698350939601
+    -0.007845818119205348
+      -0.0650710151194696
+       0.3223802943621038
+ 4.35e+10    
+       0.3224981559632858
+     -0.06545875912638048
+       0.3305987226878792
+    -0.007869437732630597
+     -0.03006943026474447
+       0.3296603722896223
+     -0.00296168636393231
+    -0.007872402035327099
+     -0.06524574923240828
+       0.3229640733533765
+ 4.36e+10    
+       0.3230815485687444
+     -0.06563452397878958
+       0.3312354669817454
+    -0.007895693274431745
+     -0.03016499155592295
+       0.3302952652013321
+      -0.0029463225631653
+    -0.007898809174047772
+      -0.0654205223341518
+       0.3235469179532341
+ 4.37e+10    
+        0.323664009247716
+     -0.06581032773472723
+       0.3318714921066935
+    -0.007921768838234505
+     -0.03026074044280658
+       0.3309294357696835
+    -0.002930603336944597
+    -0.007925037133700609
+     -0.06559532895626782
+       0.3241288245728563
+ 4.38e+10    
+       0.3242455343858729
+     -0.06598616498594162
+       0.3325067950912537
+    -0.007947662056425308
+        -0.03035667703837
+       0.3315628809284454
+    -0.002914525080261812
+    -0.007951083521761694
+     -0.06577016362710693
+       0.3247097896021739
+ 4.39e+10    
+       0.3248261203503555
+     -0.06616203032228837
+       0.3331413729538305
+     -0.00797337057109208
+     -0.03045280145733792
+       0.3321955976030737
+    -0.002898084196127866
+    -0.007976945955143583
+     -0.06594502087345207
+       0.3252898094111196
+ 4.4e+10     
+        0.325405763491003
+     -0.06633791833335298
+       0.3337752227034899
+    -0.007998892034306152
+     -0.03054911381620504
+       0.3328275827115207
+    -0.002881277096919086
+    -0.008002622060486481
+     -0.06611989522216373
+       0.3258688803508815
+ 4.41e+10    
+       0.3259844601415844
+     -0.06651382361007027
+       0.3344083413407477
+    -0.008024224108401007
+     -0.03064561423325519
+       0.3334588331650506
+    -0.002864100205735192
+    -0.008028109474445207
+     -0.06629478120182439
+       0.3264469987551517
+ 4.42e+10    
+       0.3265622066210221
+     -0.06668974074633986
+        0.335040725858358
+    -0.008049364466247199
+     -0.03074230282857898
+       0.3340893458690502
+    -0.002846549957769173
+    -0.008053405843973498
+     -0.06646967334437813
+       0.3270241609413763
+ 4.43e+10    
+       0.3271389992346187
+     -0.06686566434063929
+       0.3356723732421015
+    -0.008074310791524002
+     -0.03083917972408975
+       0.3347191177238401
+    -0.002828622801688398
+    -0.008078508826604639
+     -0.06664456618676606
+       0.3276003632119978
+ 4.44e+10    
+       0.3277148342752776
+      -0.0670415889976327
+       0.3363032804715764
+    -0.008099060778987432
+     -0.03093624504353909
+       0.3353481456254884
+     -0.00281031520102685
+    -0.008103416090728743
+     -0.06681945427255992
+       0.3281756018557022
+ 4.45e+10    
+       0.3282897080247247
+     -0.06721750932977645
+       0.3369334445209871
+    -0.008123612134734785
+     -0.03103349891253039
+       0.3359764264666216
+    -0.002791623635588085
+    -0.008128125315866522
+     -0.06699433215358971
+       0.3287498731486563
+ 4.46e+10    
+       0.3288636167547218
+     -0.06739341995891911
+       0.3375628623599324
+    -0.008147962576465356
+     -0.03113094145853106
+       0.3366039571372343
+    -0.002772544602858562
+    -0.008152634192939472
+     -0.06716919439156732
+       0.3293231733557467
+ 4.47e+10    
+       0.3294365567282811
+     -0.06756931551789788
+       0.3381915309541988
+    -0.008172109833737611
+     -0.03122857281088445
+       0.3372307345255006
+     -0.00275307461943096
+    -0.008176940424536856
+     -0.06734403555970515
+       0.3298954987318128
+ 4.48e+10    
+       0.3300085242008738
+     -0.06774519065212931
+       0.3388194472665431
+    -0.008196051648222891
+      -0.0313263931008195
+       0.3378567555185825
+     -0.00273321022243721
+    -0.008201041725178552
+     -0.06751885024433063
+        0.330466845522877
+ 4.49e+10    
+       0.3305795154216368
+     -0.06792104002119705
+       0.3394466082574879
+     -0.00821978577395484
+     -0.03142440246146019
+       0.3384820170034378
+    -0.002712947970990866
+    -0.008224935821574984
+     -0.06769363304649384
+       0.3310372099673725
+ 4.5e+10     
+       0.3311495266345715
+     -0.06809685830043016
+       0.3400730108861033
+    -0.008243309977575837
+     -0.03152260102783339
+       0.3391065158676266
+    -0.002692284447638362
+    -0.008248620452882684
+     -0.06786837858357096
+       0.3316065882973637
+ 4.51e+10    
+       0.3317185540797463
+     -0.06827264018248046
+       0.3406986521107966
+    -0.008266622038578843
+     -0.03162098893687559
+       0.3397302490001153
+    -0.002671216259818932
+    -0.008272093370956855
+     -0.06804308149086025
+       0.3321749767397655
+ 4.52e+10    
+       0.3322865939944828
+     -0.06844838037889006
+       0.3413235288900973
+    -0.008289719749546259
+     -0.03171956632743907
+       0.3403532132920831
+    -0.002649740041332606
+    -0.008295352340599783
+     -0.06821773642317414
+       0.3327423715175579
+ 4.53e+10    
+         0.33285364261455
+     -0.06862407362165562
+       0.3419476381834415
+    -0.008312600916384289
+     -0.03181833334029673
+       0.3409754056377212
+    -0.002627852453816205
+     -0.00831839513980568
+     -0.06839233805642214
+       0.3333087688509924
+ 4.54e+10    
+       0.3334196961753435
+     -0.06879971466478368
+       0.3425709769519548
+    -0.008335263358553887
+     -0.03191729011814576
+       0.3415968229350319
+    -0.002605550188226633
+    -0.008341219560001889
+     -0.06856688108918935
+       0.3338741649587977
+ 4.55e+10    
+        0.333984750913067
+     -0.06897529828584194
+       0.3431935421592344
+    -0.008357704909297561
+     -0.03201643680561114
+       0.3422174620866293
+    -0.002582829966331311
+     -0.00836382340628614
+     -0.06874136024430708
+       0.3344385560593793
+ 4.56e+10    
+       0.3345488030659024
+      -0.0691508192875006
+       0.3438153307721274
+    -0.008379923415862679
+     -0.03211577354924722
+        0.342837320000533
+    -0.002559688542205172
+    -0.008386204497660107
+     -0.06891577027041537
+       0.3350019383720088
+ 4.57e+10    
+       0.3351118488751815
+     -0.06932627249907038
+       0.3444363397615129
+    -0.008401916739720378
+     -0.03221530049753962
+       0.3434563935909619
+    -0.002536122703734017
+    -0.008408360667259265
+     -0.06909010594352076
+       0.3355643081180178
+ 4.58e+10    
+       0.3356738845865433
+     -0.06950165277802818
+       0.3450565661030718
+    -0.008423682756780963
+     -0.03231501780090499
+        0.344074679779124
+     -0.00251212927412358
+    -0.008430289762578681
+     -0.06926436206854319
+       0.3361256615219744
+ 4.59e+10    
+       0.3362349064510943
+       -0.069676955011541
+        0.345676006778068
+    -0.008445219357605173
+     -0.03241492561169129
+       0.3446921754940064
+    -0.002487705113414195
+    -0.008451989645695164
+     -0.06943853348085748
+       0.3366859948128638
+ 4.6e+10     
+       0.3367949107265568
+     -0.06985217411797628
+       0.3462946587741139
+    -0.008466524447611628
+     -0.03251502408417623
+       0.3453088776731604
+    -0.002462847120000345
+    -0.008473458193485521
+     -0.06961261504782527
+       0.3372453042252551
+ 4.61e+10    
+       0.3373538936784127
+     -0.07002730504840833
+       0.3469125190859446
+    -0.008487595947280137
+     -0.03261531337456608
+       0.3459247832634819
+    -0.002437552232154843
+    -0.008494693297840836
+       -0.069786601670319
+       0.3378035860004668
+ 4.62e+10    
+       0.3379118515810431
+     -0.07020234278811453
+       0.3475295847161823
+    -0.008508431792351355
+     -0.03271579364099259
+       0.3465398892219942
+    -0.002411817429557233
+    -0.008515692865877172
+     -0.06996048828423773
+       0.3383608363877245
+ 4.63e+10    
+       0.3384687807188588
+     -0.07037728235806326
+       0.3481458526761014
+    -0.008529029934022273
+     -0.03281646504351024
+       0.3471541925166231
+    -0.002385639734825863
+    -0.008536454820141846
+     -0.07013426986201365
+       0.3389170516453099
+ 4.64e+10    
+       0.3390246773874243
+      -0.0705521188163938
+       0.3487613199863899
+    -0.008549388339137601
+     -0.03291732774409235
+       0.3477676901269689
+    -0.002359016215053345
+    -0.008556977098816532
+     -0.07030794141410937
+       0.3394722280417059
+ 4.65e+10    
+       0.3395795378945764
+     -0.07072684725988609
+       0.3493759836779083
+    -0.008569504990377603
+     -0.03301838190662703
+       0.3483803790450791
+    -0.002331943983344808
+    -0.008577257655915708
+     -0.07048149799050708
+       0.3400263618567336
+ 4.66e+10    
+       0.3401333585615362
+     -0.07090146282542296
+       0.3499898407924454
+    -0.008589377886441466
+     -0.03311962769691221
+        0.348992256276212
+    -0.002304420200358674
+    -0.008597294461481877
+     -0.07065493468218652
+       0.3405794493826817
+ 4.67e+10    
+       0.3406861357240109
+     -0.07107596069144126
+       0.3506028883834706
+    -0.008609005042227186
+     -0.03322106528265031
+       0.3496033188396032
+    -0.002276442075849297
+    -0.008617085501776346
+     -0.07082824662259546
+        0.341131486925428
+ 4.68e+10    
+        0.341237865733292
+     -0.07125033607937512
+       0.3512151235168836
+    -0.008628384489006944
+     -0.03332269483344257
+       0.3502135637692195
+      -0.0022480068702113
+    -0.008636628779466533
+     -0.07100142898910852
+        0.341682470805558
+ 4.69e+10    
+       0.3417885449573445
+     -0.07142458425508849
+       0.3518265432717594
+    -0.008647514274599056
+     -0.03342451652078282
+       0.3508229881145195
+    -0.002219111896024765
+     -0.00865592231380889
+     -0.07117447700447668
+       0.3422323973594673
+ 4.7e+10     
+       0.3423381697818872
+     -0.07159870053029771
+       0.3524371447410922
+    -0.008666392463535606
+     -0.03352653051805064
+       0.3514315889412017
+    -0.002189754519601343
+    -0.008674964140828511
+     -0.07134738593826698
+       0.3427812629404659
+ 4.71e+10    
+       0.3428867366114695
+     -0.07177268026398465
+       0.3530469250325332
+    -0.008685017137226159
+     -0.03362873700050496
+       0.3520393633319538
+    -0.002159932162530236
+    -0.008693752313494247
+     -0.07152015110829094
+       0.3433290639198679
+ 4.72e+10    
+       0.3434342418705346
+     -0.07194651886379952
+       0.3536558812691256
+    -0.008703386394117666
+     -0.03373113614527627
+       0.3526463083871942
+    -0.002129642303224037
+    -0.008712284901890292
+     -0.07169276788202332
+       0.3438757966880753
+ 4.73e+10    
+         0.34398068200448
+     -0.07212021178745241
+       0.3542640105900374
+    -0.008721498349850252
+     -0.03383372813135936
+       0.3532524212258128
+    -0.002098882478463792
+    -0.008730559993383954
+     -0.07186523167800914
+       0.3444214576556558
+ 4.74e+10    
+       0.3445260534807069
+     -0.07229375454409522
+        0.354871310151287
+    -0.008739351137409283
+     -0.03393651313960529
+       0.3538576989859047
+    -0.002067650284942828
+    -0.008748575692788979
+     -0.07203753796726103
+       0.3449660432544081
+ 4.75e+10    
+       0.3450703527896631
+     -0.07246714269569211
+       0.3554777771264682
+    -0.008756942907273291
+     -0.03403949135271378
+       0.3544621388255003
+    -0.002035943380808741
+    -0.008766330122525839
+     -0.07220968227464371
+       0.3455095499384221
+ 4.76e+10    
+       0.3456135764458755
+      -0.0726403718583796
+       0.3560834087074685
+    -0.008774271827558057
+     -0.03414266295522445
+       0.3550657379232908
+    -0.002003759487203364
+    -0.008783821422777425
+     -0.07238166018024897
+         0.34605197418513
+ 4.77e+10    
+       0.3461557209889773
+     -0.07281343770381499
+       0.3566882021051846
+    -0.008791336084157003
+     -0.03424602813350892
+       0.3556684934793506
+    -0.001971096389800028
+    -0.008801047751641209
+     -0.07255346732075847
+       0.3465933124963474
+ 4.78e+10    
+       0.3466967829847243
+     -0.07298633596051393
+       0.3572921545502324
+    -0.008808133880877372
+     -0.03434958707576219
+       0.3562704027158521
+     -0.00193795194033755
+    -0.008818007285277759
+     -0.07272509939079412
+       0.3471335613993078
+ 4.79e+10    
+       0.3472367590260018
+     -0.07315906241517618
+       0.3578952632936543
+    -0.008824663439572895
+     -0.03445333997199411
+        0.356871462877779
+    -0.001904324058150724
+    -0.008834698218054941
+     -0.07289655214425893
+       0.3476727174476863
+ 4.8e+10     
+       0.3477756457338264
+     -0.07333161291400063
+       0.3584975256076215
+    -0.008840923000272229
+     -0.03455728701402094
+       0.3574716712336304
+    -0.001870210731696636
+    -0.008851118762688834
+      -0.0730678213956629
+       0.3482107772226149
+ 4.81e+10    
+       0.3483134397583353
+      -0.0735039833639874
+       0.3590989387861283
+    -0.008856910821304067
+     -0.03466142839545651
+       0.3580710250761252
+    -0.001835610020076403
+    -0.008867267150380477
+     -0.07323890302143982
+       0.3487477373336906
+ 4.82e+10    
+       0.3488501377797687
+     -0.07367616973422897
+       0.3596995001456882
+    -0.008872625179417977
+     -0.03476576431170396
+       0.3586695217228965
+    -0.001800520054551724
+    -0.008883141630949078
+     -0.07340979296124972
+       0.3492835944199699
+ 4.83e+10    
+        0.349385736509442
+     -0.07384816805718929
+       0.3602992070260199
+    -0.008888064369901808
+     -0.03487029495994707
+       0.3592671585171838
+     -0.00176493904005594
+    -0.008898740472961436
+     -0.07358048721927021
+       0.3498183451509597
+ 4.84e+10    
+       0.3499202326907099
+     -0.07401997442997028
+       0.3608980567907302
+    -0.008903226706695194
+     -0.03497502053914193
+       0.3598639328285201
+    -0.001728865256698977
+    -0.008914061963857524
+     -0.07375098186547507
+       0.3503519862275942
+ 4.85e+10    
+        0.350453623099921
+     -0.07419158501556658
+       0.3614960468279916
+    -0.008918110522499412
+      -0.0350799412500087
+       0.3604598420534114
+    -0.001692297061265682
+    -0.008929104410072584
+     -0.07392127303689976
+       0.3508845143832048
+ 4.86e+10    
+       0.3509859045473619
+     -0.07436299604410763
+       0.3620931745512168
+    -0.008932714168883431
+     -0.03518505729502337
+       0.3610548836160121
+    -0.001655232888707051
+    -0.008943866137155306
+      -0.0740913569388949
+       0.3514159263844786
+ 4.87e+10    
+       0.3515170738781938
+     -0.07453420381408714
+        0.362689437399723
+    -0.008947036016386514
+     -0.03529036887841005
+       0.3616490549687968
+    -0.001617671253624013
+    -0.008958345489882636
+     -0.07426122984636636
+       0.3519462190324107
+ 4.88e+10    
+       0.3520471279733778
+     -0.07470520469358052
+       0.3632848328393997
+    -0.008961074454616949
+     -0.03539587620613316
+       0.3622423535932229
+    -0.001579610751743002
+    -0.008972540832370693
+     -0.07443088810500272
+        0.352475389163242
+ 4.89e+10    
+       0.3525760637505921
+      -0.0748759951214488
+        0.363879358363361
+    -0.008974827892347371
+      -0.0355015794858899
+       0.3628347770003892
+    -0.001541050061382998
+    -0.008986450548182322
+     -0.07460032813248932
+       0.3530034336493905
+ 4.9e+10     
+       0.3531038781651387
+     -0.07504657160853045
+       0.3644730114926005
+    -0.008988294757606357
+     -0.03560747892710332
+       0.3634263227316918
+     -0.00150198794491352
+    -0.009000073040431038
+      -0.0747695464197099
+       0.3535303494003727
+ 4.91e+10    
+       0.3536305682108398
+      -0.0752169307388191
+       0.3650657897766362
+    -0.009001473497766765
+     -0.03571357474091531
+       0.3640169883594677
+    -0.001462423250203034
+      -0.0090134067318812
+     -0.07493853953193311
+       0.3540561333637127
+ 4.92e+10    
+       0.3541561309209269
+     -0.07538706917063062
+       0.3656576907941548
+     -0.00901436257963009
+      -0.0358198671401804
+         0.36460677148764
+    -0.001422354912057232
+    -0.009026450065045205
+     -0.07510730410998809
+        0.354580782525843
+ 4.93e+10    
+       0.3546805633689158
+     -0.07555698363775279
+       0.3662487121536406
+    -0.009026960489507978
+     -0.03592635633945918
+       0.3651956697523511
+    -0.001381781953646846
+    -0.009039201502276587
+     -0.07527583687142461
+       0.3551042939129962
+ 4.94e+10    
+       0.3552038626694767
+     -0.07572667095058742
+       0.3668388514940149
+    -0.009039265733299788
+      -0.0360330425550132
+       0.3657836808225933
+    -0.001340703487924198
+    -0.009051659525860362
+     -0.07544413461165995
+       0.3556266645920824
+ 4.95e+10    
+        0.355726025979289
+     -0.07589612799727308
+       0.3674281064852504
+    -0.009051276836567054
+     -0.03613992600479913
+       0.3663708024008324
+    -0.001299118719028448
+    -0.009063822638099361
+     -0.07561219420511282
+       0.3561478916715614
+ 4.96e+10    
+        0.356247050497891
+     -0.07606535174479953
+        0.368016474828997
+    -0.009062992344604483
+     -0.03624700690846457
+       0.3669570322236264
+    -0.001257026943678482
+    -0.009075689361397639
+     -0.07578001260632342
+       0.3566679723023023
+ 4.97e+10    
+       0.3567669334685145
+      -0.0762343392401045
+       0.3686039542591896
+    -0.009074410822507862
+     -0.03635428548734339
+       0.3675423680622357
+    -0.001214427552553382
+    -0.009087258238340362
+     -0.07594758685105753
+       0.3571869036784295
+ 4.98e+10    
+       0.3572856721789145
+     -0.07640308761116063
+       0.3691905425426592
+    -0.009085530855238253
+     -0.03646176196445208
+       0.3681268077232281
+    -0.001171320031659775
+    -0.009098527831770641
+     -0.07611491405739962
+       0.3577046830381652
+ 4.99e+10    
+       0.3578032639621838
+     -0.07657159406804542
+       0.3697762374797307
+    -0.009096351047683585
+     -0.03656943656448688
+       0.3687103490490816
+    -0.001127703963685606
+    -0.009109496724862755
+     -0.07628199142683109
+       0.3582213076646558
+ 5e+10       
+       0.3583197061975608
+      -0.0767398559039989
+       0.3703610369048178
+    -0.009106870024716543
+     -0.03667730951382045
+       0.3692929899187714
+    -0.001083579029339873
+      -0.0091201635211926
+     -0.07644881624529136
+       0.3587367748867877
+ 5.01e+10    
+       0.3588349963112236
+     -0.07690787049646809
+       0.3709449386870134
+    -0.009117086431249519
+     -0.03678538104050073
+       0.3698747282483613
+    -0.001038945008677753
+    -0.009130526844804605
+     -0.07661538588422945
+       0.3592510820799962
+ 5.02e+10    
+       0.3593491317770778
+     -0.07707563530813652
+       0.3715279407306727
+    -0.009126998932286653
+      -0.0368936513742493
+       0.3704555619915831
+   -0.0009938017824106357
+    -0.009140585340276024
+     -0.07678169780163881
+       0.3597642266670635
+ 5.03e+10    
+       0.3598621101175292
+     -0.07724314788793932
+       0.3721100409759873
+    -0.009136606212972541
+     -0.03700212074646027
+       0.3710354891404074
+   -0.0009481493332006872
+    -0.009150337672777547
+     -0.07694774954307659
+       0.3602762061188988
+ 5.04e+10    
+       0.3603739289042495
+     -0.07741040587206562
+       0.3726912373995573
+    -0.009145906978638096
+     -0.03711078939020097
+       0.3716145077256139
+   -0.0009019877469393877
+    -0.009159782528131436
+     -0.07711353874267085
+       0.3607870179553169
+ 5.05e+10    
+       0.3608845857589301
+     -0.07757740698494621
+       0.3732715280149552
+    -0.009154899954843568
+     -0.03721965754021225
+       0.3721926158173514
+   -0.0008553172140093811
+    -0.009168918612866431
+      -0.0772790631241127
+       0.3612966597458012
+ 5.06e+10    
+       0.3613940783540262
+     -0.07774414904022689
+       0.3738509108732855
+    -0.009163583887418439
+      -0.0373287254329103
+       0.3727698115256912
+   -0.0008081380305294788
+    -0.009177744654269697
+     -0.07744432050163269
+       0.3618051291102567
+ 5.07e+10    
+       0.3619024044134863
+     -0.07791062994172716
+       0.3744293840637327
+    -0.009171957542498707
+     -0.03743799330638863
+       0.3733460930011755
+    -0.000760450599582099
+    -0.009186259400436074
+     -0.07760930878096378
+       0.3623124237197503
+ 5.08e+10    
+       0.3624095617134774
+      -0.0780768476843859
+       0.3750069457141086
+    -0.009180019706561226
+     -0.03754746140042122
+       0.3739214584353576
+   -0.0007122554324226586
+    -0.009194461620314336
+     -0.07777402596028969
+        0.362818541297245
+ 5.09e+10    
+       0.3629155480830949
+     -0.07824280035519163
+       0.3755835939913917
+     -0.00918776918645535
+     -0.03765712995646647
+       0.3744959060613366
+   -0.0006635531496707143
+     -0.00920235010375073
+     -0.07793847013117766
+       0.3633234796183163
+ 5.1e+10     
+       0.3634203614050621
+     -0.07840848613409876
+       0.3761593271022589
+    -0.009195204809431938
+      -0.0377669992176719
+       0.3750694341542851
+   -0.0006143444824818762
+    -0.009209923661529795
+     -0.07810263947949744
+       0.3638272365118643
+ 5.11e+10    
+       0.3639239996164208
+     -0.07857390329492941
+       0.3767341432936094
+    -0.009202325423169604
+      -0.0378770694288796
+       0.3756420410319692
+   -0.0005646302737005989
+    -0.009217181125412468
+     -0.07826653228632469
+       0.3643298098608095
+ 5.12e+10    
+       0.3644264607092105
+      -0.0787390502062608
+       0.3773080408530872
+    -0.009209129895798612
+     -0.03798734083663306
+       0.3762137250552633
+   -0.0005144114789929302
+    -0.009224121348171535
+     -0.07843014692883055
+       0.3648311976027809
+ 5.13e+10    
+        0.364927742731134
+     -0.07890392533229822
+       0.3778810181095917
+     -0.00921561711592183
+     -0.03809781368918413
+       0.3767844846286562
+   -0.0004636891679590015
+     -0.00923074320362471
+      -0.0785934818811551
+       0.3653313977307913
+ 5.14e+10    
+       0.3654278437862163
+     -0.07906852723373299
+       0.3784530734337841
+    -0.009221785992633869
+     -0.03820848823650169
+       0.3773543182007536
+   -0.0004124645252246994
+    -0.009237045586664753
+     -0.07875653571526757
+       0.3658304082939017
+ 5.15e+10    
+       0.3659267620354503
+     -0.07923285456858693
+       0.3790242052385878
+    -0.009227635455536953
+     -0.03831936473028075
+       0.3779232242647674
+   -0.0003607388515120958
+    -0.009243027413287534
+     -0.07891930710180932
+       0.3663282273978752
+ 5.16e+10    
+        0.366424495697432
+     -0.07939690609304126
+       0.3795944119796799
+     -0.00923316445475522
+      -0.0384304434239528
+       0.3784912013590075
+   -0.0003085135646881914
+    -0.009248687620617519
+     -0.07908179481092473
+       0.3668248532058192
+ 5.17e+10    
+       0.3669210430489835
+     -0.07956068066225075
+       0.3801636921559774
+    -0.009238371960946255
+     -0.03854172457269692
+       0.3790582480673554
+   -0.0002557902007915269
+    -0.009254025166930871
+     -0.07924399771307424
+       0.3673202839388158
+ 5.18e+10    
+       0.3674164024257671
+     -0.07972417723114454
+       0.3807320443101179
+    -0.009243256965310412
+      -0.0386532084334525
+       0.3796243630197444
+   -0.0002025704150360852
+    -0.009259039031676117
+      -0.0794059147798358
+       0.3678145178765433
+ 5.19e+10    
+       0.3679105722228882
+     -0.07988739485521104
+       0.3812994670289312
+    -0.009247818479598172
+     -0.03876489526493204
+       0.3801895448926164
+   -0.0001488559827923835
+    -0.009263728215492839
+     -0.07956754508468671
+       0.3683075533578825
+ 5.2e+10     
+        0.368403550895485
+     -0.08005033269126877
+       0.3818659589439042
+     -0.00925205553611508
+      -0.0388767853276358
+       0.3807537924093877
+   -9.464880054493776e-05
+     -0.00926809174022789
+     -0.07972888780377571
+       0.3687993887815167
+ 5.21e+10    
+       0.3688953369593101
+     -0.08021298999822223
+       0.3824315187316426
+    -0.009255967187724789
+      -0.0389888788838671
+       0.3813171043408964
+    -3.99508868258291e-05
+    -0.009272128648949728
+     -0.07988994221667589
+       0.3692900226065159
+ 5.22e+10    
+       0.3693859289912984
+     -0.08037536613780352
+       0.3829961451143195
+    -0.009259552507849968
+     -0.03910117619774909
+       0.3818794795058488
+    1.523561687584375e-05
+    -0.009275838005960107
+     -0.08005070770712427
+       0.3697794533529118
+ 5.23e+10    
+       0.3698753256301267
+     -0.08053746057529883
+       0.3835598368601252
+    -0.009262810590471396
+     -0.03921367753524238
+       0.3824409167712568
+    7.090844522952876e-05
+      -0.0092792188968046
+     -0.08021118376374708
+       0.3702676796022639
+ 5.24e+10    
+       0.3703635255767604
+     -0.08069927288026055
+          0.3841225927837
+    -0.009265740550124925
+     -0.03932638316416352
+       0.3830014150528668
+    0.0001270652082035744
+    -0.009282270428280172
+     -0.08037136998076806
+       0.3707546999982087
+ 5.25e+10    
+       0.3708505275949884
+     -0.08086080272720444
+       0.3846844117465714
+    -0.009268341521896697
+     -0.03943929335420538
+       0.3835609733155849
+    0.0001837033902314586
+    -0.009284991728441563
+     -0.08053126605870352
+       0.3712405132470019
+ 5.26e+10    
+       0.3713363305119504
+     -0.08102204989629247
+        0.385245292657577
+    -0.009270612661416634
+     -0.03955240837695805
+       0.3841195905738924
+    0.0002408203494037374
+    -0.009287381946605465
+     -0.08069087180504186
+       0.3717251181180508
+ 5.27e+10    
+       0.3718209332186497
+     -0.08118301427400018
+       0.3858052344732771
+    -0.009272553144850258
+     -0.03966572850593078
+       0.3846772658922533
+    0.0002984133166864049
+    -0.009289440253352724
+     -0.08085018713490669
+       0.3722085134444288
+ 5.28e+10    
+       0.3723043346704565
+     -0.08134369585377084
+        0.386364236198375
+     -0.00927416216888842
+      -0.0397792540165763
+       0.3852339983855194
+    0.0003564793951658996
+    -0.009291165840529237
+     -0.08100921207170764
+       0.3726906981233863
+ 5.29e+10    
+       0.3727865338876014
+     -0.08150409473665331
+       0.3869222968861134
+    -0.009275438950735945
+     -0.03989298518631455
+       0.3857897872193214
+    0.0004150155593212819
+    -0.009292557921244775
+     -0.08116794674777363
+       0.3731716711168454
+ 5.3e+10     
+       0.3732675299556538
+     -0.08166421113192622
+       0.3874794156386738
+    -0.009276382728098382
+     -0.04000692229455935
+         0.38634463161046
+    0.0004740186543238864
+    -0.009293615729870038
+     -0.08132639140497225
+       0.3736514314518837
+ 5.31e+10    
+       0.3737473220259954
+     -0.08182404535770732
+       0.3880355916075675
+    -0.009276992759167275
+     -0.04012106562274513
+       0.3868985308272836
+    0.0005334853953646789
+    -0.009294338522032741
+     -0.08148454639531461
+       0.3741299782212118
+ 5.32e+10    
+       0.3742259093162766
+      -0.0819835978415476
+       0.3885908239940156
+    -0.009277268322604146
+     -0.04023541545435536
+       0.3874514841900621
+     0.000593412367009948
+    -0.009294725574611229
+     -0.08164241218154411
+       0.3746073105836314
+ 5.33e+10    
+       0.3747032911108672
+     -0.08214286912101244
+        0.389145112049329
+    -0.009277208717522932
+     -0.04034997207495253
+       0.3880034910713555
+    0.0006537960225854102
+    -0.009294776185727525
+     -0.08179998933771132
+       0.3750834277644902
+ 5.34e+10    
+       0.3751794667612911
+     -0.08230185984424579
+       0.3896984550752725
+    -0.009276813263471262
+     -0.04046473577220847
+       0.3885545508963687
+    0.0007146326835893401
+    -0.009294489674738279
+     -0.08195727854973305
+       0.3755583290561197
+ 5.35e+10    
+       0.3756544356866561
+     -0.08246057077052223
+       0.3902508524244322
+    -0.009276081300410121
+      -0.0405797068359374
+        0.389104663143306
+    0.0007759185391347184
+    -0.009293865382224709
+     -0.08211428061593744
+       0.3760320138182673
+ 5.36e+10    
+       0.3761281973740669
+      -0.0826190027707822
+       0.3908023035005662
+     -0.00927501218869276
+     -0.04069488555812886
+       0.3896538273437159
+    0.0008376496454210851
+    -0.009292902669980917
+     -0.08227099644759356
+       0.3765044814785103
+ 5.37e+10    
+       0.3766007513790304
+     -0.08277715682815488
+       0.3913528077589534
+    -0.009273605309042055
+     -0.04081027223298272
+        0.390202043082826
+    0.0008998219252361675
+    -0.009291600921001317
+     -0.08242742706942596
+       0.3769757315326668
+ 5.38e+10    
+       0.3770720973258506
+     -0.08293503403846469
+       0.3919023647067353
+    -0.009271860062527114
+     -0.04092586715694524
+       0.3907493099998756
+     0.000962431167487776
+    -0.009289959539466531
+     -0.08258357362011566
+       0.3774457635451884
+ 5.39e+10    
+       0.3775422349080102
+     -0.08309263561072537
+       0.3924509739032512
+    -0.009269775870538224
+     -0.04104167062874722
+       0.3912956277884379
+     0.001025473026765966
+    -0.009287977950728178
+     -0.08273943735278447
+        0.377914577149547
+ 5.4e+10     
+       0.3780111638885437
+     -0.08324996286761668
+       0.3929986349603603
+    -0.009267352174761764
+     -0.04115768294944164
+       0.3918409961967343
+     0.001088943022936219
+    -0.009285655601292714
+     -0.08289501963546704
+       0.3783821720486092
+ 5.41e+10    
+       0.3784788841004003
+     -0.08340701724595055
+       0.3935453475427672
+    -0.009264588437153264
+     -0.04127390442244518
+       0.3923854150279463
+     0.001152836540763498
+    -0.009282991958804018
+     -0.08305032195156545
+        0.378848548014996
+ 5.42e+10    
+       0.3789453954467916
+     -0.08356380029711931
+       0.3940911113683309
+    -0.009261484139910046
+     -0.04139033535357878
+       0.3929288841405125
+     0.001217148829567668
+    -0.009279986512025115
+     -0.08320534590029119
+       0.3793137048914382
+ 5.43e+10    
+       0.3794106979015343
+     -0.08372031368753208
+       0.3946359262083719
+    -0.009258038785443005
+     -0.04150697605111122
+       0.3934714034484278
+       0.0012818750029106
+    -0.009276638770818907
+     -0.08336009319709266
+       0.3797776425911166
+ 5.44e+10    
+       0.3798747915093808
+     -0.08387655919903625
+        0.395179791887972
+     -0.00925425189634748
+     -0.04162382682580319
+       0.3940129729215266
+      0.00134701003831497
+    -0.009272948266127937
+      -0.0835145656740657
+       0.3802403610979905
+ 5.45e+10    
+       0.3803376763863335
+     -0.08403253872932301
+       0.3957227082862634
+    -0.009250123015373576
+     -0.04174088799095282
+       0.3945535925857641
+     0.001412548777015281
+    -0.009268914549953438
+      -0.0836687652803529
+        0.380701860467119
+ 5.46e+10    
+       0.3807993527199586
+     -0.08418825429232245
+       0.3962646753367162
+    -0.009245651705395564
+     -0.04185815986244323
+       0.3950932625234892
+     0.001478485923741177
+    -0.009264537195333371
+     -0.08382269408252595
+       0.3811621408249691
+ 5.47e+10    
+       0.3812598207696802
+     -0.08434370801858009
+       0.3968056930274143
+     -0.00924083754938103
+     -0.04197564275879065
+       0.3956319828737112
+     0.001544816046533331
+    -0.009259815796320157
+     -0.08397635426495513
+       0.3816212023697141
+ 5.48e+10    
+       0.3817190808670697
+     -0.08449890215562347
+       0.3973457614013287
+    -0.009235680150359088
+     -0.04209333700119464
+        0.396169753832356
+     0.001611533576592151
+    -0.009254749967956999
+     -0.08412974813016313
+       0.3820790453715193
+ 5.49e+10    
+       0.3821771334161225
+       -0.084653839068312
+       0.3978848805565776
+    -0.009230179131388265
+     -0.04221124291358898
+       0.3967065756525182
+     0.001678632808159414
+    -0.009249339346254375
+     -0.08428287809916554
+       0.3825356701728204
+ 5.5e+10     
+        0.382633978893524
+     -0.08480852123917365
+       0.3984230506466861
+    -0.009224334135523971
+     -0.04232936082269505
+       0.3972424486447076
+     0.001746107898433164
+    -0.009243583588165103
+     -0.08443574671179743
+       0.3829910771885882
+ 5.51e+10    
+       0.3830896178489053
+     -0.08496295126872765
+       0.3989602718808348
+    -0.009218144825785446
+     -0.04244769105807528
+       0.3977773731770836
+     0.001813952867516007
+    -0.009237482371559691
+     -0.08458835662702426
+       0.3834452669065851
+ 5.52e+10    
+        0.383544050905093
+     -0.08511713187579469
+       0.3994965445241047
+    -0.009211610885122337
+     -0.04256623395218966
+       0.3983113496756872
+     0.001882161598396917
+     -0.00923103539520042
+     -0.08474071062324035
+       0.3838982398876108
+ 5.53e+10    
+       0.3839972787583392
+     -0.08527106589779046
+       0.4000318688977101
+    -0.009204732016380997
+     -0.04268498984045179
+       0.3988443786246622
+     0.001950727836966837
+    -0.009224242378715599
+     -0.08489281159855197
+       0.3843499967657346
+ 5.54e+10    
+       0.3844493021785522
+     -0.08542475629100868
+       0.4005662453792303
+    -0.009197507942270543
+     -0.04280395906128821
+       0.3993764605664739
+     0.002019645192068127
+    -0.009217103062572767
+     -0.08504466257104731
+       0.3848005382485202
+ 5.55e+10    
+        0.384900122009509
+     -0.08557820613088794
+       0.4010996744028301
+    -0.009189938405328632
+     -0.04292314195619781
+       0.3999075961021158
+     0.002088907135578198
+    -0.009209617208052164
+     -0.08519626667905257
+        0.385249865117243
+ 5.56e+10    
+       0.3853497391690621
+     -0.08573141861226638
+       0.4016321564594763
+    -0.009182023167887007
+     -0.04304253886981341
+       0.4004377858913126
+     0.002158507002527049
+    -0.009201784597219417
+     -0.08534762718137327
+       0.3856979782270902
+ 5.57e+10    
+       0.3857981546493355
+     -0.08588439704962259
+       0.4021636920971456
+     -0.00917376201203704
+      -0.0431621501499647
+       0.4009670306527158
+     0.002228437991249472
+    -0.009193605032898155
+     -0.08549874745752259
+       0.3861448785073554
+ 5.58e+10    
+       0.3862453695169096
+     -0.08603714487730298
+       0.4026942819210269
+    -0.009165154739595125
+     -0.04328197614774235
+       0.4014953311640894
+     0.002298693163571464
+    -0.009185078338642252
+     -0.08564963100793588
+       0.3865905669616218
+ 5.59e+10    
+       0.3866913849129963
+     -0.08618966564973497
+       0.4032239265937139
+    -0.009156201172067868
+     -0.04340201721756368
+       0.4020226882624942
+     0.002369265445031196
+    -0.009176204358707987
+     -0.08580028145417179
+       0.3870350446679368
+ 5.6e+10     
+       0.3871362020536063
+     -0.08634196304162856
+       0.4037526268353959
+    -0.009146901150617481
+      -0.0435222737172401
+       0.4025491028444595
+     0.002440147625134731
+    -0.009166982958025946
+     -0.08595070253909881
+       0.3874783127789743
+ 5.61e+10    
+       0.3875798222297053
+     -0.08649404084816294
+       0.4042803834240363
+    -0.009137254536027189
+     -0.04364274600804567
+       0.4030745758661522
+     0.002511332357646316
+    -0.009157414022172862
+     -0.08610089812706949
+       0.3879203725221893
+ 5.62e+10    
+       0.3880222468073576
+     -0.08664590298516048
+       0.4048071971955488
+    -0.009127261208666379
+     -0.04376343445478716
+       0.4035991083435356
+     0.002582812160913552
+    -0.009147497457343258
+     -0.08625087220408073
+       0.3883612251999601
+ 5.63e+10    
+       0.3884634772278685
+     -0.08679755348924921
+        0.405333069043965
+    -0.009116921068456373
+     -0.04388433942587581
+       0.4041227013525238
+     0.002654579418227488
+    -0.009137233190321203
+     -0.08640062887792055
+       0.3888008721897234
+ 5.64e+10    
+       0.3889035150079078
+     -0.08694899651800921
+       0.4058579999215929
+    -0.009106234034835885
+     -0.04400546129340011
+       0.4046453560291286
+     0.002726626378217455
+     -0.00912662116845191
+     -0.08655017237830231
+        0.389239314944098
+ 5.65e+10    
+       0.3893423617396278
+     -0.08710023635010848
+       0.4063819908391734
+    -0.009095200046726893
+      -0.0441268004332005
+        0.405167073569598
+     0.002798945155280918
+     -0.00911566135961327
+      -0.0866995070569844
+       0.3896765549909996
+ 5.66e+10    
+       0.3897800190907741
+     -0.08725127738542521
+       0.4069050428660279
+    -0.009083819062500711
+     -0.04424835722494531
+       0.4056878552305522
+      0.00287152773004843
+    -0.009104353752187844
+     -0.08684863738787904
+       0.3901125939337461
+ 5.67e+10    
+       0.3902164888047839
+     -0.08740212414515681
+       0.4074271571301968
+    -0.009072091059944111
+     -0.04437013205220829
+       0.4062077023291062
+     0.002944365949883336
+    -0.009092698355034366
+     -0.08699756796714543
+       0.3905474334511528
+ 5.68e+10    
+       0.3906517727008749
+      -0.0875527812719174
+       0.4079483348185757
+    -0.009060016036225959
+     -0.04449212530254743
+       0.4067266162429927
+     0.003017451529416721
+    -0.009080695197459729
+     -0.08714630351327236
+       0.3909810752976185
+ 5.69e+10    
+        0.391085872674129
+     -0.08770325352982067
+       0.4084685771770414
+    -0.009047594007864106
+     -0.04461433736758497
+       0.4072445984106728
+     0.003090776051117162
+    -0.009068344329191107
+     -0.08729484886714618
+       0.3914135213032034
+ 5.7e+10     
+       0.3915187906955622
+     -0.08785354580455285
+       0.4089878855105741
+    -0.009034825010692455
+     -0.04473676864308992
+       0.4077616503314437
+     0.003164330965895577
+    -0.009055645820347994
+      -0.0874432089921071
+       0.3918447733736951
+ 5.71e+10    
+       0.3919505288121879
+     -0.08800366310343095
+       0.4095062611833717
+    -0.009021709099828502
+     -0.04485941952906097
+        0.408277773565538
+     0.003238107593744933
+    -0.009042599761414768
+     -0.08759138897399288
+       0.3922748334906692
+ 5.72e+10    
+       0.3923810891470708
+     -0.08815361055544918
+        0.410023705618956
+     -0.00900824634964135
+     -0.04498229042981111
+       0.4087929697342158
+     0.003312097124414989
+    -0.009029206263213178
+     -0.08773939402116861
+       0.3927037037115373
+ 5.73e+10    
+       0.3928104738993737
+      -0.0883033934113145
+        0.410540220300276
+    -0.008994436853720044
+     -0.04510538175405406
+       0.4093072405198521
+     0.003386290618121721
+    -0.009015465456875184
+     -0.08788722946454547
+       0.3931313861695866
+ 5.74e+10    
+       0.3932386853443923
+     -0.08845301704346781
+       0.4110558067698017
+    -0.008980280724842204
+     -0.04522869391499178
+       0.4098205876660163
+     0.003460679006291695
+    -0.009001377493816253
+     -0.08803490075758726
+       0.3935578830740152
+ 5.75e+10    
+       0.3936657258335828
+     -0.08860248694609425
+       0.4115704666296124
+    -0.008965778094943457
+      -0.0453522273304037
+       0.4103330129775465
+     0.003535253092341065
+    -0.008986942545708677
+     -0.08818241347630268
+       0.3939831967099507
+ 5.76e+10    
+        0.394091597794584
+     -0.08875180873512184
+       0.4120842015414778
+     -0.00895092911508708
+      -0.0454759824227369
+       0.4108445183206141
+     0.003610003552489262
+    -0.008972160804455207
+     -0.08832977331922751
+       0.3944073294384675
+ 5.77e+10    
+       0.3945163037312241
+     -0.08890098814820674
+        0.412597013226937
+    -0.008935733955434146
+     -0.04559995961919892
+       0.4113551056227868
+     0.003684920936607208
+    -0.008957032482163204
+     -0.08847698610739377
+       0.3948302836965897
+ 5.78e+10    
+       0.3949398462235267
+     -0.08905003104470789
+       0.4131089034673626
+    -0.008920192805214524
+     -0.04572415935185004
+       0.4118647768730807
+     0.003759995669099893
+    -0.008941557811119128
+     -0.08862405778428623
+       0.3952520619972906
+ 5.79e+10    
+       0.3953622279277031
+     -0.08919894340565035
+       0.4136198741040284
+    -0.008904305872697783
+     -0.04584858205769936
+       0.4123735341220096
+     0.003835218049823297
+    -0.008925737043763227
+     -0.08877099441578867
+       0.3956726669294784
+ 5.8e+10     
+       0.3957834515761382
+     -0.08934773133367432
+        0.414129927038163
+    -0.008888073385165542
+     -0.04597322817880013
+       0.4128813794816256
+     0.003910578255035648
+    -0.008909570452664613
+     -0.08891780219011686
+       0.3960921011579796
+ 5.81e+10    
+       0.3962035199773692
+     -0.08949640105297588
+       0.4146390642310004
+    -0.008871495588883347
+     -0.04609809816234805
+       0.4133883151255519
+     0.003986066338382275
+      -0.0088930583304969
+     -0.08906448741773974
+       0.3965103674235083
+ 5.82e+10    
+       0.3966224360160557
+     -0.08964495890923418
+       0.4151472877038255
+    -0.008854572749074169
+     -0.04622319246078017
+       0.4138943432890151
+     0.004061672231914898
+    -0.008876200990014167
+     -0.08921105653129033
+       0.3969274685426314
+ 5.83e+10    
+       0.3970402026529391
+      -0.0897934113695282
+       0.4156545995380108
+    -0.008837305149891563
+     -0.04634851153187561
+       0.4143994662688659
+     0.004137385747144138
+    -0.008858998764027267
+     -0.08935751608546386
+       0.3973434074077239
+ 5.84e+10    
+       0.3974568229248009
+     -0.08994176502224131
+        0.416161001875048
+    -0.008819693094394242
+     -0.04647405583885759
+       0.4149036864235947
+     0.004213196576125877
+    -0.008841452005380664
+     -0.08950387275690422
+       0.3977581869869152
+ 5.85e+10    
+       0.3978722999444058
+      -0.0900900265769556
+       0.4166664969165749
+    -0.008801736904520699
+     -0.04659982585049661
+       0.4154070061733429
+     0.004289094292580806
+    -0.008823561086929691
+     -0.08965013334408112
+       0.3981718103240329
+ 5.86e+10    
+       0.3982866369004396
+     -0.09023820286433398
+       0.4171710869243931
+    -0.008783436921064654
+     -0.04672582204121556
+       0.4159094279999071
+      0.00436506835304709
+    -0.008805326401518097
+     -0.08979630476715326
+       0.3985842805385305
+ 5.87e+10    
+       0.3986998370574445
+     -0.09038630083599297
+        0.417674774220484
+    -0.008764793503651185
+     -0.04685204489119581
+       0.4164109544467344
+     0.004441108098066113
+    -0.008786748361956292
+     -0.08994239406782201
+       0.3989956008254137
+ 5.88e+10    
+        0.399111903755739
+     -0.09053432756436269
+        0.418177561187013
+    -0.008745807030713414
+     -0.04697849488648474
+       0.4169115881189174
+     0.004517202753400728
+    -0.008767827400999871
+     -0.09008840840917391
+       0.3994057744551591
+ 5.89e+10    
+       0.3995228404113353
+     -0.09068229024253686
+       0.4186794502663332
+    -0.008726477899469795
+     -0.04710517251910482
+       0.4174113316831782
+     0.004593341431286143
+    -0.008748563971328723
+     -0.09023435507551172
+         0.39981480477362
+ 5.9e+10     
+       0.3999326505158496
+     -0.09083019618411274
+         0.41918044396098
+    -0.008706806525902264
+     -0.04723207828716397
+       0.4179101878678484
+     0.004669513131712912
+    -0.008728958545526293
+     -0.09038024147217523
+       0.4002226952019308
+ 5.91e+10    
+       0.4003413376364018
+     -0.09097805282301891
+       0.4196805448336624
+    -0.008686793344734517
+     -0.04735921269496746
+       0.4184081594628436
+     0.004745706743741892
+    -0.008709011616059702
+     -0.09052607512535021
+       0.4006294492364011
+ 5.92e+10    
+       0.4007489054155132
+     -0.09112586771333472
+       0.4201797555072436
+    -0.008666438809411646
+     -0.04748657625313089
+       0.4189052493196302
+     0.004821911046851118
+    -0.008688723695260223
+     -0.09067186368186848
+       0.4010350704484039
+ 5.93e+10    
+       0.4011553575709915
+     -0.09127364852909597
+       0.4206780786647219
+    -0.008645743392079797
+     -0.04761416947869469
+       0.4194014603511895
+     0.004898114712313712
+    -0.008668095315303829
+     -0.09081761490899598
+       0.4014395624842551
+ 5.94e+10    
+       0.4015606978958141
+     -0.09142140306409449
+       0.4211755170492013
+    -0.008624707583566669
+     -0.04774199289524023
+       0.4198967955319712
+     0.004974306304607243
+    -0.008647127028192744
+     -0.09096333669421046
+       0.4018429290650871
+ 5.95e+10    
+       0.4019649302580019
+     -0.09156913923166349
+       0.4216720734638572
+    -0.008603331893362848
+     -0.04787004703300641
+        0.420391257897848
+     0.005050474282853776
+    -0.008625819405736965
+     -0.09110903704497045
+       0.4022451739867173
+ 5.96e+10    
+       0.4023680586004849
+     -0.09171686506445553
+       0.4221677507718999
+    -0.008581616849603318
+     -0.04799833242900903
+       0.4208848505460543
+     0.005126607002290504
+    -0.008604173039536697
+     -0.09125472408847099
+       0.4026463011195053
+ 5.97e+10    
+       0.4027700869409674
+     -0.09186458871420901
+       0.4226625518965264
+     -0.00855956299904998
+     -0.04812684962716017
+        0.421377576635132
+      0.00520269271577044
+    -0.008582188540964604
+     -0.09140040607139266
+       0.4030463144082084
+ 5.98e+10    
+       0.4031710193717783
+     -0.09201231845150538
+       0.4231564798208709
+    -0.008537170907074589
+     -0.04825559917838931
+       0.4218694393848605
+     0.005278719575293196
+    -0.008559866541149052
+     -0.09154609135963854
+       0.4034452178718279
+ 5.99e+10    
+       0.4035708600597237
+     -0.09216006266551671
+       0.4236495375879495
+    -0.008514441157642202
+     -0.04838458164076643
+       0.4223604420761838
+     0.005354675633565075
+    -0.008537207690957374
+     -0.09169178843806061
+       0.4038430156034472
+ 6e+10       
+       0.4039696132459253
+     -0.09230782986374196
+       0.4241417283005969
+    -0.008491374353295552
+     -0.04851379757962531
+       0.4228505880511353
+     0.005430548845588468
+     -0.00851421266097975
+     -0.09183750591017929
+       0.4042397117700707
+ 6.01e+10    
+        0.404367283245658
+     -0.09245562867173585
+       0.4246330551213999
+    -0.008467971115139368
+     -0.04864324756768881
+       0.4233398807127522
+     0.005506327070279989
+    -0.008490882141513278
+     -0.09198325249788916
+       0.4046353106124455
+ 6.02e+10    
+       0.4047638744481803
+     -0.09260346783282676
+       0.4251235212726243
+    -0.008444232082825855
+      -0.0487729321851957
+       0.4238283235249898
+     0.005581998072117117
+    -0.008467216842546584
+      -0.0921290370411591
+       0.4050298164448874
+ 6.03e+10    
+       0.4051593913165568
+     -0.09275135620782507
+       0.4256131300361371
+    -0.008420157914540432
+     -0.04890285202002782
+       0.4243159200126235
+       0.0056575495228128
+    -0.008443217493744663
+     -0.09227486849772043
+       0.4054232336550963
+ 6.04e+10    
+       0.4055538383874783
+     -0.09289930277472383
+       0.4261018847533231
+     -0.00839574928698782
+     -0.04903300766783969
+       0.4248026737611523
+     0.005732969003017841
+    -0.008418884844434002
+     -0.09242075594274558
+       0.4058155667039616
+ 6.05e+10    
+       0.4059472202710725
+     -0.09304731662838735
+       0.4265897888249939
+    -0.008371006895378985
+     -0.04916339973218839
+       0.4252885884166934
+     0.005808244004050376
+    -0.008394219663588123
+     -0.09256670856851931
+       0.4062068201253729
+ 6.06e+10    
+       0.4063395416507116
+     -0.09319540698023351
+       0.4270768457112962
+    -0.008345931453418184
+     -0.04929402882466525
+       0.4257736676858711
+     0.005883361929652395
+    -0.008369222739813416
+       -0.092712735684099
+        0.406596998526011
+ 6.07e+10    
+       0.4067308072828135
+     -0.09334358315790539
+        0.427563058931612
+    -0.008320523693290765
+     -0.04942489556502896
+       0.4262579153357026
+     0.005958310097772633
+    -0.008343894881335044
+     -0.09285884671496648
+       0.4069861065851459
+ 6.08e+10    
+       0.4071210219966377
+     -0.09349185460493455
+       0.4280484320644521
+    -0.008294784365651037
+     -0.04955600058133928
+       0.4267413351934753
+     0.006033075742375332
+    -0.008318236915983355
+     -0.09300505120267086
+        0.407374149054422
+ 6.09e+10    
+       0.4075101906940765
+     -0.09364023088039468
+       0.4285329687473474
+    -0.008268714239610944
+     -0.04968734451009232
+       0.4272239311466249
+     0.006107646015274713
+    -0.008292249691180142
+     -0.09315135880446251
+       0.4077611307576385
+ 6.1e+10     
+       0.4078983183494381
+     -0.09378872165854761
+       0.4290166726767333
+    -0.008242314102728823
+     -0.04981892799635756
+       0.4277057071426011
+     0.006182007987994622
+    -0.008265934073925623
+     -0.09329777929291863
+       0.4081470565905284
+ 6.11e+10    
+       0.4082854100092302
+     -0.09393733672848051
+       0.4294995476078318
+    -0.008215584760998557
+     -0.04995075169391518
+       0.4281866671887327
+     0.006256148653652685
+    -0.008239290950784971
+     -0.09344432255555873
+        0.408531931520528
+ 6.12e+10    
+       0.4086714707919328
+     -0.09408608599373325
+       0.4299815973545223
+    -0.008188527038838902
+     -0.05008281626539522
+       0.4286668153520862
+     0.006330054928868626
+    -0.008212321227875383
+     -0.09359099859445318
+       0.4089157605865424
+ 6.13e+10    
+       0.4090565058877688
+     -0.09423497947191892
+       0.4304628257892144
+      -0.0081611417790836
+     -0.05021512238241765
+       0.4291461557593211
+     0.006403713655696551
+    -0.008185025830853282
+     -0.09373781752582258
+         0.40929854889871
+ 6.14e+10    
+       0.4094405205584706
+     -0.09438402729433593
+       0.4309432368427124
+    -0.008133429842971064
+      -0.0503476707257337
+       0.4296246925965379
+       0.0064771116035804
+    -0.008157405704901121
+     -0.09388478957962901
+       0.4096803016381549
+ 6.15e+10    
+        0.409823520137041
+     -0.09453323970556961
+       0.4314228345040745
+    -0.008105392110134734
+     -0.05048046198536884
+       0.4301024301091228
+     0.006550235471331843
+    -0.008129461814714755
+     -0.09403192509915825
+       0.4100610240567413
+ 6.16e+10    
+       0.4102055100275078
+     -0.09468262706308908
+       0.4319016228204681
+    -0.008077029478593421
+     -0.05061349686076605
+       0.4305793726015865
+     0.006623071889130869
+    -0.008101195144490439
+     -0.09417923454059481
+       0.4104407214768184
+ 6.17e+10    
+       0.4105864957046771
+     -0.09483219983683325
+       0.4323796058970201
+    -0.008048342864741957
+     -0.05074677606093073
+       0.4310555244374003
+     0.006695607420548047
+    -0.008072606697912169
+     -0.09432672847258872
+       0.4108193992909663
+ 6.18e+10    
+       0.4109664827138811
+     -0.09498196860879085
+       0.4328567878966632
+    -0.008019333203341574
+     -0.05088030030457736
+       0.4315308900388242
+     0.006767828564587741
+    -0.008043697498138453
+      -0.0944744175758138
+       0.4111970629617289
+ 6.19e+10    
+       0.4113454766707189
+     -0.09513194407257065
+       0.4333331730399753
+    -0.007990001447510962
+     -0.05101407032027559
+       0.4320054738867309
+     0.006839721757752365
+    -0.008014468587789458
+     -0.09462231264251773
+       0.4115737180213523
+ 6.2e+10     
+       0.4117234832607986
+     -0.09528213703296594
+       0.4338087656050154
+    -0.007960348568716802
+     -0.05114808684659972
+       0.4324792805204315
+     0.006911273376126773
+    -0.007984921028933601
+     -0.09477042457606709
+       0.4119493700715114
+ 6.21e+10    
+       0.4121005082394701
+     -0.09543255840551038
+       0.4342835699271582
+    -0.007930375556764551
+     -0.05128235063227753
+       0.4329523145374856
+     0.006982469737482297
+    -0.007955055903074375
+     -0.09491876439048086
+       0.4123240247830363
+ 6.22e+10    
+       0.4124765574315559
+     -0.09558321921602519
+       0.4347575903989154
+    -0.007900083419789082
+     -0.05141686243634064
+       0.4334245805935144
+     0.007053297103399714
+    -0.007924874311136573
+     -0.09506734320995858
+       0.4126976878956337
+ 6.23e+10    
+       0.4128516367310789
+     -0.09573413060016156
+       0.4352308314697636
+    -0.007869473184245338
+     -0.05155162302827704
+         0.43389608340201
+      0.00712374168141134
+    -0.007894377373452372
+     -0.09521617226840137
+       0.4130703652176029
+ 6.24e+10    
+       0.4132257521009858
+     -0.09588530380293311
+       0.4357032976459576
+    -0.007838545894898777
+     -0.05168663318818289
+       0.4343668277341334
+     0.007193789627160472
+    -0.007863566229747265
+     -0.09536526290892451
+       0.4134420626255514
+ 6.25e+10    
+       0.4135989095728656
+     -0.09603675017824299
+       0.4361749934903471
+    -0.007807302614815497
+      -0.0518218937069171
+       0.4348368184185167
+     0.007263427046578903
+    -0.007832442039125382
+     -0.09551462658336354
+       0.4138127860641041
+ 6.26e+10    
+       0.4139711152466659
+     -0.09618848118840154
+       0.4366459236221829
+    -0.007775744425352687
+     -0.05195740538625564
+       0.4353060603410532
+     0.007332639998081029
+    -0.007801005980054611
+     -0.09566427485177205
+       0.4141825415456066
+ 6.27e+10    
+       0.4143423752904066
+     -0.09634050840364024
+        0.437116092716923
+    -0.007743872426147753
+     -0.05209316903904795
+       0.4357745584446873
+     0.007401414494774364
+    -0.007769259250351204
+     -0.09581421938191406
+       0.4145513351498333
+ 6.28e+10    
+       0.4147126959398876
+     -0.09649284350161517
+       0.4375855055060323
+    -0.007711687735108468
+     -0.05222918548937398
+       0.4362423177292021
+     0.007469736506685818
+    -0.007737203067163822
+     -0.09596447194874907
+        0.414919173023682
+ 6.29e+10    
+        0.415082083498393
+     -0.09664549826690552
+       0.4380541667767778
+    -0.007679191488401472
+      -0.0523654555727018
+       0.4367093432509959
+     0.007537591963003309
+    -0.007704838666957238
+     -0.09611504443390839
+       0.4152860613808715
+ 6.3e+10     
+       0.4154505443363982
+     -0.09679848459050561
+        0.438522081372022
+     -0.00764638484044136
+     -0.05250198013604733
+       0.4371756401228618
+      0.00760496675433176
+    -0.007672167305495182
+     -0.09626594882516748
+       0.4156520065016351
+ 6.31e+10    
+       0.4158180848912648
+      -0.0969518144693087
+       0.4389892541900086
+    -0.007613268963878617
+      -0.0526387600381338
+        0.437641213513758
+      0.00767184673496326
+    -0.007639190257822861
+     -0.09641719721590966
+       0.4160170147324085
+ 6.32e+10    
+       0.4161847116669396
+     -0.09710550000558567
+       0.4394556901841468
+    -0.007579845049587494
+     -0.05277579614955363
+       0.4381060686485785
+     0.007738217725160716
+     -0.00760590881824857
+     -0.09656880180458458
+       0.4163810924855177
+ 6.33e+10    
+       0.4165504312336464
+     -0.09725955340645573
+       0.4399213943627883
+    -0.007546114306652913
+     -0.05291308935292958
+       0.4385702108079141
+     0.007804065513454003
+    -0.007572324300324586
+     -0.09672077489415865
+       0.4167442462388614
+ 6.34e+10    
+       0.4169152502275792
+     -0.09741398698335328
+       0.4403863717890067
+    -0.007512077962357197
+     -0.05305064054307859
+       0.4390336453278146
+     0.007869375858948844
+    -0.007538438036827515
+     -0.09687312889156072
+        0.417106482535593
+ 6.35e+10    
+       0.4172791753505868
+      -0.0975688131514845
+       0.4408506275803654
+    -0.007477737262165797
+     -0.05318845062717576
+       0.4394963775995452
+     0.007934134493646876
+    -0.007504251379737471
+     -0.09702587630712095
+       0.4174678079837975
+ 6.36e+10    
+       0.4176422133698608
+     -0.09772404442928165
+       0.4413141669086845
+    -0.007443093469712322
+     -0.05332652052491896
+       0.4399584130693378
+     0.007998327124776938
+    -0.007469765700216639
+     -0.09717902975400299
+       0.4178282292561676
+ 6.37e+10    
+       0.4180043711176165
+     -0.09787969343784862
+        0.441776994999806
+     -0.00740814786678301
+     -0.05346485116869522
+         0.44041975723814
+     0.008061939437136683
+    -0.007434982388586694
+     -0.09733260194763049
+       0.4181877530896757
+ 6.38e+10    
+       0.4183656554907743
+     -0.09803577290040207
+       0.4422391171333524
+    -0.007372901753300025
+      -0.0536034435037474
+       0.4408804156613595
+     0.008124957095443999
+    -0.007399902854305499
+     -0.09748660570510773
+       0.4185463862852444
+ 6.39e+10    
+       0.4187260734506372
+      -0.0981922956417051
+       0.4427005386424819
+    -0.007337356447304341
+     -0.05374229848834221
+       0.4413403939486055
+     0.008187365746697647
+    -0.007364528525942344
+     -0.09764105394463443
+       0.4189041357074148
+ 6.4e+10     
+       0.4190856320225662
+     -0.09834927458749676
+       0.4431612649136397
+    -0.007301513284937064
+     -0.05388141709393864
+       0.4417996977634253
+     0.008249151022546281
+    -0.007328860851152596
+     -0.09779595968491492
+       0.4192610082840124
+ 6.41e+10    
+       0.4194443382956539
+     -0.09850672276391402
+       0.4436213013863078
+    -0.007265373620420388
+     -0.05402080030535789
+       0.4422583328230377
+     0.008310298541665585
+    -0.007292901296650778
+     -0.09795133604455977
+       0.4196170110058082
+ 6.42e+10    
+       0.4198021994223949
+     -0.09866465329690928
+       0.4440806535527471
+    -0.007228938826037022
+     -0.05416044912095385
+       0.4427163048980636
+     0.008370793912142535
+     -0.00725665134818262
+     -0.09810719624148537
+       0.4199721509261841
+ 6.43e+10    
+       0.4201592226183561
+     -0.09882307941166228
+       0.4445393269577402
+    -0.007192210292108722
+      -0.0543003645527844
+        0.443173619812252
+     0.008430622733866409
+    -0.007220112510495849
+     -0.09826355359230479
+       0.4203264351607868
+ 6.44e+10    
+       0.4205154151618433
+     -0.09898201443198551
+       0.4449973271983272
+    -0.007155189426973545
+     -0.05444054762678384
+       0.4436302834422025
+     0.008489770600925702
+    -0.007183286307309673
+     -0.09842042151171411
+       0.4206798708871894
+ 6.45e+10    
+       0.4208707843935666
+     -0.09914147177972547
+       0.4454546599235393
+    -0.007117877656962153
+     -0.05458099938293557
+        0.444086301717084
+     0.008548223104010814
+    -0.007146174281282789
+     -0.09857781351187472
+       0.4210324653445449
+ 6.46e+10    
+       0.4212253377163038
+     -0.09930146497415775
+       0.4459113308341289
+    -0.007080276426372357
+     -0.05472172087544667
+       0.4445416806183527
+     0.008605965832820918
+    -0.007108777993980014
+     -0.09873574320178904
+       0.4213842258332405
+ 6.47e+10    
+       0.4215790825945631
+     -0.09946200763137651
+       0.4463673456822964
+    -0.007042387197442756
+     -0.05486271317292216
+       0.4449964261794618
+     0.008662984378475427
+     -0.00707109902583745
+     -0.09889422428667048
+       0.4217351597145476
+ 6.48e+10    
+       0.4219320265542419
+     -0.09962311346368113
+       0.4468227102714151
+     -0.00700421145032463
+     -0.05500397735854103
+        0.445450544485573
+     0.008719264335928891
+    -0.007033138976126261
+     -0.09905327056731095
+       0.4220852744102757
+ 6.49e+10    
+       0.4222841771822861
+     -0.09978479627895363
+       0.4472774304557459
+    -0.006965750683052671
+     -0.05514551453023213
+       0.4459040416732605
+     0.008774791306388389
+    -0.006994899462914326
+     -0.09921289593944017
+       0.4224345774024162
+ 6.5e+10     
+       0.4226355421263471
+     -0.09994706998003544
+       0.4477315121401591
+    -0.006927006411514084
+     -0.05528732580085179
+       0.4463569239302147
+     0.008829550899733748
+    -0.006956382123026943
+     -0.09937311439308263
+       0.4227830762327949
+ 6.51e+10    
+       0.4229861290944374
+      -0.1001099485640969
+       0.4481849612798452
+      -0.0068879801694159
+     -0.05542941229836126
+       0.4468091974949408
+     0.008883528736938869
+    -0.006917588612005343
+     -0.09953394001190835
+       0.4231307785027137
+ 6.52e+10    
+       0.4233359458545861
+      -0.1002734461220022
+       0.4486377838800253
+    -0.006848673508250989
+     -0.05557177516600619
+       0.4472608686564558
+     0.008936710452494136
+    -0.006878520604063318
+     -0.09969538697257968
+        0.423477691872597
+ 6.53e+10    
+       0.4236850002344901
+      -0.1004375768376699
+        0.449089985995657
+    -0.006809087997262153
+     -0.05571441556249528
+       0.4477119437539817
+      0.00898908169682925
+    -0.006839179792042691
+      -0.0998574695440928
+       0.4238238240616347
+ 6.54e+10    
+       0.4240333001211672
+      -0.1006023549874288
+        0.449541573731139
+    -0.006769225223404585
+     -0.05585733466218084
+       0.4481624291766336
+     0.009040628138735671
+     -0.00679956788736602
+      -0.1000202020871153
+       0.4241691828474239
+ 6.55e+10    
+       0.4243808534606059
+      -0.1007677949393686
+       0.4499925532400104
+    -0.006729086791306377
+      -0.0560005336552395
+       0.4486123313631087
+     0.009091335467788056
+    -0.006759686619988147
+      -0.1001835990533189
+       0.4245137760656105
+ 6.56e+10    
+       0.4247276682574178
+      -0.1009339111526885
+       0.4504429307246502
+     -0.00668867432322726
+     -0.05614401374785418
+       0.4490616568013703
+     0.009141189396764228
+    -0.006719537738345128
+      -0.1003476749847083
+       0.4248576116095287
+ 6.57e+10    
+       0.4250737525744827
+      -0.1011007181770372
+       0.4508927124359698
+    -0.006647989459015388
+     -0.05628777616239605
+       0.4495104120283273
+     0.009190175664062879
+    -0.006679123009301515
+      -0.1005124445129453
+       0.4252006974298412
+ 6.58e+10    
+       0.4254191145325987
+      -0.1012682306518523
+       0.4513419046731046
+    -0.006607033856062179
+     -0.05643182213760753
+       0.4499586036295136
+      0.00923828003611829
+     -0.00663844421809528
+      -0.1006779223586682
+       0.4255430415341753
+ 6.59e+10    
+        0.425763762310128
+      -0.1014364633056938
+        0.451790513783104
+    -0.006565809189254859
+     -0.05657615292878608
+       0.4504062382387642
+     0.009285488309811898
+    -0.006597503168280726
+      -0.1008441233308092
+       0.4258846519867611
+ 6.6e+10     
+       0.4261077041426457
+      -0.1016054309555745
+        0.452238546160615
+    -0.006524317150927415
+     -0.05672076980796818
+       0.4508533225378857
+     0.009331786314879457
+    -0.006556301681669187
+      -0.1010110623259048
+       0.4262255369080696
+ 6.61e+10    
+       0.4264509483225797
+      -0.1017751485062835
+       0.4526860082475654
+    -0.006482559450808688
+     -0.05686567406411448
+        0.451299863256328
+     0.009377159916313559
+    -0.006514841598267006
+      -0.1011787543274044
+       0.4265657044744455
+ 6.62e+10    
+       0.4267935031988632
+       -0.101945630949711
+       0.4531329065328475
+    -0.006440537815968794
+     -0.05701086700329565
+       0.4517458671708497
+     0.009421595016760976
+    -0.006473124776212019
+      -0.1013472144049748
+       0.4269051629177462
+ 6.63e+10    
+       0.4271353771765717
+      -0.1021168933641627
+       0.4535792475519884
+    -0.006398253990763161
+     -0.05715634994887746
+       0.4521913411051846
+     0.009465077558913789
+    -0.006431153091706665
+         -0.1015164577138
+       0.4272439205249727
+ 6.64e+10    
+       0.4274765787165704
+      -0.1022889509136761
+       0.4540250378868303
+    -0.006355709736773964
+      -0.0573021242417088
+       0.4526362919297028
+     0.009507593527894103
+    -0.006388928438949485
+      -0.1016864994938782
+       0.4275819856379072
+ 6.65e+10    
+       0.4278171163351574
+      -0.1024618188473292
+       0.4544702841651996
+    -0.006312906832749304
+     -0.05744819124030777
+       0.4530807265610667
+     0.009549128953631383
+      -0.0063464527300635
+      -0.1018573550693137
+        0.427919366652744
+ 6.66e+10    
+       0.4281569986037049
+      -0.1026355124985475
+       0.4549149930605786
+    -0.006269847074540226
+     -0.05759455232105094
+       0.4535246519618952
+     0.009589669913232271
+    -0.006303727895022338
+      -0.1020290398476083
+       0.4282560720197241
+ 6.67e+10    
+       0.4284962341483027
+      -0.1028100472844071
+       0.4553591712917695
+    -0.006226532275034644
+     -0.05774120887836012
+       0.4539680751404099
+      0.00962920253334193
+    -0.006260755881573876
+      -0.1022015693189459
+       0.4285921102427694
+ 6.68e+10    
+       0.4288348316494003
+      -0.1029854387049329
+       0.4558028256225591
+    -0.006182964264089322
+     -0.05788816232489231
+        0.454411003150091
+     0.009667712992495948
+    -0.006217538655160755
+      -0.1023749590554747
+        0.428927489879113
+ 6.69e+10    
+       0.4291727998414468
+      -0.1031617023423956
+       0.4562459628613815
+     -0.00613914488845865
+     -0.05803541409172908
+       0.4548534430893284
+     0.009705187523463178
+    -0.006174078198838489
+      -0.1025492247105886
+       0.4292622195389344
+ 6.7e+10     
+       0.4295101475125351
+      -0.1033388538606034
+       0.4566885898609787
+    -0.006095076011721212
+     -0.05818296562856663
+       0.4552954021010637
+     0.009741612415578244
+     -0.00613037651319079
+      -0.1027243820182005
+       0.4295963078849893
+ 6.71e+10    
+       0.4298468835040426
+      -0.1035169090041919
+       0.4571307135180523
+    -0.006050759514203558
+     -0.05833081840390508
+       0.4557368873724395
+     0.009776974017062933
+    -0.006086435616242164
+      -0.1029004467920175
+       0.4299297636322436
+ 6.72e+10    
+       0.4301830167102697
+      -0.1036958835979085
+       0.4575723407729227
+    -0.006006197292900728
+     -0.05847897390524082
+       0.4561779061344403
+     0.009811258737336542
+    -0.006042257543367117
+        -0.10307743492481
+       0.4302625955475058
+ 6.73e+10    
+       0.4305185560780863
+      -0.1038757935458977
+       0.4580134786091815
+    -0.005961391261394642
+     -0.05862743363925715
+       0.4566184656615311
+     0.009844453049314326
+    -0.005997844347197341
+      -0.1032553623876773
+       0.4305948124490582
+ 6.74e+10    
+       0.4308535106065673
+       -0.104056654830978
+       0.4584541340533358
+    -0.005916343349769124
+     -0.05877619913201571
+       0.4570585732712996
+     0.009876543491692917
+    -0.005953198097524695
+       -0.103434245229314
+       0.4309264232062894
+ 6.75e+10    
+       0.4311878893466388
+      -0.1042384835139208
+       0.4588943141744633
+     -0.00587105550452204
+     -0.05892527192914956
+       0.4574982363240871
+     0.009907516671223075
+    -0.005908320881202556
+      -0.1036140995752683
+        0.431257436739326
+ 6.76e+10    
+       0.4315217014007146
+       -0.104421295732723
+       0.4593340260838532
+    -0.005825529688474712
+     -0.05907465359605515
+       0.4579374622226273
+     0.009937359264968868
+    -0.005863214802042932
+      -0.1037949416272028
+       0.4315878620186684
+ 6.77e+10    
+       0.4318549559223424
+      -0.1046051077018776
+       0.4597732769346489
+    -0.005779767880678081
+     -0.05922434571808514
+       0.4583762584116755
+     0.009966058022552012
+    -0.005817881980710959
+      -0.1039767876621483
+       0.4319177080648184
+ 6.78e+10    
+       0.4321876621158425
+      -0.1047899357116433
+        0.460212073921492
+     -0.00573377207631569
+      -0.0593743499007419
+       0.4588146323776362
+     0.009993599768382122
+    -0.005772324554616437
+       -0.104159654031757
+       0.4322469839479156
+ 6.79e+10    
+       0.4325198292359493
+      -0.1049757961273081
+         0.46065042428016
+    -0.005687544286603894
+     -0.05952466776987164
+       0.4592525916481972
+      0.01001997140387111
+    -0.005726544677801629
+      -0.1043435571615541
+       0.4325756987873697
+ 6.8e+10     
+       0.4328514665874547
+      -0.1051627053884533
+       0.4610883352872031
+    -0.005641086538688386
+     -0.05967530097185772
+       0.4596901437919486
+      0.01004515990963191
+     -0.00568054452082618
+      -0.1045285135501836
+       0.4329038617514931
+ 6.81e+10    
+       0.4331825835248497
+      -0.1053506800082127
+       0.4615258142595799
+    -0.005594400875538201
+     -0.05982625117381509
+       0.4601272964180116
+      0.01006915234766092
+    -0.005634326270648705
+      -0.1047145397686557
+       0.4332314820571369
+ 6.82e+10    
+       0.4335131894519672
+      -0.1055397365725314
+       0.4619628685542911
+    -0.005547489355835485
+      -0.0599775200637858
+       0.4605640571756603
+      0.01009193586350325
+    -0.005587892130504757
+      -0.1049016524595891
+       0.4335585689693215
+ 6.83e+10    
+       0.4338432938216247
+      -0.1057298917394195
+       0.4623995055680091
+    -0.005500354053863078
+     -0.06012910935093251
+       0.4610004337539385
+      0.01011349768840063
+     -0.00554124431978173
+      -0.1050898683364511
+       0.4338851318008741
+ 6.84e+10    
+       0.4341729061352674
+      -0.1059211622382059
+       0.4628357327367088
+    -0.005452997059387735
+      -0.0602810207657344
+       0.4614364338812824
+      0.01013382514142123
+    -0.005494385073890313
+       -0.105279204182798
+       0.4342111799120638
+ 6.85e+10    
+       0.4345020359426136
+       -0.106113564868789
+       0.4632715575352955
+    -0.005405420477540571
+     -0.06043325606018281
+       0.4618720653251364
+      0.01015290563157128
+    -0.005447316644132153
+        -0.10546967685151
+       0.4345367227102345
+ 6.86e+10    
+       0.4348306928412955
+      -0.1063071165008837
+       0.4637069874772276
+    -0.005357626428693946
+     -0.06058581700797611
+       0.4623073358915675
+      0.01017072665988732
+    -0.005400041297564367
+       -0.105661303264026
+       0.4348617696494435
+ 6.87e+10    
+       0.4351588864765062
+      -0.1065018340732687
+        0.464142030114146
+    -0.005309617048334459
+     -0.06073870540471631
+       0.4627422534248779
+       0.0101872758215091
+    -0.005352561316860391
+      -0.1058541004095762
+       0.4351863302300969
+ 6.88e+10    
+       0.4354866265406465
+      -0.1066977345930301
+       0.4645766930354919
+    -0.005261394486933214
+     -0.06089192306810447
+       0.4631768258072217
+       0.0102025408077327
+    -0.005304879000167181
+      -0.1060480853444129
+        0.435510413998587
+ 6.89e+10    
+       0.4358139227729667
+      -0.1068948351348034
+       0.4650109838681303
+     -0.00521296090981186
+     -0.06104547183813732
+       0.4636110609582095
+      0.01021650940804298
+    -0.005256996660958954
+      -0.1062432751910385
+       0.4358340305469308
+ 6.9e+10     
+       0.4361407849592147
+      -0.1070931528400125
+       0.4654449102759667
+    -0.005164318497005197
+     -0.06119935357730318
+       0.4640449668345215
+      0.01022916951212491
+    -0.005208916627887049
+       -0.106439687137432
+       0.4361571895124058
+ 6.91e+10    
+       0.4364672229312825
+      -0.1072927049161094
+        0.465878479959567
+    -0.005115469443120364
+     -0.06135357017077882
+       0.4644785514295132
+      0.01024050911185417
+    -0.005160641244626401
+      -0.1066373384362753
+        0.436479900577194
+ 6.92e+10    
+       0.4367932465668565
+      -0.1074935086358092
+        0.466311700655771
+    -0.005066415957192242
+     -0.06150812352662555
+        0.464911822772821
+      0.01025051630326508
+     -0.00511217286971798
+      -0.1068362464041752
+       0.4368021734680163
+ 6.93e+10    
+       0.4371188657890596
+      -0.1076955813363243
+       0.4667445801373103
+    -0.005017160262535043
+     -0.06166301557598666
+       0.4653447889299696
+      0.01025917928849688
+    -0.005063513876407853
+      -0.1070364284208861
+       0.4371240179557768
+ 6.94e+10    
+       0.4374440905661061
+      -0.1078989404185989
+       0.4671771262124181
+    -0.004967704596590402
+      -0.0618182482732834
+       0.4657774580019726
+      0.01026648637771699
+    -0.005014666652482117
+      -0.1072379019285298
+       0.4374454438552015
+ 6.95e+10    
+        0.437768930910947
+      -0.1081036033465372
+       0.4676093467244422
+    -0.004918051210771554
+      -0.0619738235964118
+       0.4662098381249346
+      0.01027242599102091
+    -0.004965633600098219
+      -0.1074406844308145
+       0.4377664610244834
+ 6.96e+10    
+       0.4380933968809221
+      -0.1083095876462351
+       0.4680412495514541
+    -0.004868202370303774
+     -0.06212974354694006
+       0.4666419374696528
+       0.0102769866603091
+    -0.004916417135612549
+      -0.1076447934922516
+       0.4380870793649209
+ 6.97e+10    
+       0.4384174985774104
+      -0.1085169109052073
+       0.4684728426058612
+    -0.004818160354061097
+      -0.0622860101503051
+        0.467073764241218
+      0.01028015703113923
+      -0.0048670196894039
+      -0.1078502467373725
+       0.4384073088205662
+ 6.98e+10    
+       0.4387412461454805
+      -0.1087255907716133
+       0.4689041338340094
+    -0.004767927454398998
+     -0.06244262545600917
+       0.4675053266786097
+      0.01028192586455451
+    -0.004817443705693309
+      -0.1080570618499425
+       0.4387271593778664
+ 6.99e+10    
+       0.4390646497735467
+      -0.1089356449534838
+       0.4693351312157943
+    -0.004717505976983383
+     -0.06259959153781679
+        0.467936633054294
+      0.01028228203888668
+    -0.004767691642359936
+      -0.1082652565721748
+       0.4390466410653109
+ 7e+10       
+       0.4393877196930168
+      -0.1091470912179421
+        0.469765842764262
+    -0.004666898240615838
+     -0.06275691049395155
+       0.4683676916738226
+      0.01028121455153443
+    -0.004717765970752869
+      -0.1084748487039423
+        0.439365763953075
* NOTE: Solution at 1e+08 Hz used as DC point.

.model c_m4lines_port_1 sp N=4 SPACING=nonuniform VALTYPE=real
+ INTERPOLATION=spline
+ INFINITY =
+    8.016335543513601e-11
+   -2.300565173929285e-11
+    8.459718257292866e-11
+   -1.858265556210685e-12
+   -1.176346435114431e-11
+    8.452718514577025e-11
+    -1.86120549715101e-13
+    -1.84837363016514e-12
+   -2.301064440037953e-11
+    8.022553825614561e-11
+ DATA = 700
+ 0           
+    8.745714244497287e-11
+   -2.212814696889387e-11
+    8.927795692543775e-11
+   -8.467390817336624e-13
+   -1.048600945697321e-11
+    8.923543991764458e-11
+   -3.056330636422667e-13
+   -8.444772721076193e-13
+    -2.21803936465989e-11
+    8.759868115078844e-11
+ 2e+08       
+    8.683981392535683e-11
+   -2.200610203744423e-11
+    8.865513547495764e-11
+   -8.494939034760619e-13
+    -1.04321586716866e-11
+    8.861454644671484e-11
+   -3.052161253392888e-13
+   -8.472590182311929e-13
+     -2.2058071082135e-11
+     8.69799168290736e-11
+ 3e+08       
+    8.647525050009691e-11
+   -2.193547403342267e-11
+    8.828622373626237e-11
+   -8.469204314857208e-13
+   -1.040316282563671e-11
+    8.824622959178165e-11
+   -3.049158301918048e-13
+   -8.446456594881739e-13
+    -2.19877000464908e-11
+    8.661460833346853e-11
+ 4e+08       
+    8.623566605767624e-11
+   -2.189167439600001e-11
+    8.804463576155199e-11
+   -8.448921161832739e-13
+   -1.038496658518787e-11
+    8.800522489309862e-11
+   -3.048357076443738e-13
+   -8.425865898003304e-13
+   -2.194417626792234e-11
+    8.637458088434692e-11
+ 5e+08       
+    8.604953077068542e-11
+   -2.185681704418195e-11
+    8.785704659641704e-11
+   -8.436368351604128e-13
+   -1.037005385747412e-11
+    8.781815822793378e-11
+   -3.045879012637334e-13
+   -8.413140052860127e-13
+    -2.19094605598687e-11
+    8.618808448728736e-11
+ 6e+08       
+    8.589372068966307e-11
+   -2.182653721677049e-11
+     8.76998447419683e-11
+   -8.427176211337245e-13
+   -1.035688506685164e-11
+    8.766139050926989e-11
+   -3.041153998269266e-13
+   -8.403829602404814e-13
+   -2.187924950232326e-11
+    8.603195612301891e-11
+ 7e+08       
+     8.57598122801371e-11
+   -2.179984363425893e-11
+    8.756453181240886e-11
+   -8.418533659551775e-13
+   -1.034515623839089e-11
+    8.752642230455287e-11
+    -3.03463223417793e-13
+   -8.395083712774953e-13
+   -2.185259386081025e-11
+    8.589776624328757e-11
+ 8e+08       
+    8.564348177330895e-11
+   -2.177629106933934e-11
+    8.744683943305225e-11
+   -8.409249137093704e-13
+   -1.033470397950519e-11
+    8.740900612646088e-11
+   -3.026868291132039e-13
+   -8.385697085701523e-13
+   -2.182906822074987e-11
+    8.578118912466996e-11
+ 9e+08       
+    8.554159737698257e-11
+   -2.175542053672015e-11
+    8.734372730336448e-11
+   -8.399001522957813e-13
+    -1.03253364205605e-11
+    8.730613667976507e-11
+   -3.018273746429759e-13
+   -8.375342817074133e-13
+   -2.180822378326449e-11
+    8.567909055315986e-11
+ 1e+09       
+    8.545151646626288e-11
+   -2.173673192754379e-11
+    8.725264117104621e-11
+   -8.387833104678768e-13
+   -1.031684463534174e-11
+    8.721530021783062e-11
+   -3.009101086466027e-13
+   -8.364058188026178e-13
+   -2.178956708964096e-11
+    8.558882477052716e-11
+ 1.1e+09     
+    8.537898684230445e-11
+    -2.17250289549019e-11
+    8.718016701559234e-11
+   -8.379326921102572e-13
+   -1.031137362032845e-11
+    8.714292497629194e-11
+    -2.99728627197578e-13
+   -8.355709999745456e-13
+     -2.1777558421059e-11
+    8.551602498428931e-11
+ 1.2e+09     
+    8.530991664075069e-11
+   -2.171283490931975e-11
+     8.71109648362162e-11
+   -8.370169156267862e-13
+   -1.030563165598015e-11
+    8.707387941349606e-11
+   -2.986212640198248e-13
+   -8.346546581294013e-13
+    -2.17652013500883e-11
+    8.544674652982053e-11
+ 1.3e+09     
+    8.524448994759453e-11
+   -2.170034610463755e-11
+    8.704523678216632e-11
+   -8.360043977962049e-13
+     -1.0299707149649e-11
+    8.700834259445373e-11
+    -2.97559669987812e-13
+   -8.336301353214107e-13
+   -2.175265164527196e-11
+    8.538115859298584e-11
+ 1.4e+09     
+    8.518271800351701e-11
+   -2.168771953874187e-11
+    8.698301166314085e-11
+   -8.348743072902544e-13
+   -1.029366915282903e-11
+    8.694632484125158e-11
+   -2.965119320370415e-13
+   -8.324805897899816e-13
+   -2.174003368960054e-11
+    8.531926004313905e-11
+ 1.5e+09     
+    8.512450165085572e-11
+   -2.167507682931222e-11
+    8.692420692583323e-11
+   -8.336154288146159e-13
+    -1.02875700484498e-11
+    8.688772959530574e-11
+   -2.954460177243315e-13
+   -8.311978655508551e-13
+   -2.172744400223442e-11
+    8.526094189999991e-11
+ 1.6e+09     
+    8.506967620580454e-11
+    -2.16625096977916e-11
+    8.686867346366327e-11
+   -8.322243464882864e-13
+   -1.028144876688317e-11
+    8.683239771360742e-11
+    -2.94332383058791e-13
+   -8.297807807787198e-13
+   -2.171495565790221e-11
+    8.520603193610958e-11
+ 1.7e+09     
+    8.501804237008339e-11
+   -2.165008559439032e-11
+    8.681622661163894e-11
+   -8.307034980514443e-13
+   -1.027533383673226e-11
+    8.678013780777862e-11
+   -2.931457848410413e-13
+   -8.282333235948307e-13
+   -2.170262268529723e-11
+    8.515432521752572e-11
+ 1.8e+09     
+    8.496938673087429e-11
+   -2.163785279049889e-11
+     8.67666667483444e-11
+   -8.290593986251667e-13
+   -1.026924598002589e-11
+    8.673074618651991e-11
+   -2.918663800848116e-13
+   -8.265630194493905e-13
+   -2.169048400827098e-11
+    8.510560422876009e-11
+ 1.9e+09     
+    8.492349483062859e-11
+   -2.162584469326755e-11
+    8.671979243937185e-11
+   -8.273011651355911e-13
+   -1.026320018434433e-11
+    8.668401940158791e-11
+   -2.904802158404028e-13
+   -8.247795846803485e-13
+    -2.16785667781403e-11
+    8.505965160706877e-11
+ 2e+09       
+    8.488015910825542e-11
+   -2.161408336005197e-11
+    8.667540841614634e-11
+   -8.254393723244762e-13
+   -1.025720729066194e-11
+    8.663976171575178e-11
+   -2.889792229659743e-13
+    -8.22893891058683e-13
+   -2.166688909394214e-11
+    8.501625780211266e-11
+ 2.1e+09     
+    8.483918339608241e-11
+   -2.160258229079561e-11
+    8.663333008275045e-11
+    -8.23485217469477e-13
+    -1.02512751755477e-11
+     8.65977891881443e-11
+     -2.8736083079883e-13
+   -8.209172178465309e-13
+   -2.165546217386383e-11
+     8.49752253455925e-11
+ 2.2e+09     
+     8.48003851613135e-11
+   -2.159134861039139e-11
+    8.659338575105291e-11
+   -8.214499464303783e-13
+    -1.02454096125149e-11
+    8.655793156983831e-11
+   -2.856273170058236e-13
+   -8.188607459768791e-13
+   -2.164429206272162e-11
+    8.493637091363693e-11
+ 2.3e+09     
+    8.476359630903524e-11
+   -2.158038475453176e-11
+    8.655541743082014e-11
+   -8.193444864280508e-13
+   -1.023961488868521e-11
+    8.652003282488664e-11
+   -2.837849982857724e-13
+    -8.16735242711909e-13
+   -2.163338096011042e-11
+    8.489952599110291e-11
+ 2.4e+09     
+    8.472866309699911e-11
+   -2.156968976028921e-11
+    8.651928073126006e-11
+   -8.171792332576831e-13
+    -1.02338942394685e-11
+    8.648395082114646e-11
+   -2.818433537692151e-13
+   -8.145508875467845e-13
+   -2.162272824444328e-11
+    8.486453668018574e-11
+ 2.5e+09     
+    8.469544552641473e-11
+   -2.155926024625489e-11
+    8.648484424135681e-11
+   -8.149639475886933e-13
+   -1.022825015035805e-11
+    8.644955654702486e-11
+   -2.798141554250774e-13
+   -8.123171968003414e-13
+   -2.161233125605763e-11
+    8.483126301064557e-11
+ 2.6e+09     
+    8.466381644601125e-11
+   -2.154909115093917e-11
+    8.645198862721802e-11
+   -8.127077236829148e-13
+    -1.02226845630933e-11
+    8.641673308271596e-11
+   -2.777106605521883e-13
+   -8.100430125920139e-13
+   -2.160218589088073e-11
+    8.479957798313685e-11
+ 2.7e+09     
+    8.463366052126717e-11
+    -2.15391762840394e-11
+    8.642060559808845e-11
+   -8.104190025655238e-13
+    -1.02171990138627e-11
+    8.638537446969617e-11
+   -2.755469025482309e-13
+   -8.077365301650289e-13
+   -2.159228704597431e-11
+    8.476936649290474e-11
+ 2.8e+09     
+    8.460487316401111e-11
+   -2.152950873354381e-11
+    8.639059683556333e-11
+   -8.081056094842732e-13
+   -1.021179472380827e-11
+    8.635538456680167e-11
+   -2.733370992776192e-13
+   -8.054053449130229e-13
+   -2.158262894987158e-11
+    8.474052422541462e-11
+ 2.9e+09     
+    8.457735948033087e-11
+   -2.152008116232012e-11
+    8.636187294334369e-11
+   -8.057748019709965e-13
+   -1.020647265652601e-11
+     8.63266759455411e-11
+   -2.710951845760588e-13
+   -8.030565065997723e-13
+   -2.157320540386384e-11
+    8.471295657904957e-11
+ 3e+09       
+    8.455103327046927e-11
+   -2.151088602049314e-11
+    8.633435245099362e-11
+   -8.034333198711488e-13
+   -1.020123355316101e-11
+    8.629916885468163e-11
+   -2.688344581780033e-13
+   -8.006965730312998e-13
+   -2.156400995502222e-11
+    8.468657764642248e-11
+ 3.1e+09     
+    8.452581609877522e-11
+   -2.150191569417122e-11
+    8.630796089003389e-11
+   -8.010874324237145e-13
+   -1.019607795272979e-11
+     8.62727902700514e-11
+   -2.665673425517244e-13
+   -7.983316589316203e-13
+   -2.155503601749539e-11
+    8.466130927077385e-11
+ 3.2e+09     
+    8.450163644187394e-11
+   -2.149316260659788e-11
+    8.628262995126825e-11
+   -7.987429800469735e-13
+   -1.019100620317453e-11
+    8.624747303684047e-11
+   -2.643052313346325e-13
+   -7.959674781723875e-13
+   -2.154627695525002e-11
+    8.463708018442248e-11
+ 3.3e+09     
+    8.447842891705596e-11
+   -2.148461928430086e-11
+    8.625829672646163e-11
+   -7.964054101460191e-13
+   -1.018601846713525e-11
+    8.622315510644432e-11
+    -2.62058412653256e-13
+   -7.936093790357521e-13
+    -2.15377261367339e-11
+    8.461382523039105e-11
+ 3.4e+09     
+    8.445613358916547e-11
+    -2.14762783980611e-11
+    8.623490303400188e-11
+   -7.940798072350813e-13
+   -1.018111472533316e-11
+    8.619977886672585e-11
+   -2.598360509207031e-13
+   -7.912623730692711e-13
+   -2.152937696977011e-11
+     8.45914846648382e-11
+ 3.5e+09     
+    8.443469535212682e-11
+   -2.146813278635385e-11
+    8.621239482611061e-11
+   -7.917709181619837e-13
+   -1.017629477966074e-11
+    8.617729056262524e-11
+   -2.576462121186179e-13
+   -7.889311585165066e-13
+   -2.152122292322203e-11
+    8.457000353595709e-11
+ 3.6e+09     
+    8.441406338012013e-11
+    -2.14601754671865e-11
+    8.619072167394003e-11
+   -7.894831733985057e-13
+   -1.017155825747182e-11
+    8.615563980277311e-11
+   -2.554959195874523e-13
+   -7.866201394353077e-13
+   -2.151325754050858e-11
+    8.454933113399714e-11
+ 3.7e+09     
+    8.439419064292567e-11
+   -2.145239964287149e-11
+    8.616983632613354e-11
+   -7.872207053443567e-13
+   -1.016690461809005e-11
+    8.613477914683179e-11
+   -2.533912295914022e-13
+   -7.843334415681662e-13
+   -2.150547444882548e-11
+    8.452942050665697e-11
+ 3.8e+09     
+    8.437503347986106e-11
+   -2.144479870114826e-11
+    8.614969433591869e-11
+   -7.849873644728483e-13
+   -1.016233316216368e-11
+    8.611466376751828e-11
+    -2.51337318134055e-13
+   -7.820749258899394e-13
+   -2.149786736689667e-11
+    8.451022803405527e-11
+ 3.9e+09     
+    8.435655122686775e-11
+   -2.143736621514661e-11
+    8.613025375140305e-11
+    -7.82786733984476e-13
+   -1.015784304415938e-11
+    8.609525118058328e-11
+   -2.493385725195812e-13
+   -7.798482005849238e-13
+   -2.149043011320723e-11
+    8.449171305766026e-11
+ 4e+09       
+    8.433870589156748e-11
+   -2.143009594392589e-11
+     8.61114748634013e-11
+   -7.806221434670719e-13
+   -1.015343328799773e-11
+    8.607650103539997e-11
+    -2.47398682900874e-13
+   -7.776566320310042e-13
+   -2.148315661592909e-11
+    8.447383755783639e-11
+ 4.1e+09     
+    8.432146187143489e-11
+   -2.142298183469636e-11
+    8.609332000480569e-11
+   -7.784966819103422e-13
+   -1.014910280558052e-11
+    8.605837495830268e-11
+    -2.45520730502943e-13
+   -7.755033552126505e-13
+      -2.147604092514e-11
+    8.445656587501476e-11
+ 4.2e+09     
+    8.430478571057856e-11
+   -2.141601802731342e-11
+     8.60757533952441e-11
+   -7.764132102969519e-13
+   -1.014485041775041e-11
+    8.604083644044178e-11
+   -2.437072703649662e-13
+    -7.73391283854016e-13
+   -2.146907722743704e-11
+    8.443986446983741e-11
+ 4.3e+09     
+    8.428864589096329e-11
+   -2.140919886121668e-11
+    8.605874102456371e-11
+    -7.74374373896268e-13
+    -1.01406748770579e-11
+    8.602385076174913e-11
+   -2.419604073351662e-13
+   -7.713231204597066e-13
+   -2.146225986266543e-11
+     8.44237017179865e-11
+ 4.4e+09     
+     8.42730126542312e-11
+   -2.140251888465685e-11
+    8.604225056858163e-11
+   -7.723826143171495e-13
+   -1.013657489159742e-11
+    8.600738494267513e-11
+   -2.402818647167293e-13
+   -7.693013663716024e-13
+   -2.145558334220686e-11
+    8.440804773572994e-11
+ 4.5e+09     
+    8.425785785057873e-11
+   -2.139597286580536e-11
+    8.602625133057427e-11
+   -7.704401813303984e-13
+   -1.013254914911306e-11
+    8.599140771569092e-11
+   -2.386730454394484e-13
+   -7.673283318915071e-13
+   -2.144904236810262e-11
+     8.43928742325359e-11
+ 4.6e+09     
+    8.424315481142242e-11
+   -2.138955580517204e-11
+    8.601071420216931e-11
+   -7.685491444440235e-13
+   -1.012859634056859e-11
+    8.597588950913915e-11
+   -2.371350859589206e-13
+   -7.654061464769406e-13
+   -2.144263185220659e-11
+      8.4378154387387e-11
+ 4.7e+09     
+    8.422887824282912e-11
+   -2.138326294865444e-11
+    8.599561163766192e-11
+   -7.667114042010299e-13
+   -1.012471518242088e-11
+    8.596080243685022e-11
+   -2.356689032963334e-13
+   -7.635367689878079e-13
+   -2.143634693456939e-11
+    8.436386274569466e-11
+ 4.8e+09     
+    8.421500413692404e-11
+   -2.137708980050806e-11
+    8.598091763629867e-11
+   -7.649287031656113e-13
+   -1.012090443692383e-11
+    8.594612028795083e-11
+    -2.34275235755978e-13
+   -7.617219979413434e-13
+   -2.143018300032212e-11
+     8.43499751339541e-11
+ 4.9e+09     
+    8.420150969868607e-11
+   -2.137103213554147e-11
+    8.596660772773753e-11
+   -7.632026365656392e-13
+   -1.011716292991368e-11
+    8.593181851243672e-11
+   -2.329546779180722e-13
+   -7.599634817197171e-13
+   -2.142413569444687e-11
+    8.433646858950662e-11
+ 5e+09       
+    8.418837328574521e-11
+   -2.136508600990379e-11
+    8.595265895666632e-11
+   -7.615346625647205e-13
+   -1.011348956567193e-11
+    8.591787419925991e-11
+   -2.317077105201336e-13
+   -7.582627286671518e-13
+   -2.141820093396695e-11
+    8.432332130298796e-11
+ 5.1e+09     
+    8.417557435897482e-11
+   -2.135924776992559e-11
+    8.593904986341069e-11
+   -7.599261121434493e-13
+   -1.010988333861949e-11
+    8.590426604485554e-11
+   -2.305347258253831e-13
+   -7.566211170105156e-13
+   -2.141237491725096e-11
+    8.431051257123621e-11
+ 5.2e+09     
+    8.416309344184839e-11
+   -2.135351405858887e-11
+    8.592576045822616e-11
+   -7.583781985757933e-13
+   -1.010634334175102e-11
+    8.589097431110384e-11
+   -2.294360490428125e-13
+   -7.550399045377402e-13
+   -2.140665413028137e-11
+    8.429802275862758e-11
+ 5.3e+09     
+    8.415091208670833e-11
+   -2.134788181932833e-11
+    8.591277218781569e-11
+   -7.568920264918554e-13
+   -1.010286877186333e-11
+    8.587798077266489e-11
+   -2.284119563185384e-13
+   -7.535202379719959e-13
+   -2.140103534988079e-11
+    8.428583326498647e-11
+ 5.4e+09     
+    8.413901284625933e-11
+   -2.134234829699103e-11
+    8.590006789339703e-11
+   -7.554686005224338e-13
+   -1.009945893175735e-11
+    8.586526865439258e-11
+    -2.27462689767796e-13
+   -7.520631619854356e-13
+   -2.139551564401001e-11
+    8.427392649840014e-11
+ 5.5e+09     
+    8.412737924877433e-11
+   -2.133691103589906e-11
+    8.588763176032265e-11
+   -7.541088335238611e-13
+   -1.009611322969248e-11
+    8.585282256010828e-11
+   -2.265884699656436e-13
+   -7.506696278041748e-13
+   -2.139009236934396e-11
+    8.426228585144449e-11
+ 5.6e+09     
+    8.411599577567321e-11
+   -2.133156787506537e-11
+    8.587544925982168e-11
+    -7.52813554383581e-13
+   -1.009283117644638e-11
+    8.584062839440473e-11
+   -2.257895062645671e-13
+    -7.49340501365076e-13
+   -2.138476316639601e-11
+     8.42508956795062e-11
+ 5.7e+09     
+    8.410484784030596e-11
+   -2.132631694069841e-11
+    8.586350708386463e-11
+   -7.515835154084678e-13
+   -1.008961238037773e-11
+    8.582867327936317e-11
+   -2.250660052606047e-13
+    -7.48076570994899e-13
+    -2.13795259524978e-11
+    8.423974128006196e-11
+ 5.8e+09     
+    8.409392176694898e-11
+   -2.132115663620051e-11
+    8.585179307444628e-11
+     -7.5041939929886e-13
+   -1.008645654090844e-11
+    8.581694546812059e-11
+   -2.244181776870468e-13
+   -7.468785545924247e-13
+   -2.137437891295444e-11
+    8.422880887195559e-11
+ 5.9e+09     
+    8.408320476919299e-11
+   -2.131608562991238e-11
+    8.584029614875631e-11
+   -7.493218257124259e-13
+   -1.008336344083868e-11
+    8.580543425716024e-11
+     -2.2384624397681e-13
+   -7.457471063040421e-13
+   -2.136932049068909e-11
+     8.42180855738867e-11
+ 6e+09       
+    8.407268492707682e-11
+   -2.131110284088986e-11
+    8.582900622176503e-11
+   -7.482913574229126e-13
+   -1.008033293788576e-11
+    8.579412989903737e-11
+   -2.233504387010526e-13
+   -7.446828226926732e-13
+   -2.136434937466988e-11
+    8.420755938149879e-11
+ 6.1e+09     
+     8.40623511624826e-11
+   -2.130620742301402e-11
+    8.581791412771849e-11
+   -7.473285060802301e-13
+   -1.007736495580204e-11
+    8.578302351702846e-11
+   -2.229310140623906e-13
+   -7.436862484082694e-13
+    -2.13594644873825e-11
+    8.419721914261903e-11
+ 6.2e+09     
+    8.405219321246896e-11
+   -2.130139874774063e-11
+    8.580701154193248e-11
+   -7.464337375795767e-13
+   -1.007445947538234e-11
+    8.577210702293411e-11
+   -2.225882425958656e-13
+   -7.427578813755676e-13
+   -2.135466497157566e-11
+    8.418705453036045e-11
+ 6.3e+09     
+    8.404220160036787e-11
+   -2.129667638579034e-11
+    8.579629090411562e-11
+   -7.456074770490609e-13
+   -1.007161652562077e-11
+    8.576137303899766e-11
+   -2.223224192090005e-13
+   -7.418981775207357e-13
+   -2.134995017647154e-11
+    8.417705601394396e-11
+ 6.4e+09     
+    8.403236760460251e-11
+   -2.129204008806826e-11
+    8.578574534426738e-11
+     -7.4485011346683e-13
+   -1.006883617522634e-11
+    8.575081482463417e-11
+     -2.2213386267375e-13
+   -7.411075550636941e-13
+   -2.134531964359473e-11
+    8.416721482722659e-11
+ 6.5e+09     
+    8.402268322530843e-11
+   -2.128748976608587e-11
+     8.57753686119911e-11
+   -7.441620039203154e-13
+   -1.006611852465613e-11
+    8.574042620842516e-11
+   -2.220229166670945e-13
+    -7.40386398406094e-13
+   -2.134077309234401e-11
+    8.415752293504203e-11
+ 6.6e+09     
+    8.401314114893963e-11
+   -2.128302547213967e-11
+    8.576515500986192e-11
+   -7.435434775216716e-13
+   -1.006346369877915e-11
+    8.573020152561304e-11
+   -2.219899504433974e-13
+   -7.397350616478736e-13
+   -2.133631040539766e-11
+    8.414797299755056e-11
+ 6.7e+09     
+    8.400373471112787e-11
+   -2.127864737947945e-11
+    8.575509933129613e-11
+   -7.429948389948097e-13
+    -1.00608718402425e-11
+    8.572013556115284e-11
+   -2.220353592098563e-13
+   -7.391538717661744e-13
+    -2.13319316140234e-11
+    8.413855833287985e-11
+ 6.8e+09     
+    8.399445785812799e-11
+   -2.127435576268067e-11
+    8.574519680319583e-11
+   -7.425163719503602e-13
+    -1.00583431035767e-11
+    8.571022349822413e-11
+   -2.221595642662112e-13
+   -7.386431314911764e-13
+   -2.132763688334015e-11
+    8.412927287838882e-11
+ 6.9e+09     
+    8.398530510722924e-11
+   -2.127015097841306e-11
+    8.573544303348888e-11
+   -7.421083418655361e-13
+   -1.005587765004689e-11
+    8.570046087199357e-11
+   -2.223630129611688e-13
+   -7.382031219127898e-13
+   -2.132342649756506e-11
+    8.412011115093204e-11
+ 7e+09       
+    8.397627150654172e-11
+   -2.126603344678013e-11
+    8.572583396355808e-11
+   -7.417709987863846e-13
+   -1.005347564323468e-11
+    8.569084352833635e-11
+   -2.226461785102806e-13
+   -7.378341048510068e-13
+   -2.131930084526827e-11
+    8.411106820651695e-11
+ 7.1e+09     
+    8.396735259457504e-11
+   -2.126200363338271e-11
+    8.571636582545317e-11
+   -7.415045797698021e-13
+   -1.005113724531661e-11
+    8.568136758716161e-11
+   -2.230095597134315e-13
+   -7.375363250211335e-13
+   -2.131526040464826e-11
+    8.410213959975539e-11
+ 7.2e+09     
+    8.395854436002553e-11
+   -2.125806203224329e-11
+    8.570703510369437e-11
+   -7.413093110825391e-13
+   -1.004886261399332e-11
+    8.567202940996029e-11
+   -2.234536806042132e-13
+   -7.373100120228306e-13
+    -2.13113057288376e-11
+     8.40933213434952e-11
+ 7.3e+09     
+    8.394984320216824e-11
+   -2.125420914970818e-11
+    8.569783850142597e-11
+   -7.411854101739964e-13
+   -1.004665190001514e-11
+    8.566282557117375e-11
+   -2.239790900584065e-13
+   -7.371553821795199e-13
+   -2.130743743124667e-11
+     8.40846098690025e-11
+ 7.4e+09     
+     8.39412458922216e-11
+   -2.125044548942691e-11
+    8.568877291063337e-11
+   -7.411330874389378e-13
+   -1.004450524524473e-11
+    8.565375283298662e-11
+   -2.245863613842014e-13
+     -7.3707264025188e-13
+   -2.130365617095342e-11
+    8.407600198702675e-11
+ 7.5e+09     
+    8.393274953601622e-11
+   -2.124677153849112e-11
+    8.567983538611721e-11
+   -7.411525477855103e-13
+   -1.004242278119625e-11
+     8.56448081231569e-11
+   -2.252760919129248e-13
+   -7.370619810462253e-13
+   -2.129996263815092e-11
+    8.406749485004858e-11
+ 7.6e+09     
+    8.392435153825634e-11
+   -2.124318775479761e-11
+    8.567102312290793e-11
+   -7.412439920230074e-13
+   -1.004040462799055e-11
+    8.563598851551821e-11
+   -2.260489026055082e-13
+   -7.371235909356736e-13
+   -2.129635753966918e-11
+    8.405908591596542e-11
+ 7.7e+09     
+    8.391604956861103e-11
+   -2.123969455568156e-11
+    8.566233343680224e-11
+   -7.414076180831209e-13
+   -1.003845089366862e-11
+    8.562729121281944e-11
+   -2.269054376868761e-13
+   -7.372576493088428e-13
+   -2.129284158459478e-11
+     8.40507729134262e-11
+ 7.8e+09     
+    8.390784152983017e-11
+   -2.123629230785105e-11
+    8.565376374771119e-11
+   -7.416436220873536e-13
+   -1.003656167380811e-11
+    8.561871353159174e-11
+   -2.278463643177892e-13
+   -7.374643299578137e-13
+    -2.12894154700203e-11
+    8.404255380898353e-11
+ 7.9e+09     
+    8.389972552802579e-11
+   -2.123298131863673e-11
+    8.564531156552494e-11
+   -7.419521992724809e-13
+   -1.003473705139326e-11
+    8.561025288877238e-11
+   -2.288723723113125e-13
+   -7.377438024143158e-13
+    -2.12860798669653e-11
+    8.403442677618888e-11
+ 8e+09       
+    8.389169984521321e-11
+   -2.122976182855327e-11
+    8.563697447821271e-11
+   -7.423335447852107e-13
+    -1.00329770968917e-11
+    8.560190678984352e-11
+   -2.299841738991009e-13
+   -7.380962332399721e-13
+   -2.128283540652059e-11
+    8.402639016671508e-11
+ 8.1e+09     
+    8.388376291416522e-11
+   -2.122663400515669e-11
+    8.562875014189735e-11
+   -7.427878543563552e-13
+   -1.003128186849778e-11
+    8.559367281827861e-11
+   -2.311825035509155e-13
+   -7.385217872741298e-13
+   -2.127968266627984e-11
+    8.401844248355927e-11
+ 8.2e+09     
+    8.387591329558746e-11
+   -2.122359793816547e-11
+    8.562063627266536e-11
+   -7.433153248642334e-13
+   -1.002965141250599e-11
+    8.558554862612046e-11
+   -2.324681178493491e-13
+   -7.390206288400696e-13
+   -2.127662215713253e-11
+    8.401058235634248e-11
+ 8.3e+09     
+     8.38681496575913e-11
+   -2.122065363580148e-11
+    8.561263063989062e-11
+   -7.439161547964369e-13
+   -1.002808576378305e-11
+    8.557753192554511e-11
+   -2.338417954204911e-13
+      -7.395929229082e-13
+   -2.127365431050391e-11
+    8.400280851869897e-11
+ 8.4e+09     
+    8.386047075740632e-11
+   -2.121780102229473e-11
+    8.560473106087371e-11
+   -7.445905446185727e-13
+   -1.002658494631175e-11
+    8.556962048129049e-11
+    -2.35304336920187e-13
+   -7.402388362129709e-13
+   -2.127077946613733e-11
+     8.39951197877263e-11
+ 8.5e+09     
+    8.385287542525068e-11
+   -2.121503993648692e-11
+    8.559693539661633e-11
+   -7.453386970580495e-13
+   -1.002514897378334e-11
+    8.556181210385505e-11
+   -2.368565650748115e-13
+   -7.409585383184265e-13
+    -2.12679978605232e-11
+    8.398751504544716e-11
+ 8.6e+09     
+    8.384536255025525e-11
+    -2.12123701314583e-11
+    8.558924154856856e-11
+   -7.461608173108354e-13
+   -1.002377785021919e-11
+    8.555410464339359e-11
+   -2.384993247747142e-13
+   -7.417522026260178e-13
+    -2.12653096160849e-11
+    8.397999322222135e-11
+ 8.7e+09     
+    8.383793106832136e-11
+   -2.120979127509761e-11
+    8.558164745620332e-11
+   -7.470571131783366e-13
+   -1.002247157060567e-11
+    8.554649598425299e-11
+   -2.402334832181024e-13
+   -7.426200073170995e-13
+   -2.126271473123716e-11
+    8.397255328203753e-11
+ 8.8e+09     
+    8.383057995178054e-11
+   -2.120730295152841e-11
+    8.557415109529152e-11
+   -7.480277951416653e-13
+   -1.002123012152925e-11
+    8.553898404011008e-11
+   -2.420599301027281e-13
+   -7.435621362221016e-13
+   -2.126021307143334e-11
+    8.396519420960458e-11
+ 8.9e+09     
+    8.382330820071646e-11
+   -2.120490466330204e-11
+    8.556675047676017e-11
+   -7.490730763798769e-13
+   -1.002005348180096e-11
+    8.553156674968231e-11
+   -2.439795778625711e-13
+   -7.445787796077783e-13
+   -2.125780436131626e-11
+    8.395791499915929e-11
+ 9e+09       
+    8.381611483580541e-11
+   -2.120259583426511e-11
+    8.555944364603437e-11
+   -7.501931727386697e-13
+   -1.001894162306234e-11
+    8.552424207299517e-11
+   -2.459933619466614e-13
+   -7.456701348741088e-13
+   -2.125548817808263e-11
+    8.395071464490432e-11
+ 9.1e+09     
+    8.380899889253005e-11
+   -2.120037581300966e-11
+    8.555222868277174e-11
+   -7.513883026557049e-13
+   -1.001789451036601e-11
+    8.551700798819543e-11
+   -2.481022411371248e-13
+   -7.468364071527385e-13
+   -2.125326394616202e-11
+    8.394359213298677e-11
+ 9.2e+09     
+    8.380195941662367e-11
+   -2.119824387681457e-11
+    8.554510370091214e-11
+   -7.526586870482263e-13
+   -1.001691210272639e-11
+    8.550986248890329e-11
+   -2.503071979038438e-13
+   -7.480778097997116e-13
+   -2.125113093329935e-11
+    8.393654643493151e-11
+ 9.3e+09     
+    8.379499546060686e-11
+   -2.119619923598937e-11
+    8.553806684897224e-11
+   -7.540045491687278e-13
+   -1.001599435363713e-11
+    8.550280358210017e-11
+    -2.52609238793172e-13
+   -7.493945647760895e-13
+   -2.124908824811377e-11
+    8.392957650243606e-11
+ 9.4e+09     
+    8.378810608128073e-11
+   -2.119424103853467e-11
+    8.553111631052644e-11
+   -7.554261144336153e-13
+   -1.001514121155295e-11
+    8.549582928654761e-11
+   -2.550093948485825e-13
+   -7.507869029116318e-13
+   -2.124713483918859e-11
+    8.392268126344279e-11
+ 9.5e+09     
+    8.378129033805217e-11
+    -2.11923683750381e-11
+    8.552425030482058e-11
+   -7.569236102299112e-13
+   -1.001435262033466e-11
+    8.548893763173071e-11
+   -2.575087220614173e-13
+   -7.522550640481005e-13
+   -2.124526949572505e-11
+    8.391585961939552e-11
+ 9.6e+09     
+    8.377454729197218e-11
+   -2.119058028372963e-11
+    8.551746708747346e-11
+    -7.58497265704469e-13
+   -1.001362851965699e-11
+    8.548212665731833e-11
+   -2.601083018503905e-13
+   -7.537992970606519e-13
+   -2.124349084976947e-11
+    8.390911044359488e-11
+ 9.7e+09     
+    8.376787600537767e-11
+   -2.118887575562587e-11
+    8.551076495122924e-11
+   -7.601473115399243e-13
+   -1.001296884537947e-11
+    8.547539441312477e-11
+    -2.62809241568875e-13
+   -7.554198597576709e-13
+   -2.124179737999783e-11
+    8.390243258056145e-11
+ 9.8e+09     
+    8.376127554203544e-11
+   -2.118725373969873e-11
+    8.550414222672634e-11
+   -7.618739797212503e-13
+   -1.001237352988081e-11
+    8.546873895955275e-11
+   -2.656126750395663e-13
+   -7.571170186613149e-13
+   -2.124018741701632e-11
+    8.389582484631768e-11
+ 9.9e+09     
+    8.375474496769834e-11
+   -2.118571314801147e-11
+    8.549759728325697e-11
+   -7.636775032964617e-13
+   -1.001184250235861e-11
+    8.546215836849665e-11
+   -2.685197631165044e-13
+   -7.588910486731447e-13
+   -2.123865915011114e-11
+    8.388928602949918e-11
+ 1e+10       
+    8.374828335098979e-11
+   -2.118425286076998e-11
+    8.549112852949293e-11
+   -7.655581161346286e-13
+   -1.001137568909523e-11
+     8.54556507246693e-11
+   -2.715316942750253e-13
+   -7.607422326310141e-13
+   -2.123721063535514e-11
+     8.38828148932047e-11
+ 1.01e+10    
+    8.374176925262979e-11
+   -2.118332705501576e-11
+    8.548486851426227e-11
+   -7.677697184886483e-13
+   -1.001128520682366e-11
+    8.544940020698455e-11
+   -2.746968601270755e-13
+   -7.629297733125297e-13
+   -2.123627897437604e-11
+    8.387628224572417e-11
+ 1.02e+10    
+    8.373529664749316e-11
+   -2.118241937361016e-11
+     8.54786657769058e-11
+    -7.70002818028213e-13
+   -1.001120430458993e-11
+    8.544320535121991e-11
+    -2.77894753098657e-13
+   -7.651389592183628e-13
+   -2.123536484949096e-11
+    8.386979108034153e-11
+ 1.03e+10    
+    8.372886577944913e-11
+   -2.118152993838519e-11
+    8.547252060195258e-11
+   -7.722572009643641e-13
+   -1.001113294492601e-11
+    8.543706647218625e-11
+   -2.811248330920193e-13
+   -7.673695777968157e-13
+   -2.123446839051573e-11
+    8.386334163938702e-11
+ 1.04e+10    
+    8.372247685659804e-11
+   -2.118065886216766e-11
+    8.546643323807506e-11
+    -7.74532650971598e-13
+   -1.001107109020586e-11
+    8.543098384906882e-11
+   -2.843865530937285e-13
+     -7.6962141381145e-13
+   -2.123358971833501e-11
+    8.385693412928849e-11
+ 1.05e+10    
+    8.371613005272023e-11
+   -2.117980624909924e-11
+    8.546040389960065e-11
+   -7.768289493928517e-13
+   -1.001101870283026e-11
+    8.542495772690379e-11
+   -2.876793596957041e-13
+   -7.718942495497908e-13
+   -2.123272894520951e-11
+     8.38505687220194e-11
+ 1.06e+10    
+    8.370982550869987e-11
+   -2.117897219495289e-11
+    8.545443276798855e-11
+   -7.791458754403795e-13
+   -1.001097574540034e-11
+    8.541898831801917e-11
+   -2.910026936058017e-13
+   -7.741878650279736e-13
+   -2.123188617508038e-11
+    8.384424555652262e-11
+ 1.07e+10    
+    8.370356333392497e-11
+   -2.117815678744548e-11
+    8.544851999326477e-11
+   -7.814832063926976e-13
+   -1.001094218087942e-11
+    8.541307580343862e-11
+   -2.943559901475637e-13
+   -7.765020381913339e-13
+   -2.123106150387046e-11
+    8.383796474011036e-11
+ 1.08e+10    
+    8.369734360766209e-11
+   -2.117736010654639e-11
+    8.544266569541997e-11
+   -7.838407177870963e-13
+   -1.001091797274363e-11
+     8.54072203342473e-11
+   -2.977386797489394e-13
+   -7.788365451106773e-13
+   -2.123025501978168e-11
+     8.38317263498388e-11
+ 1.09e+10    
+    8.369116638040468e-11
+   -2.117658222478165e-11
+    8.543686996576622e-11
+     -7.8621818360779e-13
+   -1.001090308512173e-11
+    8.540142203292125e-11
+   -3.011501884196563e-13
+   -7.811911601740746e-13
+   -2.122946680358903e-11
+    8.382553043385579e-11
+ 1.1e+10     
+    8.368503167519434e-11
+   -2.117582320753333e-11
+    8.543113286825462e-11
+   -7.886153764695289e-13
+   -1.001089748292425e-11
+    8.539568099461621e-11
+    -3.04589938217147e-13
+   -7.835656562740318e-13
+   -2.122869692893005e-11
+    8.381937701272238e-11
+ 1.11e+10    
+    8.367893948891409e-11
+   -2.117508311333432e-11
+    8.542545444075303e-11
+   -7.910320677963565e-13
+   -1.001090113196249e-11
+    8.538999728842015e-11
+   -3.080573477007608e-13
+   -7.859598049899736e-13
+   -2.122794546259005e-11
+    8.381326608070552e-11
+ 1.12e+10    
+    8.367288979355412e-11
+   -2.117436199415748e-11
+    8.541983469628288e-11
+   -7.934680279958252e-13
+   -1.001091399905729e-11
+     8.53843709585657e-11
+   -3.115518323741772e-13
+   -7.883733767659233e-13
+   -2.122721246478268e-11
+    8.380719760704292e-11
+ 1.13e+10    
+    8.366688253744692e-11
+   -2.117365989569998e-11
+    8.541427362421648e-11
+   -7.959230266280791e-13
+    -1.00109360521384e-11
+    8.537880202560398e-11
+   -3.150728051159303e-13
+   -7.908061410832167e-13
+   -2.122649798942546e-11
+    8.380117153717937e-11
+ 1.14e+10    
+    8.366091764647488e-11
+   -2.117297685766175e-11
+    8.540877119143504e-11
+    -7.98396832570198e-13
+   -1.001096726033439e-11
+    8.537329048754048e-11
+   -3.186196765979011e-13
+   -7.932578666283056e-13
+   -2.122580208441043e-11
+    8.379518779397243e-11
+ 1.15e+10    
+    8.365499502524686e-11
+   -2.117231291401836e-11
+     8.54033273434457e-11
+   -8.008892141753669e-13
+   -1.001100759405366e-11
+    8.536783632093206e-11
+     -3.2219185569181e-13
+   -7.957283214554696e-13
+   -2.122512479186938e-11
+    8.378924627886987e-11
+ 1.16e+10    
+    8.364911455824475e-11
+   -2.117166809328807e-11
+    8.539794200546076e-11
+   -8.033999394271406e-13
+   -1.001105702505665e-11
+    8.536243948194499e-11
+   -3.257887498635926e-13
+   -7.982172731445057e-13
+   -2.122446614843359e-11
+    8.378334687305586e-11
+ 1.17e+10    
+    8.364327611094051e-11
+   -2.117104241879289e-11
+    8.539261508343727e-11
+   -8.059287760884622e-13
+      -1.001111552652e-11
+    8.535709990737632e-11
+   -3.294097655557461e-13
+   -8.007244889532095e-13
+   -2.122382618548812e-11
+    8.377748943856755e-11
+ 1.18e+10    
+    8.363747953088185e-11
+   -2.117043590891351e-11
+    8.538734646507741e-11
+     -8.0847549184577e-13
+   -1.001118307309229e-11
+    8.535181751563658e-11
+   -3.330543085575726e-13
+    -8.03249735964848e-13
+   -2.122320492942028e-11
+     8.37716738193814e-11
+ 1.19e+10    
+     8.36317246487474e-11
+   -2.116984857733808e-11
+    8.538213602079279e-11
+   -8.110398544478248e-13
+   -1.001125964094264e-11
+     8.53465922076956e-11
+   -3.367217843634261e-13
+   -8.057927812303779e-13
+   -2.122260240186203e-11
+    8.376589984246764e-11
+ 1.2e+10     
+    8.362601127937182e-11
+   -2.116928043330472e-11
+    8.537698360462949e-11
+   -8.136216318394963e-13
+    -1.00113452078015e-11
+    8.534142386799184e-11
+   -3.404115985189925e-13
+   -8.083533919056063e-13
+   -2.122201861992693e-11
+    8.376016731881632e-11
+ 1.21e+10    
+    8.362033922273925e-11
+   -2.116873148183759e-11
+    8.537188905515765e-11
+   -8.162205922905108e-13
+   -1.001143975299488e-11
+    8.533631236530567e-11
+   -3.441231569556682e-13
+   -8.109313353831646e-13
+   -2.122145359644052e-11
+    8.375447604443077e-11
+ 1.22e+10    
+    8.361470826494653e-11
+    -2.11682017239766e-11
+    8.536685219632377e-11
+   -8.188365045189619e-13
+   -1.001154325747153e-11
+    8.533125755359645e-11
+   -3.478558663131449e-13
+   -8.135263794193864e-13
+   -2.122090734016473e-11
+    8.374882580129088e-11
+ 1.23e+10    
+    8.360911817913584e-11
+   -2.116769115700074e-11
+    8.536187283826917e-11
+   -8.214691378099626e-13
+   -1.001165570382406e-11
+    8.532625927280566e-11
+   -3.516091342502892e-13
+   -8.161382922561558e-13
+   -2.122037985601633e-11
+    8.374321635828725e-11
+ 1.24e+10    
+    8.360356872639647e-11
+   -2.116719977464468e-11
+    8.535695077811204e-11
+   -8.241182621291779e-13
+   -1.001177707630385e-11
+    8.532131734962491e-11
+   -3.553823697444463e-13
+   -8.187668427376402e-13
+   -2.121987114527892e-11
+    8.373764747212306e-11
+ 1.25e+10    
+    8.359805965663631e-11
+   -2.116672756730909e-11
+    8.535208580069649e-11
+   -8.267836482313694e-13
+   -1.001190736083033e-11
+    8.531643159823091e-11
+    -3.59174983379303e-13
+   -8.214118004220918e-13
+   -2.121938120580841e-11
+    8.373211888818663e-11
+ 1.26e+10    
+    8.359259070942308e-11
+   -2.116627452226423e-11
+     8.53472776793089e-11
+   -8.294650677641457e-13
+   -1.001204654499493e-11
+    8.531160182098847e-11
+   -3.629863876214255e-13
+   -8.240729356886572e-13
+   -2.121891003223301e-11
+    8.372663034139423e-11
+ 1.27e+10    
+    8.358716161479562e-11
+   -2.116584062384713e-11
+    8.534252617636073e-11
+   -8.321622933667213e-13
+   -1.001219461805971e-11
+    8.530682780911952e-11
+   -3.668159970856652e-13
+   -8.267500198393398e-13
+   -2.121845761614576e-11
+    8.372118155700189e-11
+ 1.28e+10    
+    8.358177209404479e-11
+   -2.116542585365208e-11
+    8.533783104404091e-11
+   -8.348750987640635e-13
+   -1.001235157095136e-11
+    8.530210934334303e-11
+   -3.706632287895316e-13
+   -8.294428251961498e-13
+    -2.12180239462918e-11
+    8.371577225138904e-11
+ 1.29e+10    
+     8.35764218604658e-11
+   -2.116503019071481e-11
+    8.533319202493719e-11
+   -8.376032588561212e-13
+   -1.001251739625069e-11
+    8.529744619448369e-11
+   -3.745275023968204e-13
+   -8.321511251934376e-13
+   -2.121760900874871e-11
+    8.371040213281147e-11
+ 1.3e+10     
+    8.357111062007999e-11
+   -2.116465361168997e-11
+    8.532860885262793e-11
+   -8.403465498025811e-13
+   -1.001269208817775e-11
+    8.529283812405108e-11
+      -3.784082404505e-13
+    -8.34874694465652e-13
+   -2.121721278710082e-11
+    8.370507090212625e-11
+ 1.31e+10    
+    8.356583807232856e-11
+   -2.116429609102209e-11
+    8.532408125224427e-11
+   -8.431047491029698e-13
+   -1.001287564257314e-11
+    8.528828488479031e-11
+   -3.823048685952156e-13
+   -8.376133089304193e-13
+   -2.121683526260694e-11
+    8.369977825348684e-11
+ 1.32e+10    
+    8.356060391073694e-11
+   -2.116395760111054e-11
+    8.531960894100613e-11
+   -8.458776356723291e-13
+   -1.001306805687564e-11
+    8.528378622120533e-11
+   -3.862168157894904e-13
+   -8.403667458671554e-13
+    -2.12164764143624e-11
+    8.369452387501077e-11
+ 1.33e+10    
+    8.355540782355143e-11
+   -2.116363811246744e-11
+    8.531519162872887e-11
+   -8.486649899124989e-13
+   -1.001326933009622e-11
+    8.527934187005456e-11
+    -3.90143514507849e-13
+   -8.431347839912814e-13
+   -2.121613621945426e-11
+    8.368930744941863e-11
+ 1.34e+10    
+    8.355024949434683e-11
+   -2.116333759386971e-11
+     8.53108290183051e-11
+   -8.514665937790364e-13
+    -1.00134794627892e-11
+    8.527495156082132e-11
+   -3.940844009330938e-13
+   -8.459172035239994e-13
+   -2.121581465311093e-11
+    8.368412865464531e-11
+ 1.35e+10    
+     8.35451286026074e-11
+   -2.116305601250491e-11
+    8.530652080616164e-11
+   -8.542822308440331e-13
+    -1.00136984570202e-11
+    8.527061501615894e-11
+   -3.980389151388841e-13
+   -8.487137862579655e-13
+   -2.121551168884531e-11
+    8.367898716442399e-11
+ 1.36e+10    
+    8.354004482427995e-11
+   -2.116279333411034e-11
+     8.53022666826904e-11
+   -8.571116863547647e-13
+   -1.001392631633172e-11
+     8.52663319523115e-11
+   -4.020065012628821e-13
+   -8.515243156186746e-13
+   -2.121522729859212e-11
+    8.367388264884315e-11
+ 1.37e+10    
+    8.353499783229999e-11
+   -2.116254952310657e-11
+    8.529806633265773e-11
+   -8.599547472883338e-13
+   -1.001416304570596e-11
+    8.526210207951157e-11
+   -4.059866076706037e-13
+   -8.543485767219747e-13
+   -2.121496145283911e-11
+    8.366881477487658e-11
+ 1.38e+10    
+    8.352998729709135e-11
+   -2.116232454272464e-11
+    8.529391943558964e-11
+   -8.628112024023894e-13
+   -1.001440865152572e-11
+    8.525792510235562e-11
+   -4.099786871102912e-13
+   -8.571863564274223e-13
+    -2.12147141207526e-11
+    8.366378320688798e-11
+ 1.39e+10    
+    8.352501288704034e-11
+   -2.116211835512734e-11
+     8.52898256661365e-11
+   -8.656808422821335e-13
+   -1.001466314153317e-11
+    8.525380072015763e-11
+   -4.139821968588836e-13
+   -8.600374433879594e-13
+   -2.121448527029703e-11
+    8.365878760710868e-11
+ 1.4e+10     
+    8.352007426894324e-11
+   -2.116193092152448e-11
+    8.528578469441578e-11
+   -8.685634593834486e-13
+   -1.001492652478685e-11
+    8.524972862728239e-11
+   -4.179965988594496e-13
+   -8.629016280957527e-13
+   -2.121427486834889e-11
+      8.3653827636091e-11
+ 1.41e+10    
+    8.351517110842874e-11
+   -2.116176220228258e-11
+    8.528179618633589e-11
+   -8.714588480725756e-13
+   -1.001519881161714e-11
+    8.524570851345874e-11
+   -4.220213598501717e-13
+   -8.657787029244389e-13
+   -2.121408288080487e-11
+    8.364890295313585e-11
+ 1.42e+10    
+    8.351030307035636e-11
+   -2.116161215702867e-11
+    8.527785980390047e-11
+   -8.743668046622569e-13
+   -1.001548001358036e-11
+    8.524174006407526e-11
+   -4.260559514851557e-13
+   -8.686684621677652e-13
+   -2.121390927268483e-11
+    8.364401321669632e-11
+ 1.43e+10    
+    8.350546981918961e-11
+   -2.116148074474864e-11
+    8.527397520549412e-11
+    -8.77287127444386e-13
+   -1.001577014341166e-11
+    8.523782296045572e-11
+   -4.300998504473041e-13
+     -8.7157070207486e-13
+   -2.121375400822888e-11
+    8.363915808475713e-11
+ 1.44e+10    
+     8.35006710193454e-11
+   -2.116136792387986e-11
+    8.527014204615156e-11
+   -8.802196167195355e-13
+   -1.001606921497693e-11
+    8.523395688011934e-11
+   -4.341525385533819e-13
+   -8.744852208821391e-13
+   -2.121361705098949e-11
+    8.363433721519016e-11
+ 1.45e+10    
+    8.349590633552026e-11
+   -2.116127365239872e-11
+    8.526635997780932e-11
+   -8.831640748231209e-13
+    -1.00163772432239e-11
+    8.523014149702448e-11
+   -4.382135028516008e-13
+   -8.774118188419546e-13
+   -2.121349836391825e-11
+    8.362955026608724e-11
+ 1.46e+10    
+    8.349117543299337e-11
+   -2.116119788790256e-11
+    8.526262864954212e-11
+   -8.861203061486412e-13
+    -1.00166942441325e-11
+     8.52263764817956e-11
+   -4.422822357118316e-13
+   -8.803502982481849e-13
+   -2.121339790944737e-11
+    8.362479689606999e-11
+ 1.47e+10    
+    8.348647797790722e-11
+   -2.116114058768663e-11
+    8.525894770778431e-11
+   -8.890881171678288e-13
+   -1.001702023466484e-11
+    8.522266150193715e-11
+    -4.46358234908719e-13
+   -8.833004634587062e-13
+   -2.121331564956645e-11
+    8.362007676457741e-11
+ 1.48e+10    
+    8.348181363752605e-11
+   -2.116110170881606e-11
+    8.525531679653702e-11
+   -8.920673164479485e-13
+   -1.001735523271483e-11
+    8.521899622203291e-11
+   -4.504410036979019e-13
+   -8.862621209150123e-13
+    -2.12132515458943e-11
+    8.361538953213211e-11
+ 1.49e+10    
+    8.347718208047293e-11
+   -2.116108120819258e-11
+    8.525173555756148e-11
+   -8.950577146663791e-13
+   -1.001769925705741e-11
+    8.521538030393188e-11
+   -4.545300508855042e-13
+   -8.892350791590115e-13
+   -2.121320555974563e-11
+    8.361073486058486e-11
+ 1.5e+10     
+    8.347258297694575e-11
+   -2.116107904261678e-11
+    8.524820363056014e-11
+   -8.980591246224388e-13
+   -1.001805232729808e-11
+    8.521181340692273e-11
+   -4.586248908911498e-13
+   -8.922191488470575e-13
+   -2.121317765219375e-11
+    8.360611241333859e-11
+ 1.51e+10    
+    8.346801599891318e-11
+   -2.116109516884555e-11
+    8.524472065334524e-11
+   -9.010713612467095e-13
+   -1.001841446382211e-11
+    8.520829518789559e-11
+   -4.627250438047015e-13
+   -8.952141427613815e-13
+    -2.12131677841281e-11
+    8.360152185555205e-11
+ 1.52e+10    
+    8.346348082028984e-11
+   -2.116112954364484e-11
+    8.524128626199705e-11
+   -9.040942416078464e-13
+   -1.001878568774426e-11
+    8.520482530149425e-11
+   -4.668300354368809e-13
+   -8.982198758190061e-13
+     -2.1213175916308e-11
+     8.35969628543242e-11
+ 1.53e+10    
+     8.34589771170924e-11
+   -2.116118212383816e-11
+    8.523790009100999e-11
+   -9.071275849170092e-13
+   -1.001916602085856e-11
+    8.520140340025607e-11
+   -4.709393973640096e-13
+   -9.012361650782506e-13
+   -2.121320200941137e-11
+    8.359243507885869e-11
+ 1.54e+10    
+    8.345450456757709e-11
+   -2.116125286635066e-11
+       8.523456177343e-11
+   -9.101712125300823e-13
+   -1.001955548558874e-11
+    8.519802913474558e-11
+   -4.750526669670521e-13
+   -9.042628297428636e-13
+   -2.121324602408015e-11
+    8.358793820060967e-11
+ 1.55e+10    
+    8.345006285235842e-11
+   -2.116134172824914e-11
+    8.523127094098179e-11
+   -9.132249479475961e-13
+   -1.001995410493899e-11
+    8.519470215367584e-11
+   -4.791693874651701e-13
+   -9.072996911639518e-13
+   -2.121330792096102e-11
+    8.358347189341016e-11
+ 1.56e+10    
+    8.344565165451062e-11
+   -2.116144866677793e-11
+    8.522802722418787e-11
+   -9.162886168127007e-13
+   -1.002036190244547e-11
+    8.519142210402354e-11
+   -4.832891079439459e-13
+   -9.103465728397491e-13
+   -2.121338766074267e-11
+    8.357903583358226e-11
+ 1.57e+10    
+    8.344127065965086e-11
+     -2.1161573639391e-11
+    8.522483025247911e-11
+   -9.193620469069734e-13
+   -1.002077890212854e-11
+     8.51881886311364e-11
+   -4.874113833784808e-13
+   -9.134033004133607e-13
+   -2.121348520418925e-11
+    8.357462970003014e-11
+ 1.58e+10    
+    8.343691955600744e-11
+   -2.116171660378015e-11
+     8.52216796542979e-11
+   -9.224450681445288e-13
+   -1.002120512844563e-11
+    8.518500137883216e-11
+   -4.915357746515419e-13
+   -9.164697016685348e-13
+   -2.121360051216985e-11
+    8.357025317431658e-11
+ 1.59e+10    
+    8.343259803446978e-11
+   -2.116187751789964e-11
+    8.521857505719382e-11
+   -9.255375125640989e-13
+   -1.002164060624519e-11
+     8.51818599894932e-11
+    -4.95661848566992e-13
+   -9.195456065235348e-13
+    -2.12137335456852e-11
+    8.356590594072405e-11
+ 1.6e+10     
+    8.342830578862481e-11
+   -2.116205633998745e-11
+    8.521551608791369e-11
+   -9.286392143195517e-13
+   -1.002208536072149e-11
+    8.517876410415298e-11
+    -4.99789177858574e-13
+   -9.226308470232554e-13
+    -2.12138842658902e-11
+    8.356158768629916e-11
+ 1.61e+10    
+    8.342404251477775e-11
+   -2.116225302858305e-11
+    8.521250237248417e-11
+   -9.317500096686789e-13
+    -1.00225394173704e-11
+    8.517571336257882e-11
+   -5.039173411943153e-13
+   -9.257252573296454e-13
+   -2.121405263411403e-11
+    8.355729810088364e-11
+ 1.62e+10    
+    8.341980791195817e-11
+   -2.116246754254206e-11
+     8.52095335362911e-11
+    -9.34869736960433e-13
+   -1.002300280194634e-11
+    8.517270740334846e-11
+    -5.08045923176696e-13
+   -9.288286737105331e-13
+    -2.12142386118766e-11
+    8.355303687713022e-11
+ 1.63e+10    
+    8.341560168191279e-11
+   -2.116269984104772e-11
+    8.520660920415092e-11
+   -9.379982366206953e-13
+   -1.002347554042029e-11
+    8.516974586392284e-11
+   -5.121745143387437e-13
+   -9.319409345267957e-13
+   -2.121444216090244e-11
+    8.354880371050455e-11
+ 1.64e+10    
+    8.341142352908583e-11
+    -2.11629498836198e-11
+    8.520372900037972e-11
+   -9.411353511366895e-13
+   -1.002395765893899e-11
+    8.516682838071483e-11
+   -5.163027111362154e-13
+   -9.350618802182547e-13
+   -2.121466324313161e-11
+    8.354459829927503e-11
+ 1.65e+10    
+    8.340727316058538e-11
+   -2.116321763012032e-11
+    8.520089254885743e-11
+   -9.442809250399925e-13
+   -1.002444918378541e-11
+    8.516395458915403e-11
+   -5.204301159360219e-13
+   -9.381913532880613e-13
+     -2.1214901820728e-11
+    8.354042034448893e-11
+ 1.66e+10    
+    8.340315028613955e-11
+   -2.116350304075686e-11
+    8.519809947308762e-11
+   -9.474348048883521e-13
+   -1.002495014134042e-11
+      8.5161124123748e-11
+   -5.245563370011032e-13
+   -9.413291982858418e-13
+   -2.121515785608518e-11
+    8.353626954993755e-11
+ 1.67e+10    
+    8.339905461804012e-11
+   -2.116380607608339e-11
+    8.519534939625427e-11
+   -9.505968392463511e-13
+   -1.002546055804581e-11
+    8.515833661814234e-11
+   -5.286809884718301e-13
+    -9.44475261789555e-13
+    -2.12154313118298e-11
+    8.353214562210924e-11
+ 1.68e+10    
+    8.339498587107706e-11
+   -2.116412669699882e-11
+    8.519264194127606e-11
+    -9.53766878664948e-13
+   -1.002598046036855e-11
+    8.515559170517547e-11
+   -5.328036903441446e-13
+   -9.476293923863063e-13
+    -2.12157221508228e-11
+    8.352804827013265e-11
+ 1.69e+10    
+    8.339094376246181e-11
+   -2.116446486474327e-11
+    8.518997673085692e-11
+   -9.569447756599812e-13
+   -1.002650987476661e-11
+     8.51528890169342e-11
+   -5.369240684445684e-13
+   -9.507914406519702e-13
+   -2.121603033615842e-11
+    8.352397720570882e-11
+ 1.7e+10     
+    8.338692801174209e-11
+   -2.116482054089229e-11
+    8.518735338753437e-11
+   -9.601303846897822e-13
+   -1.002704882765578e-11
+    8.515022818480524e-11
+   -5.410417544022094e-13
+   -9.539612591298366e-13
+   -2.121635583116141e-11
+    8.351993214303447e-11
+ 1.71e+10    
+    8.338293834070787e-11
+   -2.116519368734921e-11
+    8.518477153372657e-11
+   -9.633235621318045e-13
+   -1.002759734537831e-11
+    8.514760883952622e-11
+   -5.451563856179456e-13
+   -9.571387023083561e-13
+   -2.121669859938228e-11
+    8.351591279871649e-11
+ 1.72e+10    
+    8.337897447328956e-11
+   -2.116558426633589e-11
+    8.518223079177618e-11
+   -9.665241662585322e-13
+   -1.002815545417257e-11
+    8.514503061123519e-11
+   -5.492676052308739e-13
+    -9.60323626597912e-13
+   -2.121705860459089e-11
+    8.351191889167776e-11
+ 1.73e+10    
+    8.337503613544874e-11
+   -2.116599224038167e-11
+    8.517973078399384e-11
+   -9.697320572125298e-13
+   -1.002872318014439e-11
+    8.514249312951915e-11
+   -5.533750620822073e-13
+   -9.635158903068752e-13
+   -2.121743581076853e-11
+    8.350795014305543e-11
+ 1.74e+10    
+    8.337112305506239e-11
+   -2.116641757231082e-11
+    8.517727113269977e-11
+   -9.729470969808951e-13
+   -1.002930054923964e-11
+    8.513999602346165e-11
+   -5.574784106767166e-13
+   -9.667153536168269e-13
+   -2.121783018209855e-11
+    8.350400627609276e-11
+ 1.75e+10    
+    8.336723496180092e-11
+   -2.116686022522886e-11
+    8.517485146026352e-11
+     -9.7616914936901e-13
+   -1.002988758721818e-11
+    8.513753892168921e-11
+   -5.615773111418757e-13
+   -9.699218785571329e-13
+   -2.121824168295549e-11
+    8.350008701602365e-11
+ 1.76e+10    
+    8.336337158700142e-11
+    -2.11673201625076e-11
+    8.517247138914456e-11
+   -9.793980799736924e-13
+    -1.00304843196295e-11
+    8.513512145241883e-11
+   -5.656714291848039e-13
+   -9.731353289788536e-13
+   -2.121867027789351e-11
+    8.349619208995233e-11
+ 1.77e+10    
+     8.33595326635353e-11
+   -2.116779734776907e-11
+    8.517013054193029e-11
+   -9.826337561559217e-13
+   -1.003109077178932e-11
+    8.513274324350372e-11
+   -5.697604360471586e-13
+   -9.763555705280869e-13
+   -2.121911593163329e-11
+    8.349232122672725e-11
+ 1.78e+10    
+    8.335571792567292e-11
+   -2.116829174486861e-11
+    8.516782854137472e-11
+   -9.858760470129722e-13
+   -1.003170696875796e-11
+    8.513040392247982e-11
+   -5.738440084580839e-13
+   -9.795824706188243e-13
+   -2.121957860904839e-11
+    8.348847415681121e-11
+ 1.79e+10    
+    8.335192710894425e-11
+   -2.116880331787722e-11
+    8.516556501043612e-11
+   -9.891248233502322e-13
+   -1.003233293531988e-11
+    8.512810311661173e-11
+   -5.779218285853254e-13
+    -9.82815898405225e-13
+   -2.122005827515053e-11
+    8.348465061214665e-11
+ 1.8e+10     
+    8.334815994999644e-11
+   -2.116933203106304e-11
+    8.516333957231442e-11
+   -9.923799576526142e-13
+   -1.003296869596451e-11
+    8.512584045293957e-11
+   -5.819935839846339e-13
+   -9.860557247535968e-13
+   -2.122055489507446e-11
+     8.34808503260185e-11
+ 1.81e+10    
+    8.334441618645027e-11
+   -2.116987784887256e-11
+    8.516115185048917e-11
+   -9.956413240556392e-13
+   -1.003361427486872e-11
+    8.512361555832548e-11
+   -5.860589675475735e-13
+    -9.89301822213952e-13
+   -2.122106843406206e-11
+    8.347707303291371e-11
+ 1.82e+10    
+    8.334069555675415e-11
+    -2.11704407359115e-11
+    8.515900146875629e-11
+   -9.989087983162801e-13
+   -1.003426969588018e-11
+    8.512142805950091e-11
+   -5.901176774478264e-13
+   -9.925540649912172e-13
+   -2.122159885744628e-11
+    8.347331846837932e-11
+ 1.83e+10    
+    8.333699780003735e-11
+   -2.117102065692488e-11
+    8.515688805126641e-11
+    -1.00218225778355e-12
+   -1.003493498250242e-11
+    8.511927758311415e-11
+   -5.941694170861102e-13
+   -9.958123289162144e-13
+   -2.122214613063449e-11
+     8.34695863688787e-11
+ 1.84e+10    
+     8.33333226559633e-11
+   -2.117161757677771e-11
+    8.515481122256163e-11
+   -1.005461581368961e-12
+   -1.003561015788081e-11
+    8.511716375577812e-11
+   -5.982138950338171e-13
+   -9.990764914163654e-13
+   -2.122271021909172e-11
+     8.34658764716464e-11
+ 1.85e+10    
+    8.332966986458265e-11
+   -2.117223146043489e-11
+    8.515277060761397e-11
+   -1.008746649516796e-12
+   -1.003629524479001e-11
+    8.511508620411957e-11
+   -6.022508249754401e-13
+   -1.002346431486275e-12
+   -2.122329108832403e-11
+     8.34621885145439e-11
+ 1.86e+10    
+    8.332603916618734e-11
+    -2.11728622729418e-11
+    8.515076583186373e-11
+   -1.012037344174296e-12
+   -1.003699026562254e-11
+    8.511304455482786e-11
+   -6.062799256499341e-13
+   -1.005622029658101e-12
+   -2.122388870386147e-11
+    8.345852223591416e-11
+ 1.87e+10    
+    8.332243030116623e-11
+   -2.117350997940463e-11
+    8.514879652125758e-11
+    -1.01533354876184e-12
+   -1.003769524237844e-11
+    8.511103843470513e-11
+   -6.103009207910566e-13
+   -1.008903167971853e-12
+   -2.122450303124154e-11
+    8.345487737443783e-11
+ 1.88e+10    
+    8.331884300986205e-11
+   -2.117417454497122e-11
+    8.514686230228806e-11
+   -1.018635148143026e-12
+   -1.003841019665631e-11
+    8.510906747071684e-11
+   -6.143135390668015e-13
+   -1.012189729945624e-12
+   -2.122513403599267e-11
+    8.345125366899045e-11
+ 1.89e+10    
+    8.331527703243116e-11
+    -2.11748559348123e-11
+    8.514496280203296e-11
+   -1.021942028594819e-12
+   -1.003913514964515e-11
+    8.510713129004316e-11
+   -6.183175140180315e-13
+   -1.015481600545794e-12
+   -2.122578168361801e-11
+    8.344765085850143e-11
+ 1.9e+10     
+    8.331173210870621e-11
+    -2.11755541141029e-11
+      8.5143097648195e-11
+   -1.025254077777748e-12
+   -1.003987012211754e-11
+    8.510522952013033e-11
+   -6.223125839963295e-13
+   -1.018778666157221e-12
+   -2.122644593957965e-11
+    8.344406868181503e-11
+ 1.91e+10    
+    8.330820797806195e-11
+   -2.117626904800495e-11
+    8.514126646914271e-11
+    -1.02857118470618e-12
+   -1.004061513442369e-11
+    8.510336178874398e-11
+   -6.262984921012436e-13
+   -1.022080814553503e-12
+   -2.122712676928335e-11
+    8.344050687755456e-11
+ 1.92e+10    
+    8.330470437928458e-11
+   -2.117700070164963e-11
+    8.513946889395069e-11
+   -1.031893239718696e-12
+   -1.004137020648654e-11
+    8.510152772402191e-11
+   -6.302749861169303e-13
+   -1.025387934867267e-12
+   -2.122782413806374e-11
+    8.343696518398961e-11
+ 1.93e+10    
+    8.330122105044622e-11
+   -2.117774904012144e-11
+    8.513770455244195e-11
+   -1.035220134448641e-12
+   -1.004213535779787e-11
+    8.509972695452808e-11
+   -6.342418184482857e-13
+   -1.028699917560648e-12
+   -2.122853801117029e-11
+    8.343344333890679e-11
+ 1.94e+10    
+    8.329775772878286e-11
+   -2.117851402844233e-11
+    8.513597307522893e-11
+   -1.038551761794768e-12
+   -1.004291060741531e-11
+    8.509795910930693e-11
+   -6.381987460566974e-13
+   -1.032016654395761e-12
+   -2.122926835375382e-11
+    8.342994107948429e-11
+ 1.95e+10    
+    8.329431415057793e-11
+   -2.117929563155699e-11
+     8.51342740937566e-11
+   -1.041888015892241e-12
+   -1.004369597396008e-11
+    8.509622381793865e-11
+   -6.421455303953706e-13
+   -1.035338038405512e-12
+   -2.123001513085393e-11
+    8.342645814217145e-11
+ 1.96e+10    
+    8.329089005105188e-11
+   -2.118009381431925e-11
+    8.513260724034484e-11
+   -1.045228792083675e-12
+   -1.004449147561593e-11
+    8.509452071059438e-11
+   -6.460819373444619e-13
+   -1.038663963864396e-12
+   -2.123077830738724e-11
+    8.342299426257286e-11
+ 1.97e+10    
+     8.32874851642556e-11
+   -2.118090854147906e-11
+    8.513097214823211e-11
+   -1.048573986890534e-12
+   -1.004529713012849e-11
+    8.509284941809218e-11
+   -6.500077371458999e-13
+   -1.041994326259733e-12
+    -2.12315578481364e-11
+    8.341954917533763e-11
+ 1.98e+10    
+    8.328409922297173e-11
+   -2.118173977767092e-11
+    8.512936845161878e-11
+   -1.051923497984782e-12
+   -1.004611295480566e-11
+    8.509120957195358e-11
+    -6.53922704338118e-13
+   -1.045329022262912e-12
+   -2.123235371774021e-11
+    8.341612261405341e-11
+ 1.99e+10    
+    8.328073195862106e-11
+    -2.11825874874032e-11
+    8.512779578571181e-11
+   -1.055277224160832e-12
+   -1.004693896651867e-11
+    8.508960080446063e-11
+   -6.578266176906493e-13
+   -1.048667949701089e-12
+   -2.123316588068484e-11
+    8.341271431114806e-11
+ 2e+10       
+    8.327738310117629e-11
+   -2.118345163504871e-11
+    8.512625378676839e-11
+   -1.058635065307738e-12
+   -1.004777518170377e-11
+    8.508802274871207e-11
+   -6.617192601387326e-13
+   -1.052011007529015e-12
+   -2.123399430129562e-11
+     8.34093239977951e-11
+ 2.01e+10    
+    8.327405237908133e-11
+    -2.11843321848363e-11
+    8.512474209214139e-11
+   -1.061996922381827e-12
+   -1.004862161636457e-11
+    8.508647503868128e-11
+   -6.656004187178682e-13
+   -1.055358095801305e-12
+    -2.12348389437303e-11
+    8.340595140382658e-11
+ 2.02e+10    
+    8.327073951917887e-11
+   -2.118522910084387e-11
+    8.512326034032381e-11
+   -1.065362697379561e-12
+    -1.00494782860751e-11
+    8.508495730927357e-11
+   -6.694698844985396e-13
+   -1.058709115644877e-12
+   -2.123569977197357e-11
+    8.340259625765319e-11
+ 2.03e+10    
+    8.326744424664375e-11
+   -2.118614234699234e-11
+    8.512180817099406e-11
+   -1.068732293310873e-12
+   -1.005034520598339e-11
+    8.508346919638357e-11
+   -6.733274525209537e-13
+   -1.062063969231853e-12
+   -2.123657674983216e-11
+    8.339925828618923e-11
+ 2.04e+10    
+    8.326416628492502e-11
+    -2.11870718870414e-11
+    8.512038522506179e-11
+   -1.072105614172769e-12
+   -1.005122239081555e-11
+    8.508201033695293e-11
+   -6.771729217300614e-13
+   -1.065422559752754e-12
+   -2.123746984093155e-11
+    8.339593721478597e-11
+ 2.05e+10    
+     8.32609053556937e-11
+   -2.118801768458568e-11
+     8.51189911447121e-11
+     -1.0754825649234e-12
+   -1.005210985488031e-11
+    8.508058036902773e-11
+   -6.810060949107189e-13
+   -1.068784791390051e-12
+   -2.123837900871375e-11
+    8.339263276717152e-11
+ 2.06e+10    
+    8.325766117879917e-11
+   -2.118897970305317e-11
+     8.51176255734525e-11
+   -1.078863051456509e-12
+   -1.005300761207427e-11
+    8.507917893181583e-11
+   -6.848267786231238e-13
+   -1.072150569292143e-12
+   -2.123930421643597e-11
+    8.338934466539691e-11
+ 2.07e+10    
+    8.325443347223212e-11
+   -2.118995790570409e-11
+    8.511628815615715e-11
+   -1.082246980576226e-12
+   -1.005391567588733e-11
+     8.50778056657442e-11
+   -6.886347831386278e-13
+   -1.075519799547681e-12
+   -2.124024542717111e-11
+    8.338607262979157e-11
+ 2.08e+10    
+    8.325122195209608e-11
+   -2.119095225563162e-11
+    8.511497853911292e-11
+   -1.085634259972426e-12
+   -1.005483405940856e-11
+    8.507646021251618e-11
+   -6.924299223757823e-13
+   -1.078892389160335e-12
+   -2.124120260380883e-11
+    8.338281637892363e-11
+ 2.09e+10    
+    8.324802633258521e-11
+   -2.119196271576345e-11
+    8.511369637006404e-11
+   -1.089024798196381e-12
+   -1.005576277533251e-11
+    8.507514221516722e-11
+   -6.962120138368571e-13
+    -1.08226824602394e-12
+   -2.124217570905789e-11
+    8.337957562956876e-11
+ 2.1e+10     
+    8.324484632597044e-11
+   -2.119298924886504e-11
+    8.511244129825788e-11
+   -1.092418504636899e-12
+   -1.005670183596591e-11
+    8.507385131812223e-11
+   -6.999808785447412e-13
+   -1.085647278898088e-12
+   -2.124316470545018e-11
+    8.337635009668626e-11
+ 2.11e+10    
+    8.324168164259264e-11
+   -2.119403181754377e-11
+    8.511121297448927e-11
+   -1.095815289496916e-12
+   -1.005765125323439e-11
+    8.507258716725042e-11
+   -7.037363409802961e-13
+   -1.089029397384173e-12
+    -2.12441695553453e-11
+    8.337313949340265e-11
+ 2.12e+10    
+    8.323853199086306e-11
+   -2.119509038425439e-11
+    8.511001105114485e-11
+   -1.099215063770523e-12
+   -1.005861103868986e-11
+    8.507134940992116e-11
+   -7.074782290201911e-13
+   -1.092414511901793e-12
+   -2.124519022093656e-11
+    8.336994353100126e-11
+ 2.13e+10    
+    8.323539707727121e-11
+   -2.119616491130575e-11
+    8.510883518224792e-11
+    -1.10261773922045e-12
+   -1.005958120351777e-11
+    8.507013769505812e-11
+   -7.112063738752535e-13
+   -1.095802533665715e-12
+   -2.124622666425814e-11
+    8.336676191892062e-11
+ 2.14e+10    
+     8.32322766063999e-11
+   -2.119725536086869e-11
+    8.510768502350121e-11
+   -1.106023228356004e-12
+   -1.006056175854483e-11
+    8.506895167319355e-11
+   -7.149206100293589e-13
+   -1.099193374663187e-12
+   -2.124727884719327e-11
+    8.336359436475888e-11
+ 2.15e+10    
+    8.322917028094682e-11
+   -2.119836169498492e-11
+    8.510656023233108e-11
+   -1.109431444411465e-12
+   -1.006155271424678e-11
+    8.506779099652152e-11
+   -7.186207751788792e-13
+   -1.102586947631744e-12
+   -2.124834673148362e-11
+    8.336044057428566e-11
+ 2.16e+10    
+    8.322607780175365e-11
+   -2.119948387557708e-11
+    8.510546046792929e-11
+    -1.11284230132495e-12
+   -1.006255408075635e-11
+    8.506665531894987e-11
+   -7.223067101727211e-13
+   -1.105983166037506e-12
+   -2.124943027873939e-11
+    8.335730025146048e-11
+ 2.17e+10    
+    8.322299886784119e-11
+   -2.120062186446006e-11
+    8.510438539129619e-11
+   -1.116255713717701e-12
+   -1.006356586787144e-11
+    8.506554429615197e-11
+   -7.259782589529789e-13
+   -1.109381944053859e-12
+   -2.125052945045082e-11
+    8.335417309845821e-11
+ 2.18e+10    
+    8.321993317645108e-11
+   -2.120177562335277e-11
+    8.510333466528098e-11
+   -1.119671596873925e-12
+   -1.006458808506316e-11
+    8.506445758561759e-11
+   -7.296352684961951e-13
+   -1.112783196540655e-12
+   -2.125164420800041e-11
+    8.335105881570071e-11
+ 2.19e+10    
+    8.321688042309393e-11
+   -2.120294511389152e-11
+    8.510230795462354e-11
+   -1.123089866721001e-12
+   -1.006562074148431e-11
+    8.506339484670238e-11
+   -7.332775887552855e-13
+    -1.11618683902386e-12
+   -2.125277451267629e-11
+    8.334795710189519e-11
+ 2.2e+10     
+    8.321384030160306e-11
+    -2.12041302976438e-11
+    8.510130492599381e-11
+    -1.12651043981017e-12
+   -1.006666384597751e-11
+    8.506235574067587e-11
+   -7.369050726021327e-13
+   -1.119592787675669e-12
+   -2.125392032568591e-11
+    8.334486765407873e-11
+ 2.21e+10    
+    8.321081250419474e-11
+   -2.120533113612324e-11
+     8.51003252480315e-11
+   -1.129933233297728e-12
+   -1.006771740708384e-11
+    8.506133993077018e-11
+   -7.405175757708229e-13
+   -1.123000959295046e-12
+   -2.125508160817153e-11
+    8.334179016766799e-11
+ 2.22e+10    
+    8.320779672153311e-11
+   -2.120654759080522e-11
+    8.509936859138406e-11
+   -1.133358164926607e-12
+   -1.006878143305102e-11
+    8.506034708222499e-11
+   -7.441149568016197e-13
+   -1.126411271288768e-12
+    -2.12562583212253e-11
+     8.33387243365159e-11
+ 2.23e+10    
+    8.320479264280032e-11
+   -2.120777962314313e-11
+     8.50984346287445e-11
+   -1.136785153008497e-12
+   -1.006985593184195e-11
+    8.505937686233371e-11
+   -7.476970769855923e-13
+   -1.129823641652914e-12
+   -2.125745042590618e-11
+     8.33356698529724e-11
+ 2.24e+10    
+    8.320179995577254e-11
+    -2.12090271945856e-11
+    8.509752303488784e-11
+   -1.140214116406303e-12
+   -1.007094091114305e-11
+    8.505842894048702e-11
+   -7.512638003100024e-13
+   -1.133237988954792e-12
+    -2.12586578832567e-11
+    8.333262640795204e-11
+ 2.25e+10    
+    8.319881834689969e-11
+   -2.121029026659404e-11
+     8.50966334867068e-11
+   -1.143644974517151e-12
+   -1.007203637837261e-11
+    8.505750298821544e-11
+   -7.548149934043723e-13
+   -1.136654232315342e-12
+   -2.125988065432077e-11
+    8.332959369100438e-11
+ 2.26e+10    
+    8.319584750138978e-11
+   -2.121156880066094e-11
+    8.509576566324638e-11
+   -1.147077647255775e-12
+   -1.007314234068914e-11
+     8.50565986792311e-11
+   -7.583505254873017e-13
+   -1.140072291391962e-12
+   -2.126111870016205e-11
+    8.332657139039169e-11
+ 2.27e+10    
+    8.319288710329765e-11
+   -2.121286275832866e-11
+    8.509491924573745e-11
+   -1.150512055038353e-12
+   -1.007425880499958e-11
+    8.505571568946731e-11
+   -7.618702683140231e-13
+   -1.143492086361794e-12
+   -2.126237198188254e-11
+     8.33235591931684e-11
+ 2.28e+10    
+    8.318993683561694e-11
+   -2.121417210120848e-11
+    8.509409391762899e-11
+   -1.153948118766783e-12
+   -1.007538577796744e-11
+    8.505485369711731e-11
+   -7.653740961246966e-13
+   -1.146913537905449e-12
+   -2.126364046064186e-11
+    8.332055678526676e-11
+ 2.29e+10    
+    8.318699638037569e-11
+   -2.121549679100023e-11
+    8.509328936462019e-11
+   -1.157385759813356e-12
+     -1.0076523266021e-11
+    8.505401238267175e-11
+   -7.688618855934271e-13
+   -1.150336567191159e-12
+   -2.126492409767681e-11
+    8.331756385158477e-11
+ 2.3e+10     
+    8.318406541873584e-11
+   -2.121683678951225e-11
+    8.509250527468976e-11
+   -1.160824900005887e-12
+   -1.007767127536105e-11
+    8.505319142895413e-11
+   -7.723335157780683e-13
+   -1.153761095859362e-12
+   -2.126622285432136e-11
+    8.331458007607883e-11
+ 2.31e+10    
+     8.31811436310939e-11
+   -2.121819205868127e-11
+    8.509174133812542e-11
+   -1.164265461613211e-12
+   -1.007882981196902e-11
+    8.505239052115553e-11
+   -7.757888680707433e-13
+   -1.157187046007678e-12
+   -2.126753669202668e-11
+    8.331160514185864e-11
+ 2.32e+10    
+    8.317823069718572e-11
+   -2.121956256059295e-11
+     8.50909972475521e-11
+   -1.167707367331126e-12
+   -1.007999888161453e-11
+    8.505160934686702e-11
+   -7.792278261491379e-13
+   -1.160614340176377e-12
+   -2.126886557238156e-11
+    8.330863873128557e-11
+ 2.33e+10    
+    8.317532629619286e-11
+   -2.122094825750221e-11
+    8.509027269795801e-11
+   -1.171150540268691e-12
+   -1.008117848986303e-11
+    8.505084759611108e-11
+    -7.82650275928525e-13
+   -1.164042901334188e-12
+   -2.127020945713298e-11
+    8.330568052607347e-11
+ 2.34e+10    
+    8.317243010685022e-11
+   -2.122234911185361e-11
+    8.508956738672056e-11
+   -1.174594903934954e-12
+   -1.008236864208331e-11
+    8.505010496137206e-11
+   -7.860561055145582e-13
+   -1.167472652864506e-12
+   -2.127156830820664e-11
+    8.330273020739169e-11
+ 2.35e+10    
+    8.316954180755661e-11
+   -2.122376508630208e-11
+    8.508888101363015e-11
+   -1.178040382226032e-12
+   -1.008356934345485e-11
+     8.50493811376239e-11
+   -7.894452051568138e-13
+   -1.170903518552043e-12
+   -2.127294208772768e-11
+    8.329978745597046e-11
+ 2.36e+10    
+    8.316666107648537e-11
+   -2.122519614373317e-11
+    8.508821328091334e-11
+   -1.181486899412582e-12
+   -1.008478059897483e-11
+    8.504867582235687e-11
+   -7.928174672030568e-13
+   -1.174335422569856e-12
+   -2.127433075804102e-11
+    8.329685195220688e-11
+ 2.37e+10    
+    8.316378759169647e-11
+   -2.122664224728343e-11
+    8.508756389325453e-11
+   -1.184934380127628e-12
+   -1.008600241346531e-11
+    8.504798871560334e-11
+   -7.961727860542857e-13
+   -1.177768289466707e-12
+   -2.127573428173233e-11
+    8.329392337627429e-11
+ 2.38e+10    
+    8.316092103124973e-11
+   -2.122810336036071e-11
+    8.508693255781607e-11
+   -1.188382749354758e-12
+   -1.008723479157999e-11
+    8.504731951996104e-11
+    -7.99511058120494e-13
+    -1.18120204415486e-12
+   -2.127715262164787e-11
+    8.329100140823063e-11
+ 2.39e+10    
+    8.315806107331724e-11
+   -2.122957944666386e-11
+    8.508631898425754e-11
+   -1.191831932416659e-12
+   -1.008847773781086e-11
+    8.504666794061542e-11
+   -8.028321817771689e-13
+   -1.184636611898184e-12
+   -2.127858574091499e-11
+    8.328808572812875e-11
+ 2.4e+10     
+    8.315520739629753e-11
+   -2.123107047020265e-11
+    8.508572288475349e-11
+   -1.195281854964017e-12
+   -1.008973125649479e-11
+    8.504603368536008e-11
+   -8.061360573225383e-13
+   -1.188071918300686e-12
+   -2.128003360296196e-11
+    8.328517601612737e-11
+ 2.41e+10    
+    8.315235967892821e-11
+   -2.123257639531692e-11
+    8.508514397400963e-11
+   -1.198732442964732e-12
+   -1.009099535181973e-11
+    8.504541646461632e-11
+   -8.094225869355312e-13
+    -1.19150788929531e-12
+   -2.128149617153766e-11
+    8.328227195260175e-11
+ 2.42e+10    
+    8.314951760039884e-11
+   -2.123409718669569e-11
+    8.508458196927822e-11
+   -1.202183622693453e-12
+   -1.009227002783094e-11
+    8.504481599145008e-11
+   -8.126916746344625e-13
+   -1.194944451133139e-12
+    -2.12829734107308e-11
+    8.327937321825462e-11
+ 2.43e+10    
+     8.31466808404632e-11
+    -2.12356328093957e-11
+    8.508403659037192e-11
+   -1.205635320721458e-12
+   -1.009355528843696e-11
+      8.5044231981588e-11
+   -8.159432262364392e-13
+   -1.198381530372906e-12
+   -2.128446528498877e-11
+    8.327647949422693e-11
+ 2.44e+10    
+    8.314384907955074e-11
+   -2.123718322885951e-11
+    8.508350755967639e-11
+   -1.209087463906862e-12
+   -1.009485113741534e-11
+    8.504366415343254e-11
+   -8.191771493174677e-13
+   -1.201819053870829e-12
+    -2.12859717591363e-11
+    8.327359046220823e-11
+ 2.45e+10    
+    8.314102199887664e-11
+   -2.123874841093311e-11
+    8.508299460216108e-11
+   -1.212539979385046e-12
+   -1.009615757841826e-11
+     8.50431122280741e-11
+   -8.223933531732719e-13
+    -1.20525694877079e-12
+   -2.128749279839316e-11
+    8.327070580454569e-11
+ 2.46e+10    
+    8.313819928055028e-11
+   -2.124032832188296e-11
+    8.508249744538986e-11
+   -1.215992794559447e-12
+   -1.009747461497807e-11
+    8.504257592930329e-11
+   -8.255917487808134e-13
+   -1.208695142494744e-12
+   -2.128902836839199e-11
+    8.326782520435298e-11
+ 2.47e+10    
+    8.313538060768337e-11
+   -2.124192292841251e-11
+    8.508201581952898e-11
+   -1.219445837092672e-12
+   -1.009880225051224e-11
+    8.504205498361982e-11
+   -8.287722487604615e-13
+   -1.212133562733561e-12
+   -2.129057843519481e-11
+    8.326494834561716e-11
+ 2.48e+10    
+     8.31325656644947e-11
+   -2.124353219767814e-11
+    8.508154945735518e-11
+   -1.222899034897783e-12
+   -1.010014048832877e-11
+     8.50415491202425e-11
+   -8.319347673389141e-13
+   -1.215572137438027e-12
+   -2.129214296530986e-11
+     8.32620749133052e-11
+ 2.49e+10    
+    8.312975413641479e-11
+    -2.12451560973043e-11
+    8.508109809426113e-11
+   -1.226352316129965e-12
+   -1.010148933163076e-11
+     8.50410580711151e-11
+   -8.350792203127334e-13
+   -1.219010794810202e-12
+   -2.129372192570683e-11
+    8.325920459346751e-11
+ 2.5e+10     
+    8.312694571018645e-11
+   -2.124679459539812e-11
+    8.508066146826069e-11
+   -1.229805609178382e-12
+    -1.01028487835213e-11
+    8.504058157091244e-11
+   -8.382055250125691e-13
+   -1.222449463295085e-12
+   -2.129531528383224e-11
+    8.325633707334121e-11
+ 2.51e+10    
+    8.312414007396494e-11
+   -2.124844766056341e-11
+     8.50802393199928e-11
+   -1.233258842658306e-12
+   -1.010421884700791e-11
+    8.504011935704473e-11
+    -8.41313600268038e-13
+   -1.225888071572449e-12
+   -2.129692300762376e-11
+    8.325347204145026e-11
+ 2.52e+10    
+    8.312133691741458e-11
+   -2.125011526191361e-11
+     8.50798313927233e-11
+   -1.236711945403545e-12
+   -1.010559952500687e-11
+    8.503967116966022e-11
+   -8.444033663732747e-13
+   -1.229326548549038e-12
+   -2.129854506552383e-11
+      8.3250609187704e-11
+ 2.53e+10    
+     8.31185359318033e-11
+   -2.125179736908434e-11
+    8.507943743234664e-11
+   -1.240164846459063e-12
+   -1.010699082034739e-11
+    8.503923675164696e-11
+   -8.474747450530916e-13
+   -1.232764823350953e-12
+    -2.13001814264928e-11
+    8.324774820349375e-11
+ 2.54e+10    
+    8.311573681009453e-11
+   -2.125349395224514e-11
+    8.507905718738572e-11
+   -1.243617475073841e-12
+    -1.01083927357756e-11
+    8.503881584863259e-11
+    -8.50527659429792e-13
+    -1.23620282531632e-12
+   -2.130183206002095e-11
+    8.324488878178577e-11
+ 2.55e+10    
+    8.311293924703599e-11
+   -2.125520498211019e-11
+    8.507869040899092e-11
+      -1.247069760694e-12
+   -1.010980527395845e-11
+    8.503840820898384e-11
+   -8.535620339906143e-13
+   -1.239640483988198e-12
+   -2.130349693614015e-11
+    8.324203061721337e-11
+ 2.56e+10    
+    8.311014293924613e-11
+    -2.12569304299486e-11
+    8.507833685093796e-11
+   -1.250521632956097e-12
+   -1.011122843748726e-11
+    8.503801358380348e-11
+   -8.565777945557905e-13
+   -1.243077729107699e-12
+   -2.130517602543449e-11
+    8.323917340616534e-11
+ 2.57e+10    
+    8.310734758529687e-11
+   -2.125867026759341e-11
+    8.507799626962387e-11
+   -1.253973021680705e-12
+   -1.011266222888115e-11
+    8.503763172692676e-11
+   -8.595748682472078e-13
+    -1.24651449060737e-12
+   -2.130686929904997e-11
+    8.323631684687106e-11
+ 2.58e+10    
+    8.310455288579413e-11
+   -2.126042446745054e-11
+    8.507766842406381e-11
+    -1.25742385686611e-12
+   -1.011410665059064e-11
+    8.503726239491727e-11
+   -8.625531834576872e-13
+   -1.249950698604724e-12
+   -2.130857672870402e-11
+    8.323346063948449e-11
+ 2.59e+10    
+    8.310175854345487e-11
+     -2.1262193002506e-11
+    8.507735307588405e-11
+   -1.260874068682338e-12
+   -1.011556170500051e-11
+    8.503690534705985e-11
+   -8.655126698208492e-13
+   -1.253386283396081e-12
+   -2.131029828669338e-11
+    8.323060448616355e-11
+ 2.6e+10     
+    8.309896426318054e-11
+   -2.126397584633312e-11
+    8.507704998931683e-11
+   -1.264323587465233e-12
+   -1.011702739443305e-11
+    8.503656034535406e-11
+   -8.684532581815646e-13
+   -1.256821175450564e-12
+    -2.13120339459018e-11
+    8.322774809114735e-11
+ 2.61e+10    
+    8.309616975212815e-11
+   -2.126577297309839e-11
+    8.507675893119175e-11
+   -1.267772343710861e-12
+   -1.011850372115079e-11
+    8.503622715450572e-11
+   -8.713748805669945e-13
+   -1.260255305404259e-12
+   -2.131378367980665e-11
+       8.322489116083e-11
+ 2.62e+10    
+    8.309337471977711e-11
+    -2.12675843575666e-11
+    8.507647967092738e-11
+   -1.271220268070021e-12
+   -1.011999068735926e-11
+    8.503590554191756e-11
+   -8.742774701581901e-13
+   -1.263688604054657e-12
+   -2.131554746248474e-11
+    8.322203340383158e-11
+ 2.63e+10    
+    8.309057887799392e-11
+   -2.126940997510551e-11
+    8.507621198052242e-11
+   -1.274667291342948e-12
+   -1.012148829520961e-11
+    8.503559527767808e-11
+   -8.771609612622597e-13
+   -1.267121002355228e-12
+   -2.131732526861716e-11
+    8.321917453106522e-11
+ 2.64e+10    
+    8.308778194109244e-11
+   -2.127124980168916e-11
+    8.507595563454436e-11
+    -1.27811334447421e-12
+   -1.012299654680103e-11
+    8.503529613455126e-11
+     -8.8002528928511e-13
+   -1.270552431410148e-12
+   -2.131911707349381e-11
+    8.321631425580254e-11
+ 2.65e+10    
+    8.308498362589125e-11
+   -2.127310381390078e-11
+      8.5075710410119e-11
+   -1.281558358547773e-12
+   -1.012451544418306e-11
+    8.503500788796301e-11
+   -8.828703907046966e-13
+   -1.273982822469312e-12
+   -2.132092285301646e-11
+    8.321345229373329e-11
+ 2.66e+10    
+    8.308218365176821e-11
+   -2.127497198893456e-11
+    8.507547608691664e-11
+    -1.28500226478224e-12
+   -1.012604498935763e-11
+    8.503473031598794e-11
+   -8.856962030448561e-13
+   -1.277412106923409e-12
+   -2.132274258370135e-11
+    8.321058836302458e-11
+ 2.67e+10    
+    8.307938174071074e-11
+   -2.127685430459706e-11
+    8.507525244714092e-11
+   -1.288444994526207e-12
+   -1.012758518428137e-11
+    8.503446319933551e-11
+   -8.885026648496523e-13
+   -1.280840216299187e-12
+   -2.132457624268111e-11
+    8.320772218437461e-11
+ 2.68e+10    
+    8.307657761736337e-11
+   -2.127875073930731e-11
+    8.507503927551342e-11
+   -1.291886479253822e-12
+   -1.012913603086732e-11
+    8.503420632133405e-11
+   -8.912897156582519e-13
+   -1.284267082254944e-12
+   -2.132642380770537e-11
+    8.320485348106407e-11
+ 2.69e+10    
+    8.307377100907227e-11
+   -2.128066127209665e-11
+    8.507483635925981e-11
+   -1.295326650560475e-12
+   -1.013069753098681e-11
+      8.5033959467915e-11
+   -8.940572959803263e-13
+   -1.287692636576121e-12
+   -2.132828525714131e-11
+    8.320198197900486e-11
+ 2.7e+10     
+    8.307096164592542e-11
+    -2.12825858826073e-11
+    8.507464348809376e-11
+    -1.29876544015866e-12
+   -1.013226968647115e-11
+    8.503372242759604e-11
+   -8.968053472719368e-13
+    -1.29111681117103e-12
+   -2.133016056997275e-11
+    8.319910740678389e-11
+ 2.71e+10    
+    8.306814926079079e-11
+   -2.128452455109056e-11
+    8.507446045420098e-11
+   -1.302202779873921e-12
+    -1.01338524991132e-11
+    8.503349499146308e-11
+   -8.995338119119998e-13
+   -1.294539538066775e-12
+   -2.133204972579887e-11
+    8.319622949570544e-11
+ 2.72e+10    
+    8.306533358935056e-11
+   -2.128647725840413e-11
+    8.507428705222223e-11
+   -1.305638601641022e-12
+   -1.013544597066883e-11
+    8.503327695315188e-11
+   -9.022426331791441e-13
+   -1.297960749405309e-12
+   -2.133395270483194e-11
+    8.319334797982888e-11
+ 2.73e+10    
+    8.306251437013245e-11
+   -2.128844398600867e-11
+    8.507412307923573e-11
+   -1.309072837500156e-12
+    -1.01370501028583e-11
+    8.503306810882865e-11
+   -9.049317552291598e-13
+     -1.3013803774396e-12
+   -2.133586948789468e-11
+    8.319046259600434e-11
+ 2.74e+10    
+    8.305969134453787e-11
+   -2.129042471596377e-11
+    8.507396833473876e-11
+   -1.312505419593394e-12
+   -1.013866489736752e-11
+     8.50328682571709e-11
+   -9.076011230728683e-13
+   -1.304798354529961e-12
+   -2.133780005641652e-11
+    8.318757308390461e-11
+ 2.75e+10    
+    8.305686425686719e-11
+   -2.129241943092308e-11
+    8.507382262062899e-11
+   -1.315936280161154e-12
+    -1.01402903558492e-11
+    8.503267719934536e-11
+   -9.102506825545217e-13
+   -1.308214613140501e-12
+   -2.133974439242915e-11
+    8.318467918605383e-11
+ 2.76e+10    
+    8.305403285434117e-11
+    -2.12944281141289e-11
+    8.507368574118485e-11
+   -1.319365351538856e-12
+   -1.014192647992401e-11
+    8.503249473898857e-11
+   -9.128803803306173e-13
+     -1.3116290858357e-12
+   -2.134170247856189e-11
+    8.318178064785395e-11
+ 2.77e+10    
+    8.305119688712125e-11
+   -2.129645074940613e-11
+    8.507355750304537e-11
+   -1.322792566153721e-12
+   -1.014357327118143e-11
+    8.503232068218381e-11
+   -9.154901638492417e-13
+   -1.315041705277113e-12
+   -2.134367429803572e-11
+    8.317887721760706e-11
+ 2.78e+10    
+    8.304835610832514e-11
+   -2.129848732115546e-11
+    8.507343771518979e-11
+   -1.326217856521588e-12
+   -1.014523073118081e-11
+     8.50321548374391e-11
+   -9.180799813298343e-13
+   -1.318452404220189e-12
+   -2.134565983465704e-11
+    8.317596864653592e-11
+ 2.79e+10    
+     8.30455102740403e-11
+   -2.130053781434606e-11
+    8.507332618891653e-11
+   -1.329641155243972e-12
+   -1.014689886145209e-11
+    8.503199701566467e-11
+   -9.206497817434175e-13
+   -1.321861115511208e-12
+   -2.134765907281084e-11
+    8.317305468880055e-11
+ 2.8e+10     
+    8.304265914333486e-11
+   -2.130260221450758e-11
+    8.507322273782124e-11
+   -1.333062395005131e-12
+   -1.014857766349654e-11
+    8.503184703014898e-11
+   -9.231995147932895e-13
+   -1.325267772084346e-12
+   -2.134967199745309e-11
+     8.31701351015134e-11
+ 2.81e+10    
+    8.303980247826604e-11
+    -2.13046805077218e-11
+     8.50731271777752e-11
+   -1.336481508569309e-12
+   -1.015026713878754e-11
+     8.50317046965357e-11
+   -9.257291308961416e-13
+   -1.328672306958813e-12
+   -2.135169859410262e-11
+    8.316720964475004e-11
+ 2.82e+10    
+    8.303694004388531e-11
+   -2.130677268061355e-11
+    8.507303932690276e-11
+   -1.339898428778031e-12
+   -1.015196728877108e-11
+    8.503156983279836e-11
+   -9.282385811636302e-13
+   -1.332074653236145e-12
+   -2.135373884883238e-11
+    8.316427808155882e-11
+ 2.83e+10    
+    8.303407160824154e-11
+   -2.130887872034098e-11
+    8.507295900555821e-11
+   -1.343313088547558e-12
+   -1.015367811486629e-11
+    8.503144225921672e-11
+   -9.307278173843694e-13
+   -1.335474744097562e-12
+   -2.135579274826025e-11
+    8.316134017796676e-11
+ 2.84e+10    
+    8.303119694238167e-11
+    -2.13109986145858e-11
+    8.507288603630287e-11
+    -1.34672542086637e-12
+   -1.015539961846599e-11
+    8.503132179835096e-11
+   -9.331967920063692e-13
+   -1.338872512801452e-12
+   -2.135786027953932e-11
+    8.315839570298404e-11
+ 2.85e+10    
+    8.302831582034906e-11
+   -2.131313235154242e-11
+    8.507282024388157e-11
+    -1.35013535879285e-12
+   -1.015713180093709e-11
+    8.503120827501682e-11
+   -9.356454581198676e-13
+   -1.342267892680914e-12
+   -2.135994143034748e-11
+    8.315544442860457e-11
+ 2.86e+10    
+    8.302542801917942e-11
+   -2.131527991990723e-11
+    8.507276145519856e-11
+   -1.353542835452933e-12
+   -1.015887466362088e-11
+    8.503110151625948e-11
+   -9.380737694406068e-13
+    -1.34566081714148e-12
+    -2.13620361888769e-11
+      8.3152486129806e-11
+ 2.87e+10    
+    8.302253331889456e-11
+   -2.131744130886687e-11
+    8.507270949929323e-11
+   -1.356947784037962e-12
+   -1.016062820783334e-11
+    8.503100135132751e-11
+   -9.404816802935227e-13
+   -1.349051219658828e-12
+   -2.136414454382254e-11
+    8.314952058454566e-11
+ 2.88e+10    
+    8.301963150249463e-11
+   -2.131961650808673e-11
+      8.5072664207316e-11
+   -1.360350137802589e-12
+   -1.016239243486546e-11
+    8.503090761164693e-11
+   -9.428691455968066e-13
+   -1.352439033776655e-12
+   -2.136626648437085e-11
+    8.314654757375599e-11
+ 2.89e+10    
+    8.301672235594738e-11
+   -2.132180550769849e-11
+    8.507262541250328e-11
+    -1.36374983006275e-12
+   -1.016416734598332e-11
+    8.503082013079433e-11
+   -9.452361208464223e-13
+    -1.35582419310461e-12
+    -2.13684020001874e-11
+     8.31435668813363e-11
+ 2.9e+10     
+    8.301380566817614e-11
+   -2.132400829828757e-11
+    8.507259295015291e-11
+   -1.367146794193744e-12
+   -1.016595294242836e-11
+    8.503073874447004e-11
+   -9.475825621009556e-13
+   -1.359206631316347e-12
+   -2.137055108140471e-11
+    8.314057829414383e-11
+ 2.91e+10    
+    8.301088123104591e-11
+   -2.132622487088008e-11
+    8.507256665759829e-11
+    -1.37054096362841e-12
+   -1.016774922541741e-11
+    8.503066329047179e-11
+    -9.49908425966932e-13
+   -1.362586282147582e-12
+   -2.137271371860939e-11
+    8.313758160198208e-11
+ 2.92e+10    
+    8.300794883934747e-11
+   -2.132845521692983e-11
+    8.507254637418409e-11
+   -1.373932271855331e-12
+   -1.016955619614279e-11
+    8.503059360866652e-11
+   -9.522136695844642e-13
+   -1.365963079394365e-12
+    -2.13748899028288e-11
+    8.313457659758752e-11
+ 2.93e+10    
+    8.300500829078006e-11
+   -2.133069932830443e-11
+    8.507253194124006e-11
+   -1.377320652417227e-12
+   -1.017137385577235e-11
+    8.503052954096435e-11
+   -9.544982506132965e-13
+    -1.36933695691126e-12
+   -2.137707962551786e-11
+    8.313156307661417e-11
+ 2.94e+10    
+    8.300205938593253e-11
+    -2.13329571972717e-11
+    8.507252320205512e-11
+   -1.380706038909293e-12
+   -1.017320220544938e-11
+    8.503047093129014e-11
+   -9.567621272192457e-13
+   -1.372707848609776e-12
+   -2.137928287854516e-11
+    8.312854083761733e-11
+ 2.95e+10    
+    8.299910192826227e-11
+   -2.133522881648537e-11
+    8.507252000185271e-11
+   -1.384088364977708e-12
+   -1.017504124629272e-11
+    8.503041762555652e-11
+   -9.590052580609939e-13
+   -1.376075688456761e-12
+   -2.138149965417884e-11
+    8.312550968203478e-11
+ 2.96e+10    
+    8.299613572407367e-11
+   -2.133751417897083e-11
+    8.507252218776414e-11
+   -1.387467564318177e-12
+   -1.017689097939656e-11
+    8.503036947163604e-11
+   -9.612276022772732e-13
+   -1.379440410472897e-12
+   -2.138372994507241e-11
+      8.3122469414167e-11
+ 2.97e+10    
+    8.299316058249483e-11
+    -2.13398132781105e-11
+    8.507252960880256e-11
+   -1.390843570674585e-12
+   -1.017875140583036e-11
+    8.503032631933383e-11
+   -9.634291194743913e-13
+   -1.382801948731296e-12
+   -2.138597374425017e-11
+    8.311941984115571e-11
+ 2.98e+10    
+    8.299017631545251e-11
+   -2.134212610762905e-11
+    8.507254211583728e-11
+   -1.394216317837661e-12
+   -1.018062252663878e-11
+    8.503028802035947e-11
+   -9.656097697141317e-13
+   -1.386160237356116e-12
+   -2.138823104509226e-11
+    8.311636077296082e-11
+ 2.99e+10    
+    8.298718273764697e-11
+   -2.134445266157851e-11
+    8.507255956156799e-11
+   -1.397585739643782e-12
+   -1.018250434284147e-11
+    8.503025442829973e-11
+   -9.677695135020168e-13
+   -1.389515210521302e-12
+   -2.139050184132006e-11
+    8.311329202233689e-11
+ 3e+10       
+    8.298417966652462e-11
+   -2.134679293432312e-11
+    8.507258180049818e-11
+   -1.400951769973765e-12
+   -1.018439685543293e-11
+    8.503022539859044e-11
+   -9.699083117759111e-13
+   -1.392866802449362e-12
+   -2.139278612698071e-11
+     8.31102134048073e-11
+ 3.01e+10    
+    8.298116692224997e-11
+   -2.134914692052396e-11
+    8.507260868890923e-11
+   -1.404314342751842e-12
+   -1.018630006538228e-11
+    8.503020078848903e-11
+   -9.720261258949723e-13
+   -1.396214947410195e-12
+   -2.139508389643191e-11
+    8.310712473863794e-11
+ 3.02e+10    
+     8.29781443276771e-11
+   -2.135151461512377e-11
+     8.50726400848347e-11
+   -1.407673391944537e-12
+    -1.01882139736331e-11
+    8.503018045704684e-11
+    -9.74122917628958e-13
+   -1.399559579720028e-12
+   -2.139739514432659e-11
+    8.310402584480962e-11
+ 3.03e+10    
+    8.297511170831943e-11
+   -2.135389601333125e-11
+    8.507267584803353e-11
+   -1.411028851559803e-12
+   -1.019013858110312e-11
+    8.503016426508116e-11
+   -9.761986491478584e-13
+   -1.402900633740373e-12
+   -2.139971986559708e-11
+    8.310091654698962e-11
+ 3.04e+10    
+    8.297206889231923e-11
+   -2.135629111060564e-11
+    8.507271583996497e-11
+   -1.414380655646024e-12
+   -1.019207388868403e-11
+    8.503015207514808e-11
+   -9.782532830118766e-13
+   -1.406238043877072e-12
+   -2.140205805543975e-11
+    8.309779667150217e-11
+ 3.05e+10    
+    8.296901571041576e-11
+   -2.135869990264079e-11
+    8.507275992376172e-11
+    -1.41772873829124e-12
+    -1.01940198972412e-11
+    8.503014375151477e-11
+   -9.802867821617275e-13
+   -1.409571744579384e-12
+   -2.140440970929898e-11
+    8.309466604729793e-11
+ 3.06e+10    
+    8.296595199591366e-11
+   -2.136112238534984e-11
+    8.507280796420469e-11
+   -1.421073033622321e-12
+   -1.019597660761337e-11
+    8.503013916013207e-11
+   -9.822991099092851e-13
+   -1.412901670339154e-12
+   -2.140677482285147e-11
+    8.309152450592307e-11
+ 3.07e+10    
+    8.296287758464977e-11
+   -2.136355855484917e-11
+    8.507285982769706e-11
+   -1.424413475804261e-12
+   -1.019794402061246e-11
+    8.503013816860696e-11
+    -9.84290229928521e-13
+   -1.416227755690004e-12
+   -2.140915339199016e-11
+      8.3088371881487e-11
+ 3.08e+10    
+    8.295979231495973e-11
+   -2.136600840744261e-11
+    8.507291538223793e-11
+   -1.427749999039531e-12
+   -1.019992213702314e-11
+    8.503014064617586e-11
+   -9.862601062467898e-13
+    -1.41954993520662e-12
+   -2.141154541280856e-11
+    8.308520801062999e-11
+ 3.09e+10    
+    8.295669602764382e-11
+   -2.136847193960567e-11
+    8.507297449739759e-11
+   -1.431082537567407e-12
+    -1.02019109576026e-11
+    8.503014646367711e-11
+   -9.882087032364329e-13
+   -1.422868143504051e-12
+   -2.141395088158457e-11
+    8.308203273249046e-11
+ 3.1e+10     
+    8.295358856593297e-11
+   -2.137094914796992e-11
+    8.507303704429171e-11
+   -1.434411025663468e-12
+   -1.020391048308027e-11
+    8.503015549352431e-11
+    -9.90135985606653e-13
+   -1.426182315237122e-12
+   -2.141636979476456e-11
+    8.307884588867018e-11
+ 3.11e+10    
+    8.295046977545352e-11
+   -2.137344002930678e-11
+    8.507310289555542e-11
+    -1.43773539763908e-12
+   -1.020592071415739e-11
+    8.503016760967935e-11
+   -9.920419183957502e-13
+   -1.429492385099824e-12
+   -2.141880214894746e-11
+    8.307564732320102e-11
+ 3.12e+10    
+    8.294733950419223e-11
+   -2.137594458051219e-11
+    8.507317192531877e-11
+   -1.441055587840927e-12
+    -1.02079416515068e-11
+    8.503018268762583e-11
+   -9.939264669636279e-13
+   -1.432798287824803e-12
+   -2.142124794086862e-11
+    8.307243688250956e-11
+ 3.13e+10    
+    8.294419760246053e-11
+   -2.137846279859061e-11
+    8.507324400918109e-11
+   -1.444371530650611e-12
+   -1.020997329577251e-11
+    8.503020060434286e-11
+   -9.957895969846091e-13
+   -1.436099958182895e-12
+   -2.142370716738417e-11
+    8.306921441538254e-11
+ 3.14e+10    
+    8.294104392285911e-11
+   -2.138099468063943e-11
+    8.507331902418664e-11
+   -1.447683160484317e-12
+   -1.021201564756947e-11
+    8.503022123827837e-11
+   -9.976312744405397e-13
+   -1.439397330982707e-12
+   -2.142617982545487e-11
+    8.306597977293109e-11
+ 3.15e+10    
+    8.293787832024113e-11
+   -2.138354022383325e-11
+    8.507339684879887e-11
+    -1.45099041179249e-12
+   -1.021406870748314e-11
+    8.503024446932344e-11
+   -9.994514656141985e-13
+   -1.442690341070228e-12
+   -2.142866591213032e-11
+    8.306273280855527e-11
+ 3.16e+10    
+    8.293470065167712e-11
+   -2.138609942540862e-11
+    8.507347736287705e-11
+   -1.454293219059599e-12
+   -1.021613247606922e-11
+     8.50302701787862e-11
+   -1.001250137082986e-12
+    -1.44597892332851e-12
+   -2.143116542453334e-11
+    8.305947337790791e-11
+ 3.17e+10    
+    8.293151077641758e-11
+   -2.138867228264819e-11
+    8.507356044765047e-11
+   -1.457591516803898e-12
+   -1.021820695385328e-11
+    8.503029824936619e-11
+   -1.003027255712901e-12
+   -1.449263012677373e-12
+   -2.143367835984415e-11
+    8.305620133885886e-11
+ 3.18e+10    
+     8.29283085558571e-11
+   -2.139125879286555e-11
+    8.507364598569541e-11
+   -1.460885239577296e-12
+   -1.022029214133042e-11
+    8.503032856512919e-11
+   -1.004782788652782e-12
+   -1.452542544073189e-12
+   -2.143620471528473e-11
+    8.305291655145801e-11
+ 3.19e+10    
+    8.292509385349814e-11
+   -2.139385895339002e-11
+    8.507373386090997e-11
+    -1.46417432196521e-12
+   -1.022238803896496e-11
+    8.503036101148134e-11
+   -1.006516703328877e-12
+   -1.455817452508651e-12
+   -2.143874448810343e-11
+    8.304961887789977e-11
+ 3.2e+10     
+    8.292186653491374e-11
+   -2.139647276155139e-11
+    8.507382395849149e-11
+   -1.467458698586477e-12
+   -1.022449464719013e-11
+    8.503039547514518e-11
+   -1.008228967439605e-12
+   -1.459087673012645e-12
+   -2.144129767555946e-11
+    8.304630818248593e-11
+ 3.21e+10    
+    8.291862646771186e-11
+   -2.139910021466483e-11
+    8.507391616491139e-11
+   -1.470738304093369e-12
+   -1.022661196640761e-11
+    8.503043184413367e-11
+   -1.009919548950663e-12
+   -1.462353140650139e-12
+   -2.144386427490761e-11
+    8.304298433158951e-11
+ 3.22e+10    
+    8.291537352149835e-11
+   -2.140174131001617e-11
+    8.507401036789323e-11
+   -1.474013073171543e-12
+   -1.022873999698741e-11
+    8.503047000772686e-11
+   -1.011588416090351e-12
+   -1.465613790522087e-12
+   -2.144644428338323e-11
+    8.303964719361823e-11
+ 3.23e+10    
+    8.291210756784102e-11
+   -2.140439604484693e-11
+    8.507410645638841e-11
+   -1.477282940540096e-12
+   -1.023087873926734e-11
+    8.503050985644673e-11
+   -1.013235537345188e-12
+   -1.468869557765421e-12
+   -2.144903769818691e-11
+    8.303629663897796e-11
+ 3.24e+10    
+    8.290882848023348e-11
+   -2.140706441633988e-11
+    8.507420432055383e-11
+   -1.480547840951676e-12
+   -1.023302819355285e-11
+    8.503055128203367e-11
+   -1.014860881455772e-12
+   -1.472120377553039e-12
+   -2.145164451646989e-11
+    8.303293254003653e-11
+ 3.25e+10    
+     8.29055361340587e-11
+   -2.140974642160436e-11
+    8.507430385172861e-11
+   -1.483807709192585e-12
+   -1.023518836011657e-11
+    8.503059417742243e-11
+    -1.01646441741289e-12
+   -1.475366185093862e-12
+   -2.145426473531908e-11
+     8.30295547710874e-11
+ 3.26e+10    
+    8.290223040655351e-11
+   -2.141244205766219e-11
+    8.507440494241214e-11
+   -1.487062480082926e-12
+   -1.023735923919816e-11
+    8.503063843671914e-11
+   -1.018046114453889e-12
+   -1.478606915632894e-12
+   -2.145689835174265e-11
+    8.302616320831335e-11
+ 3.27e+10    
+    8.289891117677257e-11
+   -2.141515132143321e-11
+    8.507450748624126e-11
+    -1.49031208847682e-12
+   -1.023954083100389e-11
+    8.503068395517733e-11
+   -1.019605942059305e-12
+   -1.481842504451336e-12
+   -2.145954536265541e-11
+     8.30227577297509e-11
+ 3.28e+10    
+    8.289557832555325e-11
+   -2.141787420972161e-11
+    8.507461137796864e-11
+   -1.493556469262627e-12
+   -1.024173313570632e-11
+    8.503073062917567e-11
+   -1.021143869949707e-12
+   -1.485072886866765e-12
+    -2.14622057648647e-11
+     8.30193382152541e-11
+ 3.29e+10    
+    8.289223173548012e-11
+   -2.142061071920191e-11
+    8.507471651344086e-11
+   -1.496795557363184e-12
+   -1.024393615344418e-11
+    8.503077835619501e-11
+   -1.022659868082811e-12
+   -1.488297998233293e-12
+   -2.146487955505625e-11
+    8.301590454645965e-11
+ 3.3e+10     
+    8.288887129085023e-11
+   -2.142336084640539e-11
+    8.507482278957666e-11
+    -1.50002928773615e-12
+   -1.024614988432183e-11
+    8.503082703479565e-11
+     -1.0241539066508e-12
+   -1.491517773941777e-12
+   -2.146756672978014e-11
+    8.301245660675058e-11
+ 3.31e+10    
+    8.288549687763842e-11
+   -2.142612458770659e-11
+    8.507493010434587e-11
+     -1.5032575953743e-12
+    -1.02483743284092e-11
+    8.503087656459576e-11
+   -1.025625956077922e-12
+   -1.494732149420071e-12
+   -2.147026728543729e-11
+    8.300899428122209e-11
+ 3.32e+10    
+    8.288210838346275e-11
+   -2.142890193931006e-11
+    8.507503835674858e-11
+   -1.506480415305875e-12
+   -1.025060948574143e-11
+    8.503092684624942e-11
+    -1.02707598701827e-12
+   -1.497941060133315e-12
+    -2.14729812182657e-11
+    8.300551745664637e-11
+ 3.33e+10    
+    8.287870569755081e-11
+   -2.143169289723737e-11
+    8.507514744679384e-11
+   -1.509697682595027e-12
+   -1.025285535631856e-11
+    8.503097778142459e-11
+   -1.028503970353813e-12
+   -1.501144441584237e-12
+   -2.147570852432721e-11
+    8.300202602143832e-11
+ 3.34e+10    
+    8.287528871070575e-11
+   -2.143449745731406e-11
+    8.507525727547944e-11
+   -1.512909332342169e-12
+   -1.025511194010534e-11
+    8.503102927278242e-11
+    -1.02990987719266e-12
+   -1.504342229313492e-12
+   -2.147844919949434e-11
+    8.299851986562126e-11
+ 3.35e+10    
+     8.28718573152734e-11
+   -2.143731561515711e-11
+    8.507536774477193e-11
+   -1.516115299684491e-12
+   -1.025737923703099e-11
+    8.503108122395607e-11
+   -1.031293678867505e-12
+   -1.507534358900018e-12
+   -2.148120323943726e-11
+    8.299499888079283e-11
+ 3.36e+10    
+    8.286841140510841e-11
+   -2.144014736616226e-11
+    8.507547875758606e-11
+   -1.519315519796372e-12
+   -1.025965724698888e-11
+    8.503113353952958e-11
+   -1.032655346934347e-12
+   -1.510720765961446e-12
+   -2.148397063961105e-11
+    8.299146296009235e-11
+ 3.37e+10    
+    8.286495087554272e-11
+   -2.144299270549197e-11
+    8.507559021776543e-11
+   -1.522509927889937e-12
+   -1.026194596983637e-11
+    8.503118612501823e-11
+   -1.033994853171355e-12
+   -1.513901386154507e-12
+   -2.148675139524323e-11
+    8.298791199816693e-11
+ 3.38e+10    
+    8.286147562335279e-11
+   -2.144585162806322e-11
+    8.507570203006314e-11
+   -1.525698459215572e-12
+   -1.026424540539454e-11
+    8.503123888684757e-11
+   -1.035312169577988e-12
+   -1.517076155175516e-12
+    -2.14895455013212e-11
+    8.298434589113898e-11
+ 3.39e+10    
+    8.285798554672813e-11
+    -2.14487241285356e-11
+    8.507581410012206e-11
+    -1.52888104906246e-12
+     -1.0266555553448e-11
+    8.503129173233442e-11
+   -1.036607268374323e-12
+   -1.520245008760782e-12
+   -2.149235295258041e-11
+    8.298076453657411e-11
+ 3.4e+10     
+    8.285448054523943e-11
+   -2.145161020129972e-11
+    8.507592633445658e-11
+   -1.532057632759193e-12
+   -1.026887641374463e-11
+     8.50313445696664e-11
+   -1.037880122000539e-12
+   -1.523407882687166e-12
+   -2.149517374349207e-11
+    8.297716783344867e-11
+ 3.41e+10    
+    8.285096051980825e-11
+   -2.145450984046575e-11
+    8.507603864043349e-11
+   -1.535228145674361e-12
+   -1.027120798599546e-11
+     8.50313973078836e-11
+   -1.039130703116664e-12
+   -1.526564712772578e-12
+   -2.149800786825178e-11
+    8.297355568211896e-11
+ 3.42e+10    
+    8.284742537267605e-11
+   -2.145742303985213e-11
+    8.507615092625362e-11
+   -1.538392523217165e-12
+   -1.027355026987439e-11
+    8.503144985685893e-11
+   -1.040358984602467e-12
+   -1.529715434876507e-12
+   -2.150085532076786e-11
+    8.296992798428961e-11
+ 3.43e+10    
+    8.284387500737445e-11
+   -2.146034979297467e-11
+    8.507626310093408e-11
+   -1.541550700838118e-12
+   -1.027590326501801e-11
+    8.503150212727945e-11
+   -1.041564939557555e-12
+    -1.53285998490064e-12
+   -2.150371609464997e-11
+     8.29662846429831e-11
+ 3.44e+10    
+    8.284030932869535e-11
+    -2.14632900930357e-11
+    8.507637507429016e-11
+   -1.544702614029644e-12
+   -1.027826697102554e-11
+    8.503155403062852e-11
+   -1.042748541301677e-12
+   -1.535998298789406e-12
+   -2.150659018319834e-11
+    8.296262556250945e-11
+ 3.45e+10    
+    8.283672824266172e-11
+   -2.146624393291336e-11
+    8.507648675691751e-11
+   -1.547848198326841e-12
+   -1.028064138745848e-11
+    8.503160547916704e-11
+   -1.043909763375196e-12
+   -1.539130312530593e-12
+   -2.150947757939259e-11
+    8.295895064843632e-11
+ 3.46e+10    
+    8.283313165649945e-11
+   -2.146921130515141e-11
+    8.507659806017516e-11
+    -1.55098738930817e-12
+   -1.028302651384055e-11
+    8.503165638591614e-11
+   -1.045048579539748e-12
+   -1.542255962156004e-12
+   -2.151237827588142e-11
+    8.295525980756017e-11
+ 3.47e+10    
+    8.282951947860819e-11
+   -2.147219220194902e-11
+    8.507670889616842e-11
+   -1.554120122596168e-12
+   -1.028542234965757e-11
+    8.503170666463951e-11
+   -1.046164963779072e-12
+   -1.545375183742088e-12
+   -2.151529226497203e-11
+    8.295155294787682e-11
+ 3.48e+10    
+    8.282589161853416e-11
+   -2.147518661515072e-11
+    8.507681917773211e-11
+   -1.557246333858223e-12
+   -1.028782889435715e-11
+    8.503175622982528e-11
+    -1.04725889030004e-12
+   -1.548487913410638e-12
+   -2.151821953861987e-11
+    8.294782997855317e-11
+ 3.49e+10    
+    8.282224798694277e-11
+    -2.14781945362369e-11
+    8.507692881841397e-11
+   -1.560365958807348e-12
+    -1.02902461473488e-11
+    8.503180499667093e-11
+   -1.048330333533825e-12
+   -1.551594087329435e-12
+   -2.152116008841899e-11
+    8.294409080989956e-11
+ 3.5e+10     
+    8.281858849559159e-11
+   -2.148121595631412e-11
+    8.507703773245835e-11
+   -1.563478933202956e-12
+   -1.029267410800353e-11
+    8.503185288106457e-11
+   -1.049379268137274e-12
+   -1.554693641713009e-12
+    -2.15241139055919e-11
+    8.294033535334173e-11
+ 3.51e+10    
+    8.281491305730366e-11
+   -2.148425086610596e-11
+    8.507714583479034e-11
+   -1.566585192851678e-12
+   -1.029511277565393e-11
+    8.503189979956994e-11
+   -1.050405668994413e-12
+   -1.557786512823335e-12
+   -2.152708098098041e-11
+    8.293656352139427e-11
+ 3.52e+10    
+    8.281122158594237e-11
+   -2.148729925594377e-11
+    8.507725304099977e-11
+   -1.569684673608187e-12
+    -1.02975621495939e-11
+    8.503194566940963e-11
+   -1.051409511218149e-12
+   -1.560872636970574e-12
+   -2.153006130503614e-11
+    8.293277522763391e-11
+ 3.53e+10    
+    8.280751399638505e-11
+   -2.149036111575811e-11
+    8.507735926732633e-11
+   -1.572777311376006e-12
+   -1.030002222907867e-11
+    8.503199040844922e-11
+   -1.052390770152102e-12
+    -1.56395195051386e-12
+   -2.153305486781152e-11
+    8.292897038667326e-11
+ 3.54e+10    
+    8.280379020449872e-11
+   -2.149343643506984e-11
+    8.507746443064377e-11
+   -1.575863042108422e-12
+   -1.030249301332458e-11
+    8.503203393518218e-11
+    -1.05334942137261e-12
+    -1.56702438986203e-12
+   -2.153606165895085e-11
+    8.292514891413526e-11
+ 3.55e+10    
+    8.280005012711508e-11
+   -2.149652520298196e-11
+    8.507756844844535e-11
+   -1.578941801809285e-12
+   -1.030497450150908e-11
+     8.50320761687139e-11
+   -1.054285440690889e-12
+   -1.570089891474464e-12
+   -2.153908166768184e-11
+    8.292131072662808e-11
+ 3.56e+10    
+    8.279629368200636e-11
+   -2.149962740817112e-11
+    8.507767123882877e-11
+   -1.582013526533935e-12
+   -1.030746669277054e-11
+    8.503211702874695e-11
+   -1.055198804155336e-12
+   -1.573148391861855e-12
+   -2.154211488280701e-11
+    8.291745574172062e-11
+ 3.57e+10    
+     8.27925207878622e-11
+   -2.150274303887984e-11
+    8.507777272048187e-11
+   -1.585078152390098e-12
+   -1.030996958620827e-11
+    8.503215643556677e-11
+   -1.056089488053979e-12
+   -1.576199827587027e-12
+    -2.15451612926956e-11
+    8.291358387791777e-11
+ 3.58e+10    
+    8.278873136426616e-11
+   -2.150587208290873e-11
+    8.507787281266881e-11
+   -1.588135615538766e-12
+   -1.031248318088232e-11
+    8.503219431002621e-11
+   -1.056957468917084e-12
+    -1.57924413526579e-12
+   -2.154822088527563e-11
+    8.290969505463739e-11
+ 3.59e+10    
+    8.278492533167305e-11
+   -2.150901452760883e-11
+    8.507797143521551e-11
+   -1.591185852195138e-12
+   -1.031500747581353e-11
+    8.503223057353219e-11
+   -1.057802723519885e-12
+   -1.582281251567773e-12
+     -2.1551293648026e-11
+     8.29057891921861e-11
+ 3.6e+10     
+    8.278110261138652e-11
+   -2.151217035987429e-11
+     8.50780685084965e-11
+   -1.594228798629559e-12
+   -1.031754246998337e-11
+    8.503226514803121e-11
+   -1.058625228885465e-12
+   -1.585311113217285e-12
+   -2.155437956796911e-11
+    8.290186621173743e-11
+ 3.61e+10    
+    8.277726312553802e-11
+   -2.151533956613528e-11
+    8.507816395342112e-11
+   -1.597264391168445e-12
+   -1.032008816233392e-11
+     8.50322979559957e-11
+    -1.05942496228778e-12
+   -1.588333656994162e-12
+   -2.155747863166334e-11
+    8.289792603530869e-11
+ 3.62e+10    
+    8.277340679706425e-11
+   -2.151852213235097e-11
+    8.507825769142049e-11
+   -1.600292566195254e-12
+   -1.032264455176779e-11
+    8.503232892041086e-11
+   -1.060201901254786e-12
+   -1.591348819734692e-12
+   -2.156059082519613e-11
+    8.289396858573953e-11
+ 3.63e+10    
+    8.276953354968764e-11
+   -2.152171804400293e-11
+    8.507834964443438e-11
+   -1.603313260151443e-12
+   -1.032521163714811e-11
+    8.503235796476112e-11
+   -1.060956023571737e-12
+   -1.594356538332449e-12
+     -2.1563716134177e-11
+    8.288999378667032e-11
+ 3.64e+10    
+    8.276564330789467e-11
+   -2.152492728608838e-11
+    8.507843973489894e-11
+   -1.606326409537449e-12
+   -1.032778941729841e-11
+    8.503238501301716e-11
+   -1.061687307284562e-12
+   -1.597356749739262e-12
+   -2.156685454373068e-11
+    8.288600156252113e-11
+ 3.65e+10    
+    8.276173599691663e-11
+    -2.15281498431141e-11
+     8.50785278857335e-11
+   -1.609331950913669e-12
+   -1.033037789100265e-11
+    8.503240998962366e-11
+   -1.062395730703419e-12
+   -1.600349390966064e-12
+   -2.157000603849088e-11
+    8.288199183847108e-11
+ 3.66e+10    
+       8.275781154271e-11
+   -2.153138569909018e-11
+    8.507861402032903e-11
+   -1.612329820901461e-12
+   -1.033297705700512e-11
+    8.503243281948638e-11
+   -1.063081272406316e-12
+   -1.603334399083862e-12
+   -2.157317060259385e-11
+    8.287796454043843e-11
+ 3.67e+10    
+     8.27538698719372e-11
+   -2.153463483752415e-11
+     8.50786980625357e-11
+   -1.615319956184134e-12
+   -1.033558691401046e-11
+     8.50324534279599e-11
+   -1.063743911242905e-12
+   -1.606311711224635e-12
+   -2.157634821967229e-11
+    8.287391959506094e-11
+ 3.68e+10    
+    8.274991091194734e-11
+   -2.153789724141509e-11
+     8.50787799366512e-11
+   -1.618302293507972e-12
+   -1.033820746068358e-11
+    8.503247174083628e-11
+   -1.064383626338331e-12
+   -1.609281264582307e-12
+   -2.157953887284961e-11
+    8.286985692967641e-11
+ 3.69e+10    
+    8.274593459075907e-11
+   -2.154117289324848e-11
+    8.507885956740945e-11
+   -1.621276769683234e-12
+   -1.034083869564971e-11
+    8.503248768433261e-11
+   -1.065000397097253e-12
+   -1.612242996413657e-12
+   -2.158274254473403e-11
+    8.286577647230397e-11
+ 3.7e+10     
+    8.274194083704186e-11
+   -2.154446177499046e-11
+    8.507893687996863e-11
+   -1.624243321585219e-12
+   -1.034348061749425e-11
+       8.503250118508e-11
+    -1.06559420320793e-12
+   -1.615196844039298e-12
+   -2.158595921741335e-11
+    8.286167815162594e-11
+ 3.71e+10    
+     8.27379295800986e-11
+   -2.154776386808285e-11
+    8.507901179990089e-11
+    -1.62720188615524e-12
+   -1.034613322476285e-11
+    8.503251217011197e-11
+    -1.06616502464643e-12
+   -1.618142744844652e-12
+   -2.158918887244936e-11
+    8.285756189696925e-11
+ 3.72e+10    
+    8.273390074984906e-11
+    -2.15510791534383e-11
+    8.507908425318093e-11
+   -1.630152400401718e-12
+   -1.034879651596139e-11
+    8.503252056685376e-11
+   -1.066712841680958e-12
+   -1.621080636280895e-12
+    -2.15924314908731e-11
+     8.28534276382887e-11
+ 3.73e+10    
+    8.272985427681263e-11
+   -2.155440761143531e-11
+    8.507915416617546e-11
+   -1.633094801401181e-12
+   -1.035147048955592e-11
+    8.503252630311126e-11
+   -1.067237634876257e-12
+   -1.624010455865942e-12
+   -2.159568705317966e-11
+    8.284927530614917e-11
+ 3.74e+10    
+    8.272579009209238e-11
+   -2.155774922191382e-11
+    8.507922146563269e-11
+   -1.636029026299352e-12
+   -1.035415514397263e-11
+    8.503252930706054e-11
+    -1.06773938509813e-12
+   -1.626932141185454e-12
+   -2.159895553932369e-11
+     8.28451048317093e-11
+ 3.75e+10    
+    8.272170812735928e-11
+   -2.156110396417079e-11
+    8.507928607867229e-11
+   -1.638955012312175e-12
+   -1.035685047759794e-11
+    8.503252950723762e-11
+   -1.068218073518044e-12
+   -1.629845629893787e-12
+   -2.160223692871472e-11
+    8.284091614670481e-11
+ 3.76e+10    
+    8.271760831483643e-11
+   -2.156447181695589e-11
+    8.507934793277528e-11
+   -1.641872696726912e-12
+    -1.03595564887784e-11
+    8.503252683252805e-11
+   -1.068673681617834e-12
+    -1.63275085971504e-12
+   -2.160553120021297e-11
+    8.283670918343316e-11
+ 3.77e+10    
+    8.271349058728437e-11
+   -2.156785275846759e-11
+    8.507940695577413e-11
+   -1.644782016903147e-12
+   -1.036227317582068e-11
+     8.50325212121571e-11
+   -1.069106191194506e-12
+   -1.635647768444009e-12
+   -2.160883833212498e-11
+    8.283248387473718e-11
+ 3.78e+10    
+    8.270935487798585e-11
+   -2.157124676634917e-11
+    8.507946307584335e-11
+   -1.647682910273938e-12
+   -1.036500053699166e-11
+    8.503251257568041e-11
+   -1.069515584365098e-12
+   -1.638536293947214e-12
+   -2.161215830220006e-11
+    8.282824015399071e-11
+ 3.79e+10    
+     8.27052011207318e-11
+   -2.157465381768522e-11
+    8.507951622148969e-11
+   -1.650575314346825e-12
+   -1.036773857051825e-11
+    8.503250085297363e-11
+   -1.069901843571667e-12
+   -1.641416374163934e-12
+   -2.161549108762595e-11
+    8.282397795508319e-11
+ 3.8e+10     
+    8.270102924980747e-11
+   -2.157807388899798e-11
+    8.507956632154343e-11
+   -1.653459166704932e-12
+   -1.037048727458762e-11
+     8.50324859742245e-11
+   -1.070264951586332e-12
+   -1.644287947107165e-12
+   -2.161883666502575e-11
+    8.281969721240565e-11
+ 3.81e+10    
+     8.26968391999784e-11
+   -2.158150695624404e-11
+    8.507961330514896e-11
+   -1.656334405008062e-12
+   -1.037324664734702e-11
+    8.503246786992226e-11
+   -1.070604891516398e-12
+   -1.647150950864703e-12
+   -2.162219501045411e-11
+    8.281539786083663e-11
+ 3.82e+10    
+    8.269263090647737e-11
+   -2.158495299481132e-11
+    8.507965710175648e-11
+    -1.65920096699374e-12
+   -1.037601668690382e-11
+    8.503244647084987e-11
+   -1.070921646809574e-12
+    -1.65000532360014e-12
+   -2.162556609939417e-11
+    8.281107983572819e-11
+ 3.83e+10    
+    8.268840430499154e-11
+   -2.158841197951577e-11
+    8.507969764111253e-11
+    -1.66205879047836e-12
+   -1.037879739132553e-11
+    8.503242170807471e-11
+   -1.071215201259254e-12
+   -1.652851003553876e-12
+   -2.162894990675443e-11
+    8.280674307289322e-11
+ 3.84e+10    
+     8.26841593316496e-11
+   -2.159188388459886e-11
+    8.507973485325255e-11
+   -1.664907813358215e-12
+   -1.038158875863981e-11
+    8.503239351294052e-11
+   -1.071485539009851e-12
+   -1.655687929044193e-12
+   -2.163234640686569e-11
+    8.280238750859145e-11
+ 3.85e+10    
+    8.267989592300954e-11
+   -2.159536868372469e-11
+    8.507976866849197e-11
+   -1.667747973610631e-12
+   -1.038439078683441e-11
+    8.503236181705881e-11
+   -1.071732644562256e-12
+   -1.658516038468259e-12
+    -2.16357555734786e-11
+    8.279801307951796e-11
+ 3.86e+10    
+    8.267561401604713e-11
+   -2.159886634997763e-11
+    8.507979901741839e-11
+   -1.670579209295036e-12
+   -1.038720347385725e-11
+    8.503232655230082e-11
+   -1.071956502779318e-12
+   -1.661335270303144e-12
+    -2.16391773797608e-11
+    8.279361972278995e-11
+ 3.87e+10    
+    8.267131354814356e-11
+   -2.160237685585981e-11
+    8.507982583088355e-11
+    -1.67340145855409e-12
+    -1.03900268176163e-11
+    8.503228765078975e-11
+   -1.072157098891379e-12
+    -1.66414556310694e-12
+   -2.164261179829463e-11
+    8.278920737593544e-11
+ 3.88e+10    
+    8.266699445707509e-11
+   -2.160590017328916e-11
+    8.507984903999601e-11
+   -1.676214659614734e-12
+   -1.039286081597972e-11
+    8.503224504489295e-11
+   -1.072334418501939e-12
+   -1.666946855519721e-12
+   -2.164605880107486e-11
+    8.278477597688127e-11
+ 3.89e+10    
+    8.266265668100093e-11
+   -2.160943627359709e-11
+    8.507986857611305e-11
+   -1.679018750789339e-12
+   -1.039570546677578e-11
+    8.503219866721459e-11
+   -1.072488447593289e-12
+   -1.669739086264629e-12
+   -2.164951835950658e-11
+    8.278032546394183e-11
+ 3.9e+10     
+    8.265830015845356e-11
+   -2.161298512752686e-11
+    8.507988437083403e-11
+   -1.681813670476772e-12
+   -1.039856076779279e-11
+    8.503214845058759e-11
+   -1.072619172532299e-12
+   -1.672522194148923e-12
+   -2.165299044440319e-11
+    8.277585577580816e-11
+ 3.91e+10    
+    8.265392482832787e-11
+   -2.161654670523164e-11
+    8.507989635599246e-11
+   -1.684599357163514e-12
+   -1.040142671677921e-11
+    8.503209432806719e-11
+    -1.07272658007617e-12
+   -1.675296118065013e-12
+   -2.165647502598464e-11
+    8.277136685153706e-11
+ 3.92e+10    
+      8.2649530629871e-11
+   -2.162012097627311e-11
+    8.507990446364979e-11
+   -1.687375749424766e-12
+    -1.04043033114436e-11
+    8.503203623292401e-11
+     -1.0728106573783e-12
+   -1.678060796991508e-12
+   -2.165997207387599e-11
+    8.276685863054119e-11
+ 3.93e+10    
+    8.264511750267271e-11
+   -2.162370790961976e-11
+    8.507990862608774e-11
+   -1.690142785925526e-12
+   -1.040719054945455e-11
+    8.503197409863637e-11
+   -1.072871391994193e-12
+     -1.6808161699943e-12
+   -2.166348155710546e-11
+    8.276233105257806e-11
+ 3.94e+10    
+    8.264068538665605e-11
+   -2.162730747364599e-11
+    8.507990877580245e-11
+    -1.69290040542174e-12
+   -1.041008842844073e-11
+    8.503190785888427e-11
+   -1.072908771887382e-12
+   -1.683562176227599e-12
+   -2.166700344410353e-11
+    8.275778405774121e-11
+ 3.95e+10    
+    8.263623422206745e-11
+   -2.163091963613048e-11
+    8.507990484549735e-11
+   -1.695648546761367e-12
+    -1.04129969459909e-11
+    8.503183744754312e-11
+   -1.072922785435437e-12
+   -1.686298754934962e-12
+   -2.167053770270154e-11
+    8.275321758645014e-11
+ 3.96e+10    
+    8.263176394946862e-11
+   -2.163454436425554e-11
+      8.5079896768077e-11
+   -1.698387148885505e-12
+   -1.041591609965379e-11
+     8.50317627986766e-11
+   -1.072913421436004e-12
+   -1.689025845450386e-12
+   -2.167408430013064e-11
+    8.274863157944108e-11
+ 3.97e+10    
+    8.262727450972716e-11
+   -2.163818162460606e-11
+    8.507988447664117e-11
+   -1.701116150829466e-12
+   -1.041884588693814e-11
+    8.503168384653117e-11
+   -1.072880669112874e-12
+   -1.691743387199381e-12
+   -2.167764320302091e-11
+    8.274402597775838e-11
+ 3.98e+10    
+    8.262276584400843e-11
+   -2.164183138316877e-11
+    8.507986790447857e-11
+   -1.703835491723924e-12
+   -1.042178630531274e-11
+    8.503160052552975e-11
+   -1.072824518122103e-12
+   -1.694451319699962e-12
+   -2.168121437740052e-11
+    8.273940072274533e-11
+ 3.99e+10    
+    8.261823789376717e-11
+   -2.164549360533171e-11
+    8.507984698506072e-11
+   -1.706545110795995e-12
+   -1.042473735220627e-11
+    8.503151277026587e-11
+   -1.072744958558173e-12
+   -1.697149582563769e-12
+   -2.168479778869517e-11
+    8.273475575603611e-11
+ 4e+10       
+    8.261369060073994e-11
+    -2.16491682558836e-11
+    8.507982165203663e-11
+   -1.709244947370351e-12
+   -1.042769902500735e-11
+    8.503142051549814e-11
+    -1.07264198096017e-12
+   -1.699838115497102e-12
+   -2.168839340172754e-11
+    8.273009101954756e-11
+ 4.01e+10    
+    8.260912390693707e-11
+   -2.165285529901376e-11
+    8.507979183922728e-11
+   -1.711934940870277e-12
+   -1.043067132106452e-11
+    8.503132369614443e-11
+   -1.072515576318021e-12
+   -1.702516858301967e-12
+   -2.169200118071687e-11
+    8.272540645547096e-11
+ 4.02e+10    
+    8.260453775463513e-11
+   -2.165655469831146e-11
+    8.507975748061944e-11
+    -1.71461503081887e-12
+    -1.04336542376861e-11
+    8.503122224727672e-11
+   -1.072365736078727e-12
+   -1.705185750877175e-12
+    -2.16956210892788e-11
+    8.272070200626472e-11
+ 4.03e+10    
+    8.259993208637017e-11
+   -2.166026641676629e-11
+    8.507971851036144e-11
+   -1.717285156840047e-12
+   -1.043664777214031e-11
+    8.503111610411552e-11
+   -1.072192452152667e-12
+    -1.70784473321937e-12
+   -2.169925309042517e-11
+     8.27159776146469e-11
+ 4.04e+10    
+    8.259530684493025e-11
+   -2.166399041676776e-11
+    8.507967486275705e-11
+   -1.719945258659699e-12
+   -1.043965192165508e-11
+    8.503100520202521e-11
+   -1.071995716919883e-12
+   -1.710493745424089e-12
+   -2.170289714656412e-11
+    8.271123322358785e-11
+ 4.05e+10    
+    8.259066197334895e-11
+   -2.166772666010576e-11
+    8.507962647226109e-11
+   -1.722595276106775e-12
+   -1.044266668341804e-11
+    8.503088947650862e-11
+    -1.07177552323642e-12
+   -1.713132727686835e-12
+   -2.170655321950008e-11
+    8.270646877630334e-11
+ 4.06e+10    
+    8.258599741489873e-11
+   -2.167147510797072e-11
+     8.50795732734743e-11
+   -1.725235149114383e-12
+   -1.044569205457655e-11
+    8.503076886320237e-11
+   -1.071531864440681e-12
+   -1.715761620304146e-12
+   -2.171022127043416e-11
+     8.27016842162478e-11
+ 4.07e+10    
+    8.258131311308491e-11
+   -2.167523572095387e-11
+    8.507951520113866e-11
+   -1.727864817720901e-12
+    -1.04487280322375e-11
+    8.503064329787235e-11
+   -1.071264734359794e-12
+   -1.718380363674621e-12
+   -2.171390125996447e-11
+    8.269687948710804e-11
+ 4.08e+10    
+    8.257660901163868e-11
+   -2.167900845904783e-11
+    8.507945219013255e-11
+   -1.730484222071043e-12
+   -1.045177461346735e-11
+    8.503051271640876e-11
+      -1.070974127316e-12
+   -1.720988898300005e-12
+   -2.171759314808657e-11
+    8.269205453279644e-11
+ 4.09e+10    
+    8.257188505451237e-11
+   -2.168279328164731e-11
+    8.507938417546672e-11
+   -1.733093302416997e-12
+   -1.045483179529204e-11
+    8.503037705482205e-11
+   -1.070660038133065e-12
+   -1.723587164786265e-12
+   -2.172129689419415e-11
+    8.268720929744551e-11
+ 4.1e+10     
+    8.256714118587284e-11
+   -2.168659014754963e-11
+    8.507931109227955e-11
+   -1.735691999119497e-12
+   -1.045789957469688e-11
+    8.503023624923833e-11
+   -1.070322462142696e-12
+    -1.72617510384459e-12
+   -2.172501245707972e-11
+    8.268234372540182e-11
+ 4.11e+10    
+    8.256237735009641e-11
+   -2.169039901495571e-11
+    8.507923287583278e-11
+   -1.738280252648901e-12
+   -1.046097794862651e-11
+    8.503009023589536e-11
+   -1.069961395190965e-12
+   -1.728752656292501e-12
+   -2.172873979493532e-11
+    8.267745776121955e-11
+ 4.12e+10    
+    8.255759349176334e-11
+   -2.169421984147086e-11
+    8.507914946150755e-11
+    -1.74085800358632e-12
+   -1.046406691398481e-11
+     8.50299389511387e-11
+   -1.069576833644758e-12
+   -1.731319763054901e-12
+   -2.173247886535372e-11
+    8.267255134965665e-11
+ 4.13e+10    
+    8.255278955565289e-11
+   -2.169805258410601e-11
+    8.507906078480079e-11
+   -1.743425192624695e-12
+   -1.046716646763479e-11
+    8.502978233141708e-11
+   -1.069168774398209e-12
+   -1.733876365165115e-12
+   -2.173622962532916e-11
+    8.266762443566782e-11
+ 4.14e+10    
+    8.254796548673832e-11
+   -2.170189719927863e-11
+     8.50789667813204e-11
+   -1.745981760569873e-12
+    -1.04702766063985e-11
+    8.502962031327934e-11
+   -1.068737214879167e-12
+    -1.73642240376596e-12
+   -2.173999203125877e-11
+    8.266267696440075e-11
+ 4.15e+10    
+    8.254312123018174e-11
+   -2.170575364281419e-11
+     8.50788673867826e-11
+    -1.74852764834171e-12
+   -1.047339732705699e-11
+    8.502945283337044e-11
+   -1.068282153055631e-12
+   -1.738957820110798e-12
+   -2.174376603894367e-11
+    8.265770888119062e-11
+ 4.16e+10    
+    8.253825673133029e-11
+   -2.170962186994727e-11
+    8.507876253700712e-11
+   -1.751062796975151e-12
+    -1.04765286263501e-11
+    8.502927982842781e-11
+   -1.067803587442228e-12
+   -1.741482555564569e-12
+   -2.174755160359038e-11
+    8.265272013155528e-11
+ 4.17e+10    
+      8.2533371935711e-11
+   -2.171350183532321e-11
+    8.507865216791497e-11
+   -1.753587147621325e-12
+   -1.047967050097642e-11
+    8.502910123527806e-11
+   -1.067301517106665e-12
+   -1.743996551604896e-12
+   -2.175134867981228e-11
+     8.26477106611912e-11
+ 4.18e+10    
+    8.252846678902674e-11
+   -2.171739349299946e-11
+    8.507853621552356e-11
+   -1.756100641548612e-12
+   -1.048282294759317e-11
+     8.50289169908335e-11
+    -1.06677594167616e-12
+   -1.746499749823079e-12
+   -2.175515722163108e-11
+    8.264268041596851e-11
+ 4.19e+10    
+    8.252354123715251e-11
+   -2.172129679644748e-11
+    8.507841461594502e-11
+   -1.758603220143739e-12
+   -1.048598596281606e-11
+    8.502872703208893e-11
+   -1.066226861343926e-12
+   -1.748992091925208e-12
+   -2.175897718247868e-11
+    8.263762934192755e-11
+ 4.2e+10     
+    8.251859522613115e-11
+   -2.172521169855413e-11
+    8.507828730538131e-11
+   -1.761094824912873e-12
+   -1.048915954321909e-11
+    8.502853129611859e-11
+   -1.065654276875584e-12
+   -1.751473519733156e-12
+   -2.176280851519863e-11
+    8.263255738527388e-11
+ 4.21e+10    
+    8.251362870216937e-11
+   -2.172913815162377e-11
+    8.507815422012284e-11
+   -1.763575397482659e-12
+   -1.049234368533462e-11
+    8.502832972007309e-11
+   -1.065058189615614e-12
+   -1.753943975185667e-12
+   -2.176665117204833e-11
+     8.26274644923756e-11
+ 4.22e+10    
+    8.250864161163462e-11
+   -2.173307610737991e-11
+    8.507801529654372e-11
+   -1.766044879601337e-12
+   -1.049553838565296e-11
+    8.502812224117645e-11
+    -1.06443860149377e-12
+   -1.756403400339408e-12
+   -2.177050510470058e-11
+    8.262235060975839e-11
+ 4.23e+10    
+    8.250363390105143e-11
+   -2.173702551696749e-11
+    8.507787047110036e-11
+   -1.768503213139805e-12
+    -1.04987436406224e-11
+    8.502790879672334e-11
+   -1.063795515031504e-12
+       -1.75885173737e-12
+   -2.177437026424588e-11
+    8.261721568410289e-11
+ 4.24e+10    
+     8.24986055170979e-11
+   -2.174098633095472e-11
+    8.507771968032781e-11
+   -1.770950340092683e-12
+   -1.050195944664903e-11
+    8.502768932407626e-11
+   -1.063128933348358e-12
+   -1.761288928573085e-12
+   -2.177824660119439e-11
+    8.261205966224095e-11
+ 4.25e+10    
+    8.249355640660269e-11
+   -2.174495849933524e-11
+    8.507756286083731e-11
+   -1.773386202579412e-12
+   -1.050518580009652e-11
+     8.50274637606632e-11
+   -1.062438860168342e-12
+   -1.763714916365346e-12
+   -2.178213406547817e-11
+    8.260688249115209e-11
+ 4.26e+10    
+    8.248848651654214e-11
+   -2.174894197153066e-11
+    8.507739994931371e-11
+   -1.775810742845296e-12
+   -1.050842269728601e-11
+    8.502723204397484e-11
+   -1.061725299826304e-12
+   -1.766129643285594e-12
+   -2.178603260645356e-11
+    8.260168411796116e-11
+ 4.27e+10    
+    8.248339579403672e-11
+   -2.175293669639244e-11
+    8.507723088251299e-11
+   -1.778223903262598e-12
+   -1.051167013449586e-11
+    8.502699411156216e-11
+    -1.06098825727428e-12
+   -1.768533051995796e-12
+    -2.17899421729033e-11
+    8.259646448993435e-11
+ 4.28e+10    
+    8.247828418634912e-11
+   -2.175694262220464e-11
+    8.507705559725974e-11
+    -1.78062562633158e-12
+   -1.051492810796156e-11
+    8.502674990103433e-11
+   -1.060227738087817e-12
+   -1.770925085282105e-12
+   -2.179386271303929e-11
+    8.259122355447739e-11
+ 4.29e+10    
+    8.247315164088079e-11
+   -2.176095969668627e-11
+     8.50768740304449e-11
+   -1.783015854681593e-12
+   -1.051819661387551e-11
+    8.502649935005607e-11
+    -1.05944374847227e-12
+   -1.773305686055925e-12
+   -2.179779417450471e-11
+     8.25859612591316e-11
+ 4.3e+10     
+    8.246799810517026e-11
+   -2.176498786699388e-11
+    8.507668611902357e-11
+    -1.78539453107215e-12
+   -1.052147564838673e-11
+      8.5026242396346e-11
+    -1.05863629526909e-12
+   -1.775674797354964e-12
+   -2.180173650437708e-11
+    8.258067755157279e-11
+ 4.31e+10    
+    8.246282352688971e-11
+   -2.176902707972409e-11
+    8.507649180001275e-11
+   -1.787761598393962e-12
+   -1.052476520760079e-11
+    8.502597897767424e-11
+   -1.057805385962065e-12
+   -1.778032362344258e-12
+   -2.180568964917056e-11
+    8.257537237960759e-11
+ 4.32e+10    
+    8.245762785384334e-11
+    -2.17730772809164e-11
+     8.50762910104892e-11
+   -1.790116999670009e-12
+   -1.052806528757953e-11
+    8.502570903186046e-11
+   -1.056951028683552e-12
+   -1.780378324317221e-12
+    -2.18096535548389e-11
+    8.257004569117165e-11
+ 4.33e+10    
+    8.245241103396537e-11
+     -2.1777138416056e-11
+    8.507608368758795e-11
+   -1.792460678056626e-12
+   -1.053137588434084e-11
+      8.5025432496772e-11
+   -1.056073232220664e-12
+   -1.782712626696697e-12
+    -2.18136281667781e-11
+    8.256469743432713e-11
+ 4.34e+10    
+    8.244717301531736e-11
+   -2.178121043007649e-11
+    8.507586976849977e-11
+   -1.794792576844545e-12
+   -1.053469699385847e-11
+    8.502514931032242e-11
+   -1.055172006021441e-12
+   -1.785035213035992e-12
+    -2.18176134298296e-11
+    8.255932755726111e-11
+ 4.35e+10    
+    8.244191374608667e-11
+   -2.178529326736289e-11
+    8.507564919046963e-11
+   -1.797112639459939e-12
+   -1.053802861206176e-11
+    8.502485941046908e-11
+   -1.054247360200972e-12
+   -1.787346027019908e-12
+   -2.182160928828279e-11
+    8.255393600828299e-11
+ 4.36e+10    
+    8.243663317458427e-11
+   -2.178938687175443e-11
+    8.507542189079499e-11
+   -1.799420809465514e-12
+   -1.054137073483537e-11
+    8.502456273521205e-11
+   -1.053299305547486e-12
+   -1.789645012465825e-12
+   -2.182561568587852e-11
+    8.254852273582317e-11
+ 4.37e+10    
+    8.243133124924361e-11
+   -2.179349118654801e-11
+    8.507518780682417e-11
+   -1.801717030561541e-12
+   -1.054472335801917e-11
+    8.502425922259256e-11
+   -1.052327853528426e-12
+   -1.791932113324682e-12
+   -2.182963256581185e-11
+    8.254308768843063e-11
+ 4.38e+10    
+    8.242600791861828e-11
+   -2.179760615450086e-11
+    8.507494687595481e-11
+   -1.804001246586921e-12
+   -1.054808647740777e-11
+    8.502394881069093e-11
+   -1.051333016296456e-12
+   -1.794207273682093e-12
+   -2.183365987073532e-11
+    8.253763081477192e-11
+ 4.39e+10    
+     8.24206631313809e-11
+    -2.18017317178339e-11
+    8.507469903563203e-11
+   -1.806273401520244e-12
+   -1.055146008875046e-11
+    8.502363143762585e-11
+   -1.050314806695438e-12
+   -1.796470437759282e-12
+    -2.18376975427623e-11
+    8.253215206362915e-11
+ 4.4e+10     
+    8.241529683632121e-11
+   -2.180586781823501e-11
+     8.50744442233474e-11
+   -1.808533439480809e-12
+   -1.055484418775083e-11
+    8.502330704155256e-11
+    -1.04927323826639e-12
+   -1.798721549914259e-12
+   -2.184174552346998e-11
+    8.252665138389871e-11
+ 4.41e+10    
+    8.240990898234549e-11
+   -2.181001439686227e-11
+    8.507418237663726e-11
+   -1.810781304729748e-12
+    -1.05582387700665e-11
+     8.50229755606618e-11
+   -1.048208325253357e-12
+   -1.800960554642744e-12
+   -2.184580375390305e-11
+    8.252112872458978e-11
+ 4.42e+10    
+    8.240449951847453e-11
+   -2.181417139434733e-11
+    8.507391343308169e-11
+   -1.813016941671018e-12
+   -1.056164383130888e-11
+     8.50226369331788e-11
+   -1.047120082609285e-12
+   -1.803187396579251e-12
+   -2.184987217457698e-11
+    8.251558403482328e-11
+ 4.43e+10    
+     8.23990683938428e-11
+   -2.181833875079873e-11
+    8.507363733030301e-11
+   -1.815240294852469e-12
+    -1.05650593670428e-11
+    8.502229109736146e-11
+   -1.046008526001816e-12
+   -1.805402020498144e-12
+   -2.185395072548129e-11
+    8.251001726383012e-11
+ 4.44e+10    
+    8.239361555769707e-11
+   -2.182251640580547e-11
+    8.507335400596496e-11
+   -1.817451308966893e-12
+   -1.056848537278628e-11
+    8.502193799150004e-11
+   -1.044873671819046e-12
+   -1.807604371314668e-12
+   -2.185803934608336e-11
+    8.250442836095087e-11
+ 4.45e+10    
+    8.238814095939587e-11
+   -2.182670429844051e-11
+    8.507306339777138e-11
+   -1.819649928853086e-12
+   -1.057192184401023e-11
+    8.502157755391587e-11
+   -1.043715537175234e-12
+   -1.809794394085973e-12
+    -2.18621379753319e-11
+    8.249881727563408e-11
+ 4.46e+10    
+    8.238264454840814e-11
+   -2.183090236726424e-11
+     8.50727654434648e-11
+   -1.821836099496897e-12
+   -1.057536877613801e-11
+    8.502120972296017e-11
+   -1.042534139916476e-12
+   -1.811972034012153e-12
+   -2.186624655166049e-11
+    8.249318395743567e-11
+ 4.47e+10    
+     8.23771262743125e-11
+   -2.183511055032827e-11
+    8.507246008082675e-11
+   -1.824009766032232e-12
+    -1.05788261645453e-11
+    8.502083443701358e-11
+   -1.041329498626287e-12
+   -1.814137236437337e-12
+   -2.187036501299138e-11
+    8.248752835601815e-11
+ 4.48e+10    
+    8.237158608679637e-11
+   -2.183932878517879e-11
+    8.507214724767499e-11
+   -1.826170873742208e-12
+   -1.058229400455958e-11
+    8.502045163448525e-11
+   -1.040101632631159e-12
+   -1.816289946850645e-12
+   -2.187449329673918e-11
+    8.248185042114933e-11
+ 4.49e+10    
+    8.236602393565564e-11
+   -2.184355700886079e-11
+    8.507182688186456e-11
+   -1.828319368060063e-12
+   -1.058577229145991e-11
+    8.502006125381185e-11
+   -1.038850562006087e-12
+   -1.818430110887322e-12
+    -2.18786313398146e-11
+    8.247615010270231e-11
+ 4.5e+10     
+    8.236043977079313e-11
+   -2.184779515792124e-11
+    8.507149892128556e-11
+   -1.830455194570327e-12
+   -1.058926102047657e-11
+    8.501966323345728e-11
+    -1.03757630757997e-12
+   -1.820557674329701e-12
+   -2.188277907862839e-11
+    8.247042735065434e-11
+ 4.51e+10    
+    8.235483354221956e-11
+    -2.18520431684134e-11
+    8.507116330386318e-11
+   -1.832578299009795e-12
+   -1.059276018679059e-11
+    8.501925751191146e-11
+   -1.036278890941027e-12
+   -1.822672583108298e-12
+     -2.1886936449095e-11
+    8.246468211508632e-11
+ 4.52e+10    
+     8.23492052000511e-11
+   -2.185630097590027e-11
+    8.507081996755677e-11
+   -1.834688627268606e-12
+   -1.059626978553359e-11
+    8.501884402769059e-11
+   -1.034958334442101e-12
+    -1.82477478330283e-12
+   -2.189110338663684e-11
+    8.245891434618266e-11
+ 4.53e+10    
+    8.234355469451065e-11
+   -2.186056851545888e-11
+    8.507046885035949e-11
+   -1.836786125391281e-12
+   -1.059978981178725e-11
+    8.501842271933596e-11
+   -1.033614661205931e-12
+   -1.826864221143264e-12
+   -2.189527982618787e-11
+    8.245312399423035e-11
+ 4.54e+10    
+    8.233788197592624e-11
+   -2.186484572168384e-11
+    8.507010989029718e-11
+   -1.838870739577782e-12
+   -1.060332026058295e-11
+    8.501799352541356e-11
+   -1.032247895130352e-12
+   -1.828940843010861e-12
+   -2.189946570219794e-11
+    8.244731100961901e-11
+ 4.55e+10    
+    8.233218699473157e-11
+   -2.186913252869166e-11
+    8.506974302542861e-11
+    -1.84094241618452e-12
+   -1.060686112690147e-11
+    8.501755638451392e-11
+   -1.030858060893441e-12
+   -1.831004595439226e-12
+   -2.190366094863663e-11
+    8.244147534284044e-11
+ 4.56e+10    
+    8.232646970146507e-11
+   -2.187342887012446e-11
+    8.506936819384424e-11
+   -1.843001101725485e-12
+   -1.061041240567247e-11
+    8.501711123525168e-11
+   -1.029445183958566e-12
+   -1.833055425115344e-12
+   -2.190786549899729e-11
+    8.243561694448802e-11
+ 4.57e+10    
+    8.232073004677036e-11
+   -2.187773467915443e-11
+    8.506898533366681e-11
+     -1.8450467428732e-12
+   -1.061397409177428e-11
+    8.501665801626524e-11
+   -1.028009290579426e-12
+   -1.835093278880645e-12
+   -2.191207928630147e-11
+    8.242973576525738e-11
+ 4.58e+10    
+    8.231496798139541e-11
+   -2.188204988848741e-11
+    8.506859438304969e-11
+   -1.847079286459846e-12
+   -1.061754618003324e-11
+    8.501619666621635e-11
+    -1.02655040780496e-12
+   -1.837118103732021e-12
+    -2.19163022431028e-11
+     8.24238317559453e-11
+ 4.59e+10    
+    8.230918345619296e-11
+   -2.188637443036757e-11
+    8.506819528017789e-11
+   -1.849098679478256e-12
+   -1.062112866522349e-11
+    8.501572712379019e-11
+   -1.025068563484237e-12
+   -1.839129846822911e-12
+   -2.192053430149131e-11
+    8.241790486745042e-11
+ 4.6e+10     
+    8.230337642212035e-11
+   -2.189070823658113e-11
+    8.506778796326681e-11
+    -1.85110486908301e-12
+   -1.062472154206644e-11
+    8.501524932769526e-11
+   -1.023563786271254e-12
+   -1.841128455464322e-12
+    -2.19247753930977e-11
+     8.24119550507728e-11
+ 4.61e+10    
+    8.229754683023916e-11
+   -2.189505123846082e-11
+    8.506737237056266e-11
+   -1.853097802591441e-12
+   -1.062832480523041e-11
+    8.501476321666271e-11
+   -1.022036105629651e-12
+   -1.843113877125897e-12
+    -2.19290254490975e-11
+    8.240598225701397e-11
+ 4.62e+10    
+     8.22916946317159e-11
+   -2.189940336689008e-11
+    8.506694844034197e-11
+   -1.855077427484719e-12
+   -1.063193844933011e-11
+    8.501426872944692e-11
+   -1.020485551837384e-12
+   -1.845086059436971e-12
+   -2.193328440021554e-11
+    8.239998643737732e-11
+ 4.63e+10    
+    8.228581977782164e-11
+   -2.190376455230724e-11
+    8.506651611091156e-11
+   -1.857043691408907e-12
+    -1.06355624689263e-11
+    8.501376580482516e-11
+     -1.0189121559913e-12
+   -1.847044950187585e-12
+   -2.193755217673021e-11
+    8.239396754316782e-11
+ 4.64e+10    
+    8.227992221993231e-11
+   -2.190813472470994e-11
+    8.506607532060846e-11
+   -1.858996542175972e-12
+   -1.063919685852517e-11
+    8.501325438159745e-11
+    -1.01731595001164e-12
+   -1.848990497329629e-12
+   -2.194182870847772e-11
+    8.238792552579239e-11
+ 4.65e+10    
+    8.227400190952875e-11
+   -2.191251381365932e-11
+    8.506562600779989e-11
+   -1.860935927764898e-12
+   -1.064284161257809e-11
+    8.501273439858719e-11
+   -1.015696966646479e-12
+    -1.85092264897778e-12
+   -2.194611392485679e-11
+    8.238186033676025e-11
+ 4.66e+10    
+    8.226805879819734e-11
+   -2.191690174828454e-11
+    8.506516811088329e-11
+    -1.86286179632268e-12
+   -1.064649672548096e-11
+     8.50122057946405e-11
+    -1.01405523947607e-12
+   -1.852841353410677e-12
+   -2.195040775483276e-11
+    8.237577192768309e-11
+ 4.67e+10    
+    8.226209283762973e-11
+   -2.192129845728705e-11
+    8.506470156828625e-11
+   -1.864774096165434e-12
+   -1.065016219157385e-11
+    8.501166850862724e-11
+   -1.012390802917124e-12
+   -1.854746559071897e-12
+   -2.195471012694228e-11
+      8.2369660250275e-11
+ 4.68e+10    
+    8.225610397962342e-11
+   -2.192570386894503e-11
+     8.50642263184669e-11
+   -1.866672775779405e-12
+   -1.065383800514048e-11
+    8.501112247944027e-11
+   -1.010703692227009e-12
+   -1.856638214571064e-12
+   -2.195902096929778e-11
+     8.23635252563537e-11
+ 4.69e+10    
+    8.225009217608215e-11
+   -2.193011791111787e-11
+    8.506374229991359e-11
+   -1.868557783822065e-12
+    -1.06575241604077e-11
+    8.501056764599625e-11
+   -1.008993943507841e-12
+   -1.858516268684895e-12
+   -2.196334020959176e-11
+    8.235736689783985e-11
+ 4.7e+10     
+    8.224405737901616e-11
+   -2.193454051125056e-11
+    8.506324945114539e-11
+   -1.870429069123161e-12
+   -1.066122065154503e-11
+    8.501000394723582e-11
+   -1.007261593710552e-12
+   -1.860380670358266e-12
+   -2.196766777510165e-11
+    8.235118512675832e-11
+ 4.71e+10    
+    8.223799954054274e-11
+   -2.193897159637826e-11
+    8.506274771071219e-11
+   -1.872286580685762e-12
+   -1.066492747266415e-11
+    8.500943132212385e-11
+   -1.005506680638809e-12
+   -1.862231368705293e-12
+   -2.197200359269414e-11
+     8.23449798952383e-11
+ 4.72e+10    
+    8.223191861288652e-11
+   -2.194341109313074e-11
+    8.506223701719491e-11
+   -1.874130267687332e-12
+    -1.06686446178184e-11
+    8.500884970964965e-11
+   -1.003729242952877e-12
+   -1.864068313010374e-12
+   -2.197634758882989e-11
+    8.233875115551358e-11
+ 4.73e+10    
+    8.222581454837994e-11
+   -2.194785892773696e-11
+    8.506171730920584e-11
+   -1.875960079480794e-12
+   -1.067237208100222e-11
+    8.500825904882758e-11
+   -1.001929320173419e-12
+   -1.865891452729314e-12
+   -2.198069968956803e-11
+    8.233249885992374e-11
+ 4.74e+10    
+    8.221968729946388e-11
+   -2.195231502602959e-11
+    8.506118852538878e-11
+   -1.877775965595607e-12
+   -1.067610985615067e-11
+    8.500765927869719e-11
+   -1.000106952685166e-12
+   -1.867700737490327e-12
+   -2.198505982057094e-11
+    8.232622296091385e-11
+ 4.75e+10    
+    8.221353681868828e-11
+    -2.19567793134496e-11
+    8.506065060441965e-11
+   -1.879577875738817e-12
+   -1.067985793713888e-11
+    8.500705033832381e-11
+   -9.982621817405329e-13
+   -1.869496117095176e-12
+   -2.198942790710875e-11
+    8.231992341103562e-11
+ 4.76e+10    
+    8.220736305871218e-11
+   -2.196125171505086e-11
+    8.506010348500663e-11
+   -1.881365759796108e-12
+   -1.068361631778152e-11
+     8.50064321667989e-11
+   -9.963950494631221e-13
+   -1.871277541520228e-12
+   -2.199380387406406e-11
+    8.231360016294796e-11
+ 4.77e+10    
+    8.220116597230524e-11
+   -2.196573215550473e-11
+    8.505954710589074e-11
+   -1.883139567832934e-12
+   -1.068738499183223e-11
+    8.500580470324063e-11
+   -9.945055988511728e-13
+   -1.873044960917517e-12
+   -2.199818764593665e-11
+    8.230725316941734e-11
+ 4.78e+10    
+    8.219494551234755e-11
+   -2.197022055910472e-11
+    8.505898140584595e-11
+   -1.884899250095523e-12
+   -1.069116395298309e-11
+    8.500516788679434e-11
+   -9.925938737808692e-13
+   -1.874798325615873e-12
+   -2.200257914684812e-11
+    8.230088238331873e-11
+ 4.79e+10    
+    8.218870163183033e-11
+     -2.1974716849771e-11
+    8.505840632367996e-11
+   -1.886644757012022e-12
+   -1.069495319486406e-11
+    8.500452165663338e-11
+   -9.906599190095886e-13
+   -1.876537586121967e-12
+   -2.200697830054679e-11
+    8.229448775763622e-11
+ 4.8e+10     
+     8.21824342838571e-11
+   -2.197922095105533e-11
+    8.505782179823477e-11
+   -1.888376039193491e-12
+   -1.069875271104244e-11
+    8.500386595195904e-11
+   -9.887037801790652e-13
+   -1.878262693121424e-12
+   -2.201138503041212e-11
+    8.228806924546357e-11
+ 4.81e+10    
+    8.217614342164388e-11
+   -2.198373278614541e-11
+    8.505722776838668e-11
+   -1.890093047435063e-12
+   -1.070256249502223e-11
+    8.500320071200191e-11
+   -9.867255038184404e-13
+   -1.879973597479903e-12
+   -2.201579925945978e-11
+    8.228162680000531e-11
+ 4.82e+10    
+    8.216982899852018e-11
+   -2.198825227786981e-11
+    8.505662417304753e-11
+   -1.891795732716977e-12
+   -1.070638254024362e-11
+    8.500252587602195e-11
+    -9.84725137347224e-13
+   -1.881670250244198e-12
+   -2.202022091034616e-11
+    8.227516037457704e-11
+ 4.83e+10    
+    8.216349096792956e-11
+   -2.199277934870253e-11
+    8.505601095116457e-11
+   -1.893484046205675e-12
+   -1.071021284008235e-11
+    8.500184138330933e-11
+   -9.827027290781551e-13
+   -1.883352602643353e-12
+   -2.202464990537329e-11
+    8.226866992260643e-11
+ 4.84e+10    
+    8.215712928343029e-11
+   -2.199731392076777e-11
+    8.505538804172175e-11
+   -1.895157939254895e-12
+   -1.071405338784921e-11
+    8.500114717318538e-11
+     -9.8065832821999e-13
+    -1.88502060608971e-12
+   -2.202908616649363e-11
+    8.226215539763429e-11
+ 4.85e+10    
+    8.215074389869661e-11
+   -2.200185591584465e-11
+    8.505475538373961e-11
+    -1.89681736340676e-12
+    -1.07179041767893e-11
+    8.500044318500283e-11
+   -9.785919848801622e-13
+   -1.886674212180092e-12
+   -2.203352961531473e-11
+    8.225561675331471e-11
+ 4.86e+10    
+    8.214433476751885e-11
+   -2.200640525537195e-11
+    8.505411291627685e-11
+   -1.898462270392848e-12
+    -1.07217652000816e-11
+    8.499972935814685e-11
+   -9.765037500673622e-13
+   -1.888313372696825e-12
+   -2.203798017310423e-11
+    8.224905394341651e-11
+ 4.87e+10    
+    8.213790184380456e-11
+   -2.201096186045276e-11
+    8.505346057842977e-11
+   -1.900092612135318e-12
+   -1.072563645083821e-11
+    8.499900563203588e-11
+   -9.743936756940144e-13
+   -1.889938039608924e-12
+   -2.204243776079452e-11
+    8.224246692182399e-11
+ 4.88e+10    
+    8.213144508157934e-11
+   -2.201552565185932e-11
+    8.505279830933423e-11
+    -1.90170834074799e-12
+   -1.072951792210382e-11
+    8.499827194612198e-11
+    -9.72261814578659e-13
+   -1.891548165073153e-12
+   -2.204690229898757e-11
+    8.223585564253734e-11
+ 4.89e+10    
+    8.212496443498757e-11
+   -2.202009655003779e-11
+    8.505212604816548e-11
+   -1.903309408537437e-12
+   -1.073340960685507e-11
+    8.499752823989206e-11
+   -9.701082204482189e-13
+   -1.893143701435155e-12
+    -2.20513737079599e-11
+    8.222922005967401e-11
+ 4.9e+10     
+     8.21184598582933e-11
+   -2.202467447511294e-11
+    8.505144373413933e-11
+   -1.904895768004099e-12
+   -1.073731149799993e-11
+    8.499677445286873e-11
+   -9.679329479401914e-13
+   -1.894724601230613e-12
+   -2.205585190766731e-11
+    8.222256012746956e-11
+ 4.91e+10    
+    8.211193130588097e-11
+   -2.202925934689289e-11
+    8.505075130651262e-11
+   -1.906467371843404e-12
+   -1.074122358837702e-11
+     8.49960105246106e-11
+    -9.65736052604708e-13
+   -1.896290817186293e-12
+   -2.206033681774967e-11
+     8.22158758002782e-11
+ 4.92e+10    
+    8.210537873225648e-11
+   -2.203385108487413e-11
+    8.505004870458457e-11
+   -1.908024172946827e-12
+    -1.07451458707551e-11
+     8.49952363947139e-11
+   -9.635175909065056e-13
+   -1.897842302221247e-12
+   -2.206482835753592e-11
+    8.220916703257401e-11
+ 4.93e+10    
+    8.209880209204784e-11
+   -2.203844960824585e-11
+    8.504933586769648e-11
+   -1.909566124403059e-12
+   -1.074907833783227e-11
+     8.49944520028127e-11
+   -9.612776202268126e-13
+   -1.899379009447886e-12
+   -2.206932644604882e-11
+    8.220243377895192e-11
+ 4.94e+10    
+    8.209220134000632e-11
+   -2.204305483589528e-11
+     8.50486127352341e-11
+   -1.911093179499085e-12
+   -1.075302098223543e-11
+    8.499365728858021e-11
+   -9.590161988650819e-13
+   -1.900900892173174e-12
+    -2.20738310020098e-11
+     8.21956759941282e-11
+ 4.95e+10    
+    8.208557643100686e-11
+   -2.204766668641192e-11
+    8.504787924662676e-11
+   -1.912605291721301e-12
+   -1.075697379651957e-11
+    8.499285219172943e-11
+   -9.567333860406834e-13
+   -1.902407903899699e-12
+   -2.207834194384384e-11
+    8.218889363294192e-11
+ 4.96e+10    
+    8.207892732004962e-11
+   -2.205228507809283e-11
+    8.504713534134965e-11
+   -1.914102414756655e-12
+   -1.076093677316716e-11
+     8.49920366520144e-11
+   -9.544292418944321e-13
+   -1.903899998326859e-12
+   -2.208285918968449e-11
+    8.218208665035588e-11
+ 4.97e+10    
+    8.207225396226021e-11
+   -2.205690992894692e-11
+    8.504638095892368e-11
+   -1.915584502493769e-12
+   -1.076490990458746e-11
+    8.499121060923087e-11
+   -9.521038274900493e-13
+   -1.905377129351983e-12
+   -2.208738265737837e-11
+    8.217525500145685e-11
+ 4.98e+10    
+    8.206555631289114e-11
+   -2.206154115670023e-11
+    8.504561603891703e-11
+   -1.917051509024024e-12
+   -1.076889318311581e-11
+    8.499037400321725e-11
+   -9.497572048154978e-13
+   -1.906839251071505e-12
+   -2.209191226449036e-11
+    8.216839864145749e-11
+ 4.99e+10    
+    8.205883432732235e-11
+   -2.206617867880041e-11
+    8.504484052094588e-11
+   -1.918503388642753e-12
+    -1.07728866010131e-11
+    8.498952677385606e-11
+   -9.473894367842098e-13
+   -1.908286317782081e-12
+   -2.209644792830846e-11
+    8.216151752569687e-11
+ 5e+10       
+    8.205208796106235e-11
+   -2.207082241242155e-11
+    8.504405434467486e-11
+   -1.919940095850331e-12
+   -1.077689015046487e-11
+    8.498866886107409e-11
+   -9.450005872362235e-13
+    -1.90971828398178e-12
+   -2.210098956584829e-11
+    8.215461160964115e-11
+ 5.01e+10    
+    8.204531716974905e-11
+   -2.207547227446904e-11
+    8.504325744981869e-11
+   -1.921361585353326e-12
+   -1.078090382358085e-11
+     8.49878002048442e-11
+   -9.425907209391944e-13
+   -1.911135104371198e-12
+   -2.210553709385838e-11
+    8.214768084888499e-11
+ 5.02e+10    
+    8.203852190915077e-11
+   -2.208012818158442e-11
+    8.504244977614278e-11
+    -1.92276781206563e-12
+   -1.078492761239415e-11
+    8.498692074518615e-11
+   -9.401599035893025e-13
+   -1.912536733854686e-12
+   -2.211009042882491e-11
+    8.214072519915274e-11
+ 5.03e+10    
+    8.203170213516704e-11
+   -2.208479005014998e-11
+    8.504163126346416e-11
+   -1.924158731109625e-12
+   -1.078896150886057e-11
+    8.498603042216713e-11
+   -9.377082018120413e-13
+   -1.913923127541459e-12
+   -2.211464948697642e-11
+    8.213374461629876e-11
+ 5.04e+10    
+    8.202485780382956e-11
+   -2.208945779629363e-11
+    8.504080185165226e-11
+   -1.925534297817297e-12
+   -1.079300550485794e-11
+    8.498512917590339e-11
+    -9.35235683162929e-13
+   -1.915294240746778e-12
+    -2.21192141842887e-11
+    8.212673905630863e-11
+ 5.05e+10    
+    8.201798887130317e-11
+   -2.209413133589377e-11
+    8.503996148063041e-11
+   -1.926894467731413e-12
+   -1.079705959218542e-11
+     8.49842169465612e-11
+   -9.327424161280585e-13
+   -1.916650028993155e-12
+   -2.212378443648988e-11
+    8.211970847530046e-11
+ 5.06e+10    
+    8.201109529388702e-11
+   -2.209881058458399e-11
+     8.50391100903766e-11
+   -1.928239196606661e-12
+    -1.08011237625628e-11
+    8.498329367435764e-11
+    -9.30228470124581e-13
+     -1.9179904480115e-12
+   -2.212836015906495e-11
+    8.211265282952579e-11
+ 5.07e+10    
+    8.200417702801481e-11
+   -2.210349545775772e-11
+    8.503824762092419e-11
+   -1.929568440410818e-12
+   -1.080519800762974e-11
+     8.49823592995621e-11
+    -9.27693915501055e-13
+   -1.919315453742315e-12
+   -2.213294126726079e-11
+    8.210557207537009e-11
+ 5.08e+10    
+    8.199723403025652e-11
+   -2.210818587057323e-11
+    8.503737401236324e-11
+   -1.930882155325899e-12
+    -1.08092823189451e-11
+    8.498141376249685e-11
+    -9.25138823537686e-13
+   -1.920625002336882e-12
+   -2.213752767609101e-11
+     8.20984661693545e-11
+ 5.09e+10    
+     8.19902662573189e-11
+   -2.211288173795821e-11
+    8.503648920484151e-11
+   -1.932180297749335e-12
+   -1.081337668798625e-11
+    8.498045700353861e-11
+   -9.225632664464625e-13
+   -1.921919050158455e-12
+   -2.214211930034062e-11
+    8.209133506813616e-11
+ 5.1e+10     
+    8.198327366604643e-11
+   -2.211758297461463e-11
+    8.503559313856565e-11
+   -1.933462824295124e-12
+    -1.08174811061483e-11
+    8.497948896311945e-11
+   -9.199673173711697e-13
+   -1.923197553783443e-12
+   -2.214671605457106e-11
+    8.208417872850956e-11
+ 5.11e+10    
+    8.197625621342234e-11
+   -2.212228949502342e-11
+    8.503468575380159e-11
+   -1.934729691795016e-12
+   -1.082159556474339e-11
+    8.497850958172784e-11
+   -9.173510503872877e-13
+   -1.924460470002629e-12
+   -2.215131785312482e-11
+    8.207699710740747e-11
+ 5.12e+10    
+    8.196921385656969e-11
+    -2.21270012134492e-11
+    8.503376699087642e-11
+   -1.935980857299701e-12
+        -1.0825720055e-11
+    8.497751879991006e-11
+   -9.147145405017937e-13
+   -1.925707755822337e-12
+   -2.215592461013046e-11
+    8.206979016190188e-11
+ 5.13e+10    
+     8.19621465527518e-11
+   -2.213171804394506e-11
+    8.503283679017899e-11
+   -1.937216278079931e-12
+   -1.082985456806217e-11
+    8.497651655827101e-11
+   -9.120578636528313e-13
+     -1.9269393684657e-12
+   -2.216053623950713e-11
+    8.206255784920496e-11
+ 5.14e+10    
+    8.195505425937366e-11
+   -2.213643990035725e-11
+    8.503189509216095e-11
+   -1.938435911627808e-12
+   -1.083399909498879e-11
+    8.497550279747556e-11
+   -9.093810967092694e-13
+   -1.928155265373801e-12
+   -2.216515265496965e-11
+     8.20553001266701e-11
+ 5.15e+10    
+    8.194793693398268e-11
+   -2.214116669632991e-11
+     8.50309418373383e-11
+   -1.939639715657844e-12
+   -1.083815362675286e-11
+    8.497447745824951e-11
+   -9.066843174701566e-13
+   -1.929355404206928e-12
+   -2.216977377003305e-11
+    8.204801695179283e-11
+ 5.16e+10    
+    8.194079453426966e-11
+   -2.214589834530979e-11
+     8.50299769662918e-11
+   -1.940827648108265e-12
+   -1.084231815424079e-11
+    8.497344048138104e-11
+   -9.039676046640514e-13
+   -1.930539742845792e-12
+   -2.217439949801745e-11
+     8.20407082822118e-11
+ 5.17e+10    
+    8.193362701806944e-11
+   -2.215063476055082e-11
+    8.502900041966837e-11
+   -1.941999667142116e-12
+   -1.084649266825153e-11
+    8.497239180772134e-11
+   -9.012310379482441e-13
+   -1.931708239392745e-12
+   -2.217902975205275e-11
+    8.203337407570976e-11
+ 5.18e+10    
+      8.1926434343362e-11
+   -2.215537585511894e-11
+    8.502801213818241e-11
+   -1.943155731148523e-12
+   -1.085067715949603e-11
+    8.497133137818681e-11
+   -8.984746979078453e-13
+   -1.932860852172992e-12
+   -2.218366444508362e-11
+    8.202601429021457e-11
+ 5.19e+10    
+    8.191921646827368e-11
+   -2.216012154189676e-11
+    8.502701206261668e-11
+   -1.944295798743854e-12
+    -1.08548716185963e-11
+    8.497025913375887e-11
+   -8.956986660547941e-13
+   -1.933997539735842e-12
+   -2.218830348987374e-11
+    8.201862888379996e-11
+ 5.2e+10     
+    8.191197335107727e-11
+   -2.216487173358804e-11
+    8.502600013382313e-11
+   -1.945419828772953e-12
+   -1.085907603608477e-11
+    8.496917501548623e-11
+   -8.929030248267117e-13
+   -1.935118260855929e-12
+   -2.219294679901104e-11
+    8.201121781468683e-11
+ 5.21e+10    
+    8.190470495019377e-11
+   -2.216962634272259e-11
+    8.502497629272482e-11
+   -1.946527780310322e-12
+   -1.086329040240349e-11
+    8.496807896448539e-11
+   -8.900878575856674e-13
+   -1.936222974534483e-12
+   -2.219759428491209e-11
+    8.200378104124384e-11
+ 5.22e+10    
+    8.189741122419258e-11
+   -2.217438528166067e-11
+    8.502394048031597e-11
+   -1.947619612661353e-12
+   -1.086751470790338e-11
+    8.496697092194227e-11
+    -8.87253248616809e-13
+   -1.937311640000508e-12
+   -2.220224585982683e-11
+    8.199631852198829e-11
+ 5.23e+10    
+    8.189009213179287e-11
+   -2.217914846259779e-11
+    8.502289263766428e-11
+   -1.948695285363544e-12
+   -1.087174894284355e-11
+    8.496585082911331e-11
+   -8.843992831268888e-13
+   -1.938384216712115e-12
+   -2.220690143584341e-11
+    8.198883021558759e-11
+ 5.24e+10    
+    8.188274763186425e-11
+   -2.218391579756922e-11
+    8.502183270591067e-11
+   -1.949754758187713e-12
+   -1.087599309739036e-11
+    8.496471862732626e-11
+   -8.815260472426872e-13
+   -1.939440664357691e-12
+   -2.221156092489266e-11
+    8.198131608085967e-11
+ 5.25e+10    
+    8.187537768342727e-11
+   -2.218868719845453e-11
+    8.502076062627171e-11
+   -1.950797991139211e-12
+    -1.08802471616169e-11
+    8.496357425798195e-11
+   -8.786336280092725e-13
+   -1.940480942857207e-12
+   -2.221622423875283e-11
+    8.197377607677378e-11
+ 5.26e+10    
+    8.186798224565497e-11
+   -2.219346257698235e-11
+    8.501967634004026e-11
+   -1.951824944459158e-12
+   -1.088451112550202e-11
+    8.496241766255523e-11
+      -8.757221133882e-13
+   -1.941505012363466e-12
+   -2.222089128905428e-11
+    8.196621016245214e-11
+ 5.27e+10    
+    8.186056127787323e-11
+   -2.219824184473469e-11
+    8.501857978858586e-11
+   -1.952835578625705e-12
+   -1.088878497892963e-11
+    8.496124878259593e-11
+   -8.727915922555567e-13
+   -1.942512833263344e-12
+   -2.222556198728395e-11
+    8.195861829716998e-11
+ 5.28e+10    
+    8.185311473956166e-11
+    -2.22030249131517e-11
+    8.501747091335729e-11
+   -1.953829854355212e-12
+   -1.089306871168801e-11
+    8.496006755973065e-11
+   -8.698421543999059e-13
+   -1.943504366179087e-12
+   -2.223023624479014e-11
+    8.195100044035693e-11
+ 5.29e+10    
+    8.184564259035468e-11
+   -2.220781169353606e-11
+    8.501634965588264e-11
+   -1.954807732603525e-12
+   -1.089736231346893e-11
+    8.495887393566316e-11
+   -8.668738905201204e-13
+   -1.944479571969581e-12
+   -2.223491397278695e-11
+    8.194335655159777e-11
+ 5.3e+10     
+    8.183814479004195e-11
+    -2.22126020970576e-11
+     8.50152159577707e-11
+   -1.955769174567215e-12
+   -1.090166577386696e-11
+    8.495766785217646e-11
+   -8.638868922230682e-13
+   -1.945438411731576e-12
+   -2.223959508235888e-11
+    8.193568659063307e-11
+ 5.31e+10    
+    8.183062129856945e-11
+   -2.221739603475769e-11
+     8.50140697607124e-11
+   -1.956714141684806e-12
+   -1.090597908237867e-11
+    8.495644925113337e-11
+    -8.60881252021228e-13
+    -1.94638084680105e-12
+   -2.224427948446548e-11
+    8.192799051736059e-11
+ 5.32e+10    
+    8.182307207604023e-11
+   -2.222219341755375e-11
+     8.50129110064815e-11
+   -1.957642595638033e-12
+   -1.091030222840182e-11
+    8.495521807447777e-11
+   -8.578570633301529e-13
+   -1.947306838754407e-12
+   -2.224896708994575e-11
+    8.192026829183555e-11
+ 5.33e+10    
+    8.181549708271517e-11
+   -2.222699415624382e-11
+    8.501173963693625e-11
+   -1.958554498353098e-12
+   -1.091463520123468e-11
+    8.495397426423635e-11
+   -8.548144204658295e-13
+   -1.948216349409817e-12
+   -2.225365780952273e-11
+    8.191251987427182e-11
+ 5.34e+10    
+    8.180789627901346e-11
+   -2.223179816151077e-11
+    8.501055559401966e-11
+   -1.959449812001942e-12
+   -1.091897799007513e-11
+    8.495271776251908e-11
+   -8.517534186419048e-13
+   -1.949109340828493e-12
+   -2.225835155380803e-11
+    8.190474522504248e-11
+ 5.35e+10    
+    8.180026962551412e-11
+   -2.223660534392708e-11
+    8.500935881976203e-11
+    -1.96032849900345e-12
+   -1.092333058402003e-11
+    8.495144851152077e-11
+   -8.486741539668516e-13
+   -1.949985775315975e-12
+   -2.226304823330615e-11
+    8.189694430468105e-11
+ 5.36e+10    
+    8.179261708295594e-11
+   -2.224141561395883e-11
+    8.500814925628079e-11
+   -1.961190522024784e-12
+   -1.092769297206434e-11
+     8.49501664535226e-11
+    -8.45576723440936e-13
+   -1.950845615423424e-12
+   -2.226774775841923e-11
+    8.188911707388177e-11
+ 5.37e+10    
+    8.178493861223858e-11
+   -2.224622888197044e-11
+    8.500692684578203e-11
+   -1.962035843982586e-12
+   -1.093206514310036e-11
+    8.494887153089252e-11
+   -8.424612249531435e-13
+    -1.95168882394893e-12
+   -2.227245003945113e-11
+    8.188126349350083e-11
+ 5.38e+10    
+     8.17772341744235e-11
+   -2.225104505822881e-11
+    8.500569153056198e-11
+   -1.962864428044314e-12
+   -1.093644708591696e-11
+    8.494756368608712e-11
+   -8.393277572779196e-13
+   -1.952515363938841e-12
+   -2.227715498661214e-11
+     8.18733835245568e-11
+ 5.39e+10    
+    8.176950373073412e-11
+   -2.225586405290787e-11
+    8.500444325300807e-11
+    -1.96367623762942e-12
+   -1.094083878919889e-11
+    8.494624286165267e-11
+   -8.361764200718763e-13
+   -1.953325198689018e-12
+    -2.22818625100232e-11
+     8.18654771282316e-11
+ 5.4e+10     
+    8.176174724255712e-11
+   -2.226068577609266e-11
+    8.500318195559946e-11
+   -1.964471236410732e-12
+   -1.094524024152582e-11
+    8.494490900022598e-11
+   -8.330073138703131e-13
+   -1.954118291746184e-12
+   -2.228657251972042e-11
+    8.185754426587144e-11
+ 5.41e+10    
+    8.175396467144289e-11
+    -2.22655101377839e-11
+    8.500190758090894e-11
+   -1.965249388315663e-12
+   -1.094965143137172e-11
+    8.494356204453611e-11
+   -8.298205400836448e-13
+   -1.954894606909222e-12
+   -2.229128492565935e-11
+      8.1849584898987e-11
+ 5.42e+10    
+    8.174615597910586e-11
+   -2.227033704790205e-11
+    8.500062007160374e-11
+   -1.966010657527505e-12
+   -1.095407234710404e-11
+    8.494220193740508e-11
+   -8.266162009937346e-13
+   -1.955654108230508e-12
+    -2.22959996377192e-11
+    8.184159898925475e-11
+ 5.43e+10    
+    8.173832112742593e-11
+   -2.227516641629174e-11
+    8.499931937044637e-11
+   -1.966755008486734e-12
+    -1.09585029769829e-11
+     8.49408286217495e-11
+   -8.233943997500886e-13
+   -1.956396760017205e-12
+   -2.230071656570755e-11
+    8.183358649851737e-11
+ 5.44e+10    
+    8.173046007844869e-11
+   -2.227999815272608e-11
+    8.499800542029658e-11
+   -1.967482405892281e-12
+   -1.096294330916036e-11
+    8.493944204058141e-11
+   -8.201552403659418e-13
+   -1.957122526832619e-12
+   -2.230543561936414e-11
+    8.182554738878453e-11
+ 5.45e+10    
+    8.172257279438566e-11
+   -2.228483216691053e-11
+     8.49966781641114e-11
+   -1.968192814702826e-12
+    -1.09673933316796e-11
+    8.493804213700945e-11
+   -8.168988277142309e-13
+   -1.957831373497497e-12
+   -2.231015670836549e-11
+    8.181748162223339e-11
+ 5.46e+10    
+    8.171465923761583e-11
+   -2.228966836848757e-11
+    8.499533754494714e-11
+   -1.968886200138086e-12
+   -1.097185303247418e-11
+    8.493662885424027e-11
+   -8.136252675234664e-13
+   -1.958523265091358e-12
+   -2.231487974232901e-11
+    8.180938916120968e-11
+ 5.47e+10    
+     8.17067193706855e-11
+   -2.229450666704051e-11
+    8.499398350595996e-11
+   -1.969562527680129e-12
+   -1.097632239936724e-11
+    8.493520213557958e-11
+    -8.10334666373461e-13
+   -1.959198166953869e-12
+   -2.231960463081727e-11
+    8.180126996822811e-11
+ 5.48e+10    
+    8.169875315630942e-11
+   -2.229934697209787e-11
+    8.499261599040758e-11
+   -1.970221763074655e-12
+   -1.098080142007078e-11
+    8.493376192443338e-11
+   -8.070271316909794e-13
+   -1.959856044686112e-12
+   -2.232433128334222e-11
+    8.179312400597292e-11
+ 5.49e+10    
+    8.169076055737101e-11
+   -2.230418919313746e-11
+    8.499123494164944e-11
+   -1.970863872332294e-12
+   -1.098529008218476e-11
+    8.493230816430876e-11
+   -8.037027717452519e-13
+   -1.960496864151978e-12
+   -2.232905960936925e-11
+    8.178495123729875e-11
+ 5.5e+10     
+    8.168274153692323e-11
+   -2.230903323959047e-11
+    8.498984030314893e-11
+   -1.971488821729927e-12
+   -1.098978837319652e-11
+    8.493084079881564e-11
+   -8.003616956433894e-13
+   -1.961120591479462e-12
+   -2.233378951832151e-11
+    8.177675162523118e-11
+ 5.51e+10    
+    8.167469605818869e-11
+   -2.231387902084549e-11
+    8.498843201847346e-11
+   -1.972096577811993e-12
+   -1.099429628047979e-11
+    8.492935977166747e-11
+   -7.970040133256621e-13
+   -1.961727193062057e-12
+   -2.233852091958391e-11
+    8.176852513296727e-11
+ 5.52e+10    
+    8.166662408456109e-11
+   -2.231872644625281e-11
+    8.498701003129635e-11
+   -1.972687107391778e-12
+   -1.099881379129411e-11
+    8.492786502668267e-11
+   -7.936298355607159e-13
+   -1.962316635560049e-12
+   -2.234325372250737e-11
+    8.176027172387646e-11
+ 5.53e+10    
+    8.165852557960471e-11
+   -2.232357542512821e-11
+    8.498557428539753e-11
+   -1.973260377552736e-12
+   -1.100334089278396e-11
+     8.49263565077854e-11
+   -7.902392739406216e-13
+   -1.962888885901913e-12
+   -2.234798783641269e-11
+    8.175199136150064e-11
+ 5.54e+10    
+     8.16504005070557e-11
+   -2.232842586675717e-11
+    8.498412472466463e-11
+   -1.973816355649807e-12
+   -1.100787757197801e-11
+    8.492483415900707e-11
+   -7.868324408758515e-13
+   -1.963443911285606e-12
+    -2.23527231705948e-11
+    8.174368400955496e-11
+ 5.55e+10    
+    8.164224883082226e-11
+   -2.233327768039872e-11
+    8.498266129309416e-11
+    -1.97435500931073e-12
+   -1.101242381578837e-11
+    8.492329792448731e-11
+   -7.834094495901327e-13
+   -1.963981679179978e-12
+    -2.23574596343268e-11
+    8.173534963192885e-11
+ 5.56e+10    
+    8.163407051498508e-11
+   -2.233813077528951e-11
+    8.498118393479258e-11
+   -1.974876306437347e-12
+   -1.101697961100979e-11
+    8.492174774847507e-11
+   -7.799704141151916e-13
+   -1.964502157326083e-12
+    -2.23621971368638e-11
+    8.172698819268587e-11
+ 5.57e+10    
+    8.162586552379822e-11
+   -2.234298506064772e-11
+    8.497969259397727e-11
+   -1.975380215206947e-12
+   -1.102154494431898e-11
+    8.492018357532978e-11
+   -7.765154492853985e-13
+   -1.965005313738562e-12
+   -2.236693558744702e-11
+    8.171859965606458e-11
+ 5.58e+10    
+    8.161763382168929e-11
+   -2.234784044567706e-11
+    8.497818721497782e-11
+   -1.975866704073569e-12
+   -1.102611980227375e-11
+    8.491860534952232e-11
+   -7.730446707322714e-13
+   -1.965491116706985e-12
+   -2.237167489530774e-11
+    8.171018398647885e-11
+ 5.59e+10    
+    8.160937537325989e-11
+   -2.235269683957058e-11
+    8.497666774223684e-11
+   -1.976335741769323e-12
+   -1.103070417131232e-11
+    8.491701301563637e-11
+   -7.695581948789352e-13
+   -1.965959534797216e-12
+    -2.23764149696713e-11
+     8.17017411485188e-11
+ 5.6e+10     
+    8.160109014328603e-11
+   -2.235755415151452e-11
+      8.4975134120311e-11
+   -1.976787297305713e-12
+   -1.103529803775251e-11
+    8.491540651836931e-11
+   -7.660561389344025e-13
+   -1.966410536852776e-12
+   -2.238115571976083e-11
+    8.169327110695078e-11
+ 5.61e+10    
+    8.159277809671909e-11
+   -2.236241229069234e-11
+    8.497358629387235e-11
+   -1.977221339974993e-12
+   -1.103990138779107e-11
+    8.491378580253338e-11
+    -7.62538620887803e-13
+   -1.966844091996211e-12
+   -2.238589705480129e-11
+    8.168477382671834e-11
+ 5.62e+10    
+    8.158443919868514e-11
+   -2.236727116628822e-11
+    8.497202420770904e-11
+   -1.977637839351437e-12
+   -1.104451420750283e-11
+     8.49121508130568e-11
+    -7.59005759502472e-13
+   -1.967260169630435e-12
+   -2.239063888402329e-11
+    8.167624927294209e-11
+ 5.63e+10    
+    8.157607341448659e-11
+   -2.237213068749127e-11
+     8.49704478067267e-11
+   -1.978036765292732e-12
+   -1.104913648284004e-11
+    8.491050149498459e-11
+   -7.554576743099536e-13
+   -1.967658739440129e-12
+   -2.239538111666686e-11
+    8.166769741092074e-11
+ 5.64e+10    
+    8.156768070960201e-11
+   -2.237699076349903e-11
+    8.496885703594906e-11
+   -1.978418087941248e-12
+   -1.105376819963157e-11
+    8.490883779348013e-11
+   -7.518944856038883e-13
+    -1.96803977139309e-12
+   -2.240012366198535e-11
+    8.165911820613124e-11
+ 5.65e+10    
+     8.15592610496862e-11
+    -2.23818513035212e-11
+    8.496725184051916e-11
+   -1.978781777725405e-12
+   -1.105840934358215e-11
+    8.490715965382561e-11
+   -7.483163144338202e-13
+   -1.968403235741568e-12
+   -2.240486642924907e-11
+    8.165051162422911e-11
+ 5.66e+10    
+    8.155081440057109e-11
+   -2.238671221678355e-11
+    8.496563216570073e-11
+   -1.979127805361005e-12
+   -1.106305990027172e-11
+    8.490546702142366e-11
+   -7.447232825988486e-13
+   -1.968749103023709e-12
+   -2.240960932774926e-11
+    8.164187763104908e-11
+ 5.67e+10    
+    8.154234072826602e-11
+   -2.239157341253146e-11
+    8.496399795687834e-11
+   -1.979456141852537e-12
+   -1.106771985515459e-11
+    8.490375984179791e-11
+   -7.411155126412457e-13
+   -1.969077344064856e-12
+   -2.241435226680151e-11
+    8.163321619260536e-11
+ 5.68e+10    
+    8.153383999895764e-11
+   -2.239643480003372e-11
+    8.496234915955925e-11
+   -1.979766758494523e-12
+   -1.107238919355881e-11
+    8.490203806059433e-11
+   -7.374931278399207e-13
+   -1.969387929978942e-12
+   -2.241909515574978e-11
+    8.162452727509199e-11
+ 5.69e+10    
+    8.152531217901085e-11
+   -2.240129628858595e-11
+    8.496068571937372e-11
+   -1.980059626872871e-12
+   -1.107706790068526e-11
+    8.490030162358212e-11
+    -7.33856252203804e-13
+    -1.96968083216988e-12
+   -2.242383790396982e-11
+    8.161581084488337e-11
+ 5.7e+10     
+    8.151675723496872e-11
+   -2.240615778751454e-11
+    8.495900758207653e-11
+   -1.980334718866181e-12
+   -1.108175596160717e-11
+     8.48985504766547e-11
+   -7.302050104651336e-13
+     -1.9699560223329e-12
+    -2.24285804208729e-11
+    8.160706686853428e-11
+ 5.71e+10    
+    8.150817513355291e-11
+   -2.241101920617996e-11
+    8.495731469354779e-11
+   -1.980592006647084e-12
+   -1.108645336126922e-11
+    8.489678456583101e-11
+   -7.265395280726343e-13
+   -1.970213472455952e-12
+   -2.243332261590954e-11
+    8.159829531278064e-11
+ 5.72e+10    
+    8.149956584166373e-11
+   -2.241588045398041e-11
+    8.495560699979358e-11
+   -1.980831462683579e-12
+   -1.109116008448687e-11
+    8.489500383725601e-11
+   -7.228599311845988e-13
+   -1.970453154821067e-12
+   -2.243806439857286e-11
+    8.158949614453954e-11
+ 5.73e+10    
+    8.149092932638093e-11
+   -2.242074144035548e-11
+    8.495388444694725e-11
+   -1.981053059740391e-12
+   -1.109587611594564e-11
+      8.4893208237202e-11
+   -7.191663466618824e-13
+   -1.970675042005691e-12
+   -2.244280567840229e-11
+    8.158066933090936e-11
+ 5.74e+10    
+    8.148226555496365e-11
+   -2.242560207478953e-11
+    8.495214698127054e-11
+   -1.981256770880255e-12
+   -1.110060144020041e-11
+    8.489139771206951e-11
+   -7.154589020607873e-13
+   -1.970879106884136e-12
+   -2.244754636498715e-11
+    8.157181483917079e-11
+ 5.75e+10    
+    8.147357449485031e-11
+   -2.243046226681513e-11
+    8.495039454915386e-11
+    -1.98144256946528e-12
+   -1.110533604167471e-11
+    8.488957220838854e-11
+   -7.117377256258607e-13
+   -1.971065322628879e-12
+   -2.245228636797002e-11
+    8.156293263678624e-11
+ 5.76e+10    
+    8.146485611365966e-11
+   -2.243532192601668e-11
+    8.494862709711772e-11
+     -1.9816104291583e-12
+   -1.111007990465997e-11
+     8.48877316728188e-11
+   -7.080029462825956e-13
+   -1.971233662711967e-12
+   -2.245702559705028e-11
+    8.155402269140087e-11
+ 5.77e+10    
+    8.145611037919025e-11
+   -2.244018096203373e-11
+     8.49468445718137e-11
+    -1.98176032392415e-12
+   -1.111483301331491e-11
+    8.488587605215155e-11
+   -7.042546936300295e-13
+   -1.971384100906368e-12
+   -2.246176396198761e-11
+    8.154508497084204e-11
+ 5.78e+10    
+    8.144733725942109e-11
+   -2.244503928456432e-11
+    8.494504692002495e-11
+   -1.981892228031078e-12
+   -1.111959535166471e-11
+    8.488400529330995e-11
+   -7.004930979332651e-13
+   -1.971516611287364e-12
+   -2.246650137260528e-11
+    8.153611944312042e-11
+ 5.79e+10    
+    8.143853672251156e-11
+   -2.244989680336862e-11
+     8.49432340886677e-11
+   -1.982006116051976e-12
+   -1.112436690360052e-11
+    8.488211934335007e-11
+   -6.967182901158938e-13
+    -1.97163116823391e-12
+   -2.247123773879363e-11
+    8.152712607642944e-11
+ 5.8e+10     
+     8.14297087368019e-11
+   -2.245475342827192e-11
+    8.494140602479142e-11
+   -1.982101962865814e-12
+   -1.112914765287854e-11
+     8.48802181494624e-11
+   -6.929304017523111e-13
+   -1.971727746429984e-12
+   -2.247597297051357e-11
+    8.151810483914615e-11
+ 5.81e+10    
+    8.142085327081298e-11
+   -2.245960906916818e-11
+    8.493956267558018e-11
+   -1.982179743658885e-12
+   -1.113393758311949e-11
+    8.487830165897151e-11
+   -6.891295650599873e-13
+   -1.971806320865969e-12
+    -2.24807069777995e-11
+    8.150905569983082e-11
+ 5.82e+10    
+    8.141197029324697e-11
+   -2.246446363602328e-11
+    8.493770398835363e-11
+   -1.982239433926192e-12
+   -1.113873667780789e-11
+    8.487636981933825e-11
+     -6.8531591289158e-13
+   -1.971866866840024e-12
+   -2.248543967076311e-11
+    8.149997862722772e-11
+ 5.83e+10    
+    8.140305977298683e-11
+   -2.246931703887828e-11
+    8.493582991056728e-11
+   -1.982281009472718e-12
+   -1.114354492029136e-11
+    8.487442257815998e-11
+   -6.814895787270243e-13
+   -1.971909359959427e-12
+   -2.249017095959634e-11
+    8.149087359026471e-11
+ 5.84e+10    
+    8.139412167909704e-11
+   -2.247416918785262e-11
+    8.493394038981406e-11
+   -1.982304446414803e-12
+   -1.114836229378003e-11
+     8.48724598831715e-11
+   -6.776506966655049e-13
+   -1.971933776141953e-12
+   -2.249490075457467e-11
+    8.148174055805376e-11
+ 5.85e+10    
+     8.13851559808237e-11
+   -2.247901999314741e-11
+    8.493203537382467e-11
+   -1.982309721181441e-12
+   -1.115318878134577e-11
+    8.487048168224607e-11
+   -6.737994014173403e-13
+   -1.971940091617232e-12
+    -2.24996289660605e-11
+    8.147257949989118e-11
+ 5.86e+10    
+    8.137616264759386e-11
+   -2.248386936504848e-11
+    8.493011481046851e-11
+   -1.982296810515595e-12
+   -1.115802436592159e-11
+    8.486848792339643e-11
+   -6.699358282957906e-13
+   -1.971928282928095e-12
+   -2.250435550450622e-11
+    8.146339038525746e-11
+ 5.87e+10    
+    8.136714164901668e-11
+   -2.248871721392969e-11
+    8.492817864775488e-11
+   -1.982265691475523e-12
+   -1.116286903030104e-11
+    8.486647855477496e-11
+   -6.660601132087818e-13
+   -1.971898326931932e-12
+   -2.250908028045728e-11
+    8.145417318381739e-11
+ 5.88e+10    
+    8.135809295488279e-11
+   -2.249356345025595e-11
+    8.492622683383316e-11
+   -1.982216341436103e-12
+   -1.116772275713744e-11
+     8.48644535246753e-11
+   -6.621723926505491e-13
+   -1.971850200802053e-12
+   -2.251380320455559e-11
+    8.144492786542056e-11
+ 5.89e+10    
+    8.134901653516445e-11
+   -2.249840798458627e-11
+    8.492425931699395e-11
+   -1.982148738090127e-12
+   -1.117258552894328e-11
+    8.486241278153281e-11
+   -6.582728036931823e-13
+   -1.971783882029044e-12
+   -2.251852418754234e-11
+    8.143565440010106e-11
+ 5.9e+10     
+    8.133991236001612e-11
+   -2.250325072757708e-11
+    8.492227604567002e-11
+   -1.982062859449638e-12
+   -1.117745732808966e-11
+     8.48603562739254e-11
+   -6.543614839781112e-13
+   -1.971699348422083e-12
+   -2.252324314026128e-11
+    8.142635275807759e-11
+ 5.91e+10    
+     8.13307803997736e-11
+   -2.250809158998488e-11
+    8.492027696843696e-11
+   -1.981958683847194e-12
+   -1.118233813680558e-11
+    8.485828395057455e-11
+   -6.504385717075104e-13
+   -1.971596578110312e-12
+   -2.252795997366169e-11
+    8.141702290975378e-11
+ 5.92e+10    
+    8.132162062495508e-11
+   -2.251293048266966e-11
+    8.491826203401367e-11
+   -1.981836189937235e-12
+   -1.118722793717732e-11
+    8.485619576034567e-11
+   -6.465042056356021e-13
+   -1.971475549544188e-12
+   -2.253267459880138e-11
+    8.140766482571806e-11
+ 5.93e+10    
+    8.131243300626037e-11
+   -2.251776731659755e-11
+    8.491623119126365e-11
+   -1.981695356697335e-12
+   -1.119212671114786e-11
+    8.485409165224939e-11
+   -6.425585250599187e-13
+   -1.971336241496773e-12
+   -2.253738692684974e-11
+    8.139827847674371e-11
+ 5.94e+10    
+    8.130321751457126e-11
+   -2.252260200284404e-11
+    8.491418438919532e-11
+   -1.981536163429506e-12
+    -1.11970344405162e-11
+      8.4851971575442e-11
+   -6.386016698124542e-13
+   -1.971178633065125e-12
+   -2.254209686909063e-11
+    8.138886383378894e-11
+ 5.95e+10    
+    8.129397412095161e-11
+   -2.252743445259672e-11
+    8.491212157696287e-11
+   -1.981358589761531e-12
+   -1.120195110693681e-11
+    8.484983547922654e-11
+   -6.346337802507675e-13
+   -1.971002703671579e-12
+   -2.254680433692548e-11
+    8.137942086799693e-11
+ 5.96e+10    
+    8.128470279664686e-11
+   -2.253226457715825e-11
+    8.491004270386726e-11
+   -1.981162615648204e-12
+   -1.120687669191903e-11
+    8.484768331305283e-11
+   -6.306549972489893e-13
+   -1.970808433065131e-12
+   -2.255150924187586e-11
+    8.136994955069574e-11
+ 5.97e+10    
+    8.127540351308469e-11
+   -2.253709228794923e-11
+    8.490794771935662e-11
+   -1.980948221372648e-12
+   -1.121181117682641e-11
+    8.484551502651918e-11
+   -6.266654621887927e-13
+   -1.970595801322695e-12
+   -2.255621149558671e-11
+     8.13604498533984e-11
+ 5.98e+10    
+    8.126607624187437e-11
+   -2.254191749651111e-11
+    8.490583657302704e-11
+     -1.9807153875476e-12
+   -1.121675454287618e-11
+    8.484333056937274e-11
+    -6.22665316950241e-13
+   -1.970364788850471e-12
+   -2.256091100982908e-11
+    8.135092174780293e-11
+ 5.99e+10    
+    8.125672095480727e-11
+   -2.254674011450894e-11
+    8.490370921462333e-11
+   -1.980464095116668e-12
+   -1.122170677113867e-11
+    8.484112989150963e-11
+   -6.186547039026169e-13
+   -1.970115376385227e-12
+   -2.256560769650278e-11
+    8.134136520579209e-11
+ 6e+10       
+    8.124733762385631e-11
+   -2.255156005373408e-11
+    8.490156559403964e-11
+   -1.980194325355639e-12
+   -1.122666784253668e-11
+    8.483891294297673e-11
+   -6.146337658951506e-13
+   -1.969847544995639e-12
+   -2.257030146763944e-11
+    8.133178019943376e-11
+ 6.01e+10    
+    8.123792622117596e-11
+   -2.255637722610708e-11
+    8.489940566132022e-11
+   -1.979906059873708e-12
+   -1.123163773784493e-11
+    8.483667967397137e-11
+   -6.106026462476934e-13
+   -1.969561276083571e-12
+     -2.2574992235405e-11
+    8.132216670098043e-11
+ 6.02e+10    
+    8.122848671910259e-11
+   -2.256119154368043e-11
+    8.489722936666009e-11
+   -1.979599280614773e-12
+   -1.123661643768954e-11
+    8.483443003484287e-11
+   -6.065614887413219e-13
+   -1.969256551385375e-12
+   -2.257967991210264e-11
+    8.131252468286931e-11
+ 6.03e+10    
+    8.121901909015396e-11
+   -2.256600291864117e-11
+     8.48950366604056e-11
+   -1.979273969858692e-12
+   -1.124160392254741e-11
+    8.483216397609247e-11
+   -6.025104376088853e-13
+   -1.968933352973221e-12
+   -2.258436441017548e-11
+    8.130285411772269e-11
+ 6.04e+10    
+    8.120952330702927e-11
+   -2.257081126331363e-11
+    8.489282749305518e-11
+   -1.978930110222521e-12
+   -1.124660017274572e-11
+     8.48298814483745e-11
+   -5.984496375254708e-13
+   -1.968591663256326e-12
+   -2.258904564220906e-11
+    8.129315497834692e-11
+ 6.05e+10    
+    8.119999934260901e-11
+   -2.257561649016201e-11
+     8.48906018152598e-11
+   -1.978567684661789e-12
+   -1.125160516846134e-11
+    8.482758240249676e-11
+   -5.943792335988422e-13
+   -1.968231464982282e-12
+   -2.259372352093421e-11
+    8.128342723773337e-11
+ 6.06e+10    
+    8.119044716995487e-11
+   -2.258041851179305e-11
+    8.488835957782386e-11
+   -1.978186676471716e-12
+   -1.125661888972034e-11
+     8.48252667894215e-11
+   -5.902993713597668e-13
+   -1.967852741238329e-12
+   -2.259839795922956e-11
+    8.127367086905739e-11
+ 6.07e+10    
+    8.118086676230963e-11
+   -2.258521724095866e-11
+    8.488610073170568e-11
+   -1.977787069288468e-12
+   -1.126164131639741e-11
+    8.482293456026554e-11
+   -5.862101967523346e-13
+   -1.967455475452607e-12
+    -2.26030688701241e-11
+    8.126388584567894e-11
+ 6.08e+10    
+    8.117125809309699e-11
+   -2.259001259055846e-11
+    8.488382522801811e-11
+   -1.977368847090373e-12
+    -1.12666724282154e-11
+    8.482058566630114e-11
+     -5.8211185612419e-13
+   -1.967039651395446e-12
+   -2.260773616679982e-11
+    8.125407214114214e-11
+ 6.09e+10    
+    8.116162113592147e-11
+   -2.259480447364222e-11
+    8.488153301802889e-11
+   -1.976931994199169e-12
+   -1.127171220474472e-11
+    8.481822005895698e-11
+   -5.780044962167154e-13
+   -1.966605253180587e-12
+   -2.261239976259417e-11
+    8.124422972917501e-11
+ 6.1e+10     
+    8.115195586456815e-11
+   -2.259959280341245e-11
+    8.487922405316154e-11
+   -1.976476495281211e-12
+   -1.127676062540291e-11
+    8.481583768981826e-11
+   -5.738882641551487e-13
+   -1.966152265266482e-12
+   -2.261705957100268e-11
+    8.123435858368963e-11
+ 6.11e+10    
+    8.114226225300267e-11
+   -2.260437749322696e-11
+    8.487689828499618e-11
+   -1.976002335348684e-12
+   -1.128181766945416e-11
+    8.481343851062731e-11
+   -5.697633074386763e-13
+   -1.965680672457504e-12
+   -2.262171550568125e-11
+    8.122445867878184e-11
+ 6.12e+10    
+    8.113254027537088e-11
+   -2.260915845660115e-11
+     8.48745556652692e-11
+   -1.975509499760793e-12
+   -1.128688331600868e-11
+    8.481102247328428e-11
+   -5.656297739304429e-13
+   -1.965190459905184e-12
+    -2.26263674804487e-11
+    8.121452998873089e-11
+ 6.13e+10    
+    8.112278990599878e-11
+    -2.26139356072105e-11
+    8.487219614587462e-11
+   -1.974997974224998e-12
+   -1.129195754402235e-11
+    8.480858952984791e-11
+   -5.614878118475175e-13
+   -1.964681613109495e-12
+   -2.263101540928923e-11
+    8.120457248799978e-11
+ 6.14e+10    
+    8.111301111939222e-11
+    -2.26187088588931e-11
+    8.486981967886445e-11
+   -1.974467744798174e-12
+   -1.129704033229616e-11
+    8.480613963253569e-11
+    -5.57337569750828e-13
+   -1.964154117919996e-12
+   -2.263565920635477e-11
+    8.119458615123451e-11
+ 6.15e+10    
+    8.110320389023697e-11
+   -2.262347812565175e-11
+    8.486742621644895e-11
+    -1.97391879788782e-12
+   -1.130213165947581e-11
+    8.480367273372468e-11
+   -5.531791965350258e-13
+   -1.963607960537098e-12
+   -2.264029878596724e-11
+    8.118457095326424e-11
+ 6.16e+10    
+      8.1093368193398e-11
+   -2.262824332165651e-11
+    8.486501571099732e-11
+   -1.973351120253196e-12
+   -1.130723150405121e-11
+     8.48011887859519e-11
+   -5.490128414183228e-13
+   -1.963043127513256e-12
+   -2.264493406262104e-11
+     8.11745268691009e-11
+ 6.17e+10    
+    8.108350400391985e-11
+   -2.263300436124696e-11
+    8.486258811503839e-11
+   -1.972764699006556e-12
+   -1.131233984435602e-11
+      8.4798687741915e-11
+    -5.44838653932249e-13
+   -1.962459605754191e-12
+   -2.264956495098532e-11
+    8.116445387393944e-11
+ 6.18e+10    
+    8.107361129702597e-11
+   -2.263776115893448e-11
+    8.486014338126061e-11
+   -1.972159521614223e-12
+    -1.13174566585672e-11
+    8.479616955447258e-11
+    -5.40656783911432e-13
+   -1.961857382520041e-12
+   -2.265419136590615e-11
+    8.115435194315675e-11
+ 6.19e+10    
+    8.106369004811862e-11
+   -2.264251362940451e-11
+    8.485768146251324e-11
+   -1.971535575897826e-12
+   -1.132258192470458e-11
+    8.479363417664453e-11
+   -5.364673814832477e-13
+   -1.961236445426588e-12
+    -2.26588132224088e-11
+     8.11442210523123e-11
+ 6.2e+10     
+    8.105374023277882e-11
+   -2.264726168751874e-11
+     8.48552023118059e-11
+   -1.970892850035395e-12
+   -1.132771562063044e-11
+    8.479108156161311e-11
+   -5.322705970575168e-13
+   -1.960596782446385e-12
+   -2.266343043570011e-11
+    8.113406117714751e-11
+ 6.21e+10    
+    8.104376182676579e-11
+   -2.265200524831742e-11
+     8.48527058823102e-11
+   -1.970231332562507e-12
+   -1.133285772404911e-11
+    8.478851166272294e-11
+   -5.280665813160889e-13
+   -1.959938381909961e-12
+   -2.266804292117056e-11
+    8.112387229358544e-11
+ 6.22e+10    
+    8.103375480601686e-11
+   -2.265674422702141e-11
+    8.485019212735891e-11
+   -1.969551012373404e-12
+   -1.133800821250644e-11
+    8.478592443348132e-11
+   -5.238554852024448e-13
+   -1.959261232506972e-12
+   -2.267265059439633e-11
+    8.111365437773086e-11
+ 6.23e+10    
+    8.102371914664731e-11
+   -2.266147853903443e-11
+    8.484766100044745e-11
+   -1.968851878722132e-12
+   -1.134316706338958e-11
+    8.478331982755919e-11
+   -5.196374599112263e-13
+   -1.958565323287314e-12
+   -2.267725337114162e-11
+    8.110340740586952e-11
+ 6.24e+10    
+    8.101365482494977e-11
+   -2.266620809994508e-11
+    8.484511245523362e-11
+   -1.968133921223631e-12
+   -1.134833425392641e-11
+      8.4780697798791e-11
+   -5.154126568777528e-13
+    -1.95785064366231e-12
+   -2.268185116736068e-11
+    8.109313135446851e-11
+ 6.25e+10    
+    8.100356181739433e-11
+   -2.267093282552913e-11
+    8.484254644553846e-11
+    -1.96739712985482e-12
+   -1.135350976118528e-11
+    8.477805830117578e-11
+   -5.111812277674888e-13
+   -1.957117183405786e-12
+   -2.268644389919994e-11
+    8.108282620017546e-11
+ 6.26e+10    
+    8.099344010062791e-11
+   -2.267565263175126e-11
+    8.483996292534638e-11
+   -1.966641494955746e-12
+   -1.135869356207451e-11
+    8.477540128887701e-11
+   -5.069433244654875e-13
+   -1.956364932655219e-12
+   -2.269103148299992e-11
+    8.107249191981832e-11
+ 6.27e+10    
+    8.098328965147435e-11
+   -2.268036743476748e-11
+     8.48373618488056e-11
+   -1.965867007230566e-12
+   -1.136388563334211e-11
+      8.4772726716223e-11
+   -5.026990990658121e-13
+   -1.955593881912849e-12
+   -2.269561383529745e-11
+     8.10621284904056e-11
+ 6.28e+10    
+    8.097311044693377e-11
+   -2.268507715092687e-11
+    8.483474317022875e-11
+    -1.96507365774871e-12
+   -1.136908595157543e-11
+    8.477003453770788e-11
+   -4.984487038609114e-13
+   -1.954804022046759e-12
+   -2.270019087282753e-11
+    8.105173588912532e-11
+ 6.29e+10    
+    8.096290246418232e-11
+   -2.268978169677364e-11
+    8.483210684409284e-11
+    -1.96426143794587e-12
+   -1.137429449320069e-11
+    8.476732470799123e-11
+    -4.94192291330986e-13
+   -1.953995344291952e-12
+   -2.270476251252531e-11
+    8.104131409334527e-11
+ 6.3e+10     
+    8.095266568057213e-11
+   -2.269448098904918e-11
+    8.482945282503996e-11
+   -1.963430339625096e-12
+   -1.137951123448276e-11
+    8.476459718189895e-11
+   -4.899300141333141e-13
+   -1.953167840251453e-12
+   -2.270932867152818e-11
+    8.103086308061261e-11
+ 6.31e+10    
+    8.094240007363068e-11
+   -2.269917494469389e-11
+    8.482678106787759e-11
+    -1.96258035495779e-12
+   -1.138473615152475e-11
+    8.476185191442328e-11
+   -4.856620250915611e-13
+   -1.952321501897354e-12
+   -2.271388926717741e-11
+    8.102038282865317e-11
+ 6.32e+10    
+    8.093210562106072e-11
+   -2.270386348084912e-11
+    8.482409152757872e-11
+   -1.961711476484774e-12
+   -1.138996922026772e-11
+    8.475908886072364e-11
+   -4.813884771850629e-13
+   -1.951456321571865e-12
+   -2.271844421702039e-11
+    8.100987331537186e-11
+ 6.33e+10    
+    8.092178230073967e-11
+   -2.270854651485897e-11
+    8.482138415928218e-11
+   -1.960823697117259e-12
+   -1.139521041649034e-11
+     8.47563079761263e-11
+   -4.771095235381004e-13
+   -1.950572291988357e-12
+   -2.272299343881214e-11
+    8.099933451885148e-11
+ 6.34e+10    
+    8.091143009071979e-11
+   -2.271322396427245e-11
+    8.481865891829338e-11
+   -1.959917010137883e-12
+   -1.140045971580854e-11
+    8.475350921612515e-11
+   -4.728253174091372e-13
+    -1.94966940623241e-12
+   -2.272753685051738e-11
+    8.098876641735325e-11
+ 6.35e+10    
+    8.090104896922696e-11
+   -2.271789574684486e-11
+    8.481591576008424e-11
+   -1.958991409201686e-12
+   -1.140571709367534e-11
+    8.475069253638194e-11
+   -4.685360121800412e-13
+   -1.948747657762795e-12
+   -2.273207437031231e-11
+    8.097816898931581e-11
+ 6.36e+10    
+     8.08906389146615e-11
+   -2.272256178053992e-11
+    8.481315464029315e-11
+   -1.958046888337095e-12
+    -1.14109825253804e-11
+    8.474785789272642e-11
+   -4.642417613453131e-13
+   -1.947807040412497e-12
+   -2.273660591658631e-11
+    8.096754221335529e-11
+ 6.37e+10    
+    8.088019990559678e-11
+   -2.272722198353143e-11
+    8.481037551472629e-11
+   -1.957083441946892e-12
+   -1.141625598604985e-11
+    8.474500524115669e-11
+   -4.599427185012649e-13
+   -1.946847548389715e-12
+   -2.274113140794371e-11
+    8.095688606826471e-11
+ 6.38e+10    
+     8.08697319207793e-11
+   -2.273187627420503e-11
+    8.480757833935682e-11
+   -1.956101064809139e-12
+   -1.142153745064595e-11
+    8.474213453783967e-11
+   -4.556390373352221e-13
+    -1.94586917627883e-12
+   -2.274565076320557e-11
+    8.094620053301369e-11
+ 6.39e+10    
+    8.085923493912868e-11
+   -2.273652457115994e-11
+    8.480476307032579e-11
+   -1.955099752078183e-12
+    -1.14268268939669e-11
+    8.473924573911116e-11
+    -4.51330871614678e-13
+   -1.944871919041359e-12
+    -2.27501639014114e-11
+    8.093548558674836e-11
+ 6.4e+10     
+    8.084870893973663e-11
+   -2.274116679321069e-11
+    8.480192966394195e-11
+   -1.954079499285509e-12
+   -1.143212429064647e-11
+      8.4736338801476e-11
+   -4.470183751764712e-13
+   -1.943855772016942e-12
+    -2.27546707418208e-11
+    8.092474120879068e-11
+ 6.41e+10    
+    8.083815390186704e-11
+   -2.274580285938868e-11
+    8.479907807668241e-11
+   -1.953040302340723e-12
+   -1.143742961515388e-11
+    8.473341368160846e-11
+   -4.427017019159294e-13
+   -1.942820730924253e-12
+   -2.275917120391497e-11
+    8.091396737863799e-11
+ 6.42e+10    
+    8.082756980495536e-11
+    -2.27504326889439e-11
+    8.479620826519262e-11
+    -1.95198215753241e-12
+   -1.144274284179348e-11
+    8.473047033635256e-11
+   -4.383810057760233e-13
+   -1.941766791861932e-12
+   -2.276366520739865e-11
+     8.09031640759632e-11
+ 6.43e+10    
+     8.08169566286084e-11
+   -2.275505620134666e-11
+    8.479332018628669e-11
+   -1.950905061529041e-12
+   -1.144806394470455e-11
+    8.472750872272215e-11
+   -4.340564407364991e-13
+   -1.940693951309514e-12
+   -2.276815267220149e-11
+     8.08923312806138e-11
+ 6.44e+10    
+    8.080631435260389e-11
+    -2.27596733162889e-11
+    8.479041379694738e-11
+   -1.949809011379844e-12
+   -1.145339289786116e-11
+     8.47245287979011e-11
+   -4.297281608030349e-13
+   -1.939602206128299e-12
+   -2.277263351847957e-11
+    8.088146897261169e-11
+ 6.45e+10    
+    8.079564295689014e-11
+   -2.276428395368613e-11
+    8.478748905432662e-11
+   -1.948694004515676e-12
+   -1.145872967507175e-11
+    8.472153051924343e-11
+   -4.253963199963533e-13
+   -1.938491553562262e-12
+   -2.277710766661718e-11
+     8.08705771321529e-11
+ 6.46e+10    
+    8.078494242158547e-11
+   -2.276888803367866e-11
+    8.478454591574531e-11
+   -1.947560038749863e-12
+   -1.146407424997919e-11
+    8.471851384427387e-11
+   -4.210610723413743e-13
+   -1.937361991238915e-12
+   -2.278157503722817e-11
+    8.085965573960743e-11
+ 6.47e+10    
+    8.077421272697811e-11
+   -2.277348547663323e-11
+    8.478158433869388e-11
+   -1.946407112279029e-12
+   -1.146942659606041e-11
+    8.471547873068744e-11
+    -4.16722571856348e-13
+    -1.93621351717015e-12
+   -2.278603555115742e-11
+    8.084870477551799e-11
+ 6.48e+10    
+    8.076345385352573e-11
+   -2.277807620314474e-11
+    8.477860428083253e-11
+   -1.945235223683925e-12
+   -1.147478668662632e-11
+    8.471242513635022e-11
+   -4.123809725419914e-13
+   -1.935046129753112e-12
+   -2.279048912948251e-11
+     8.08377242206008e-11
+ 6.49e+10    
+    8.075266578185459e-11
+   -2.278266013403717e-11
+    8.477560569999046e-11
+   -1.944044371930209e-12
+    -1.14801544948216e-11
+    8.470935301929903e-11
+   -4.080364283706362e-13
+   -1.933859827770967e-12
+   -2.279493569351493e-11
+    8.082671405574409e-11
+ 6.5e+10     
+    8.074184849275999e-11
+   -2.278723719036561e-11
+    8.477258855416715e-11
+   -1.942834556369289e-12
+   -1.148552999362456e-11
+    8.470626233774182e-11
+    -4.03689093275374e-13
+   -1.932654610393785e-12
+   -2.279937516480163e-11
+    8.081567426200855e-11
+ 6.51e+10    
+    8.073100196720505e-11
+   -2.279180729341734e-11
+    8.476955280153204e-11
+   -1.941605776739035e-12
+   -1.149091315584692e-11
+    8.470315305005776e-11
+   -3.993391211392061e-13
+   -1.931430477179287e-12
+   -2.280380746512643e-11
+     8.08046048206265e-11
+ 6.52e+10    
+    8.072012618632087e-11
+   -2.279637036471335e-11
+    8.476649840042446e-11
+   -1.940358033164581e-12
+   -1.149630395413383e-11
+    8.470002511479718e-11
+   -3.949866657842295e-13
+   -1.930187428073616e-12
+   -2.280823251651131e-11
+    8.079350571300137e-11
+ 6.53e+10    
+    8.070922113140586e-11
+   -2.280092632600966e-11
+      8.4763425309354e-11
+   -1.939091326159053e-12
+    -1.15017023609636e-11
+     8.46968784906821e-11
+   -3.906318809607932e-13
+   -1.928925463412157e-12
+   -2.281265024121781e-11
+    8.078237692070766e-11
+ 6.54e+10    
+    8.069828678392528e-11
+   -2.280547509929871e-11
+    8.476033348700039e-11
+   -1.937805656624284e-12
+   -1.150710834864761e-11
+    8.469371313660593e-11
+   -3.862749203366977e-13
+     -1.9276445839202e-12
+   -2.281706056174834e-11
+    8.077121842549023e-11
+ 6.55e+10    
+     8.06873231255109e-11
+   -2.281001660681059e-11
+     8.47572228922138e-11
+    -1.93650102585156e-12
+   -1.151252188933022e-11
+    8.469052901163355e-11
+   -3.819159374863881e-13
+   -1.926344790713761e-12
+   -2.282146340084744e-11
+    8.076003020926405e-11
+ 6.56e+10    
+    8.067633013796091e-11
+    -2.28145507710146e-11
+    8.475409348401492e-11
+   -1.935177435522283e-12
+    -1.15179429549887e-11
+    8.468732607500176e-11
+   -3.775550858801756e-13
+   -1.925026085300234e-12
+   -2.282585868150315e-11
+    8.074881225411375e-11
+ 6.57e+10    
+    8.066530780323891e-11
+   -2.281907751462013e-11
+    8.475094522159486e-11
+   -1.933834887708669e-12
+   -1.152337151743309e-11
+    8.468410428611892e-11
+   -3.731925188734698e-13
+   -1.923688469579114e-12
+   -2.283024632694818e-11
+     8.07375645422932e-11
+ 6.58e+10    
+    8.065425610347383e-11
+   -2.282359676057825e-11
+    8.474777806431517e-11
+   -1.932473384874401e-12
+   -1.152880754830615e-11
+    8.468086360456525e-11
+   -3.688283896960323e-13
+   -1.922331945842668e-12
+   -2.283462626066106e-11
+    8.072628705622507e-11
+ 6.59e+10    
+    8.064317502095955e-11
+   -2.282810843208277e-11
+    8.474459197170822e-11
+   -1.931092929875277e-12
+   -1.153425101908328e-11
+    8.467760399009288e-11
+   -3.644628514412412e-13
+     -1.9209565167766e-12
+   -2.283899840636757e-11
+    8.071497977850016e-11
+ 6.6e+10     
+    8.063206453815449e-11
+   -2.283261245257157e-11
+    8.474138690347693e-11
+    -1.92969352595986e-12
+   -1.153970190107248e-11
+    8.467432540262587e-11
+    -3.60096057055392e-13
+    -1.91956218546072e-12
+   -2.284336268804169e-11
+    8.070364269187768e-11
+ 6.61e+10    
+    8.062092463768069e-11
+   -2.283710874572752e-11
+    8.473816281949473e-11
+   -1.928275176770047e-12
+   -1.154516016541425e-11
+    8.467102780226003e-11
+   -3.557281593270041e-13
+   -1.918148955369527e-12
+   -2.284771902990684e-11
+    8.069227577928389e-11
+ 6.62e+10    
+     8.06097553023242e-11
+   -2.284159723548004e-11
+    8.473491967980612e-11
+     -1.9268378863417e-12
+   -1.155062578308167e-11
+    8.466771114926309e-11
+   -3.513593108761682e-13
+   -1.916716830372887e-12
+   -2.285206735643703e-11
+    8.068087902381248e-11
+ 6.63e+10    
+    8.059855651503411e-11
+   -2.284607784600585e-11
+     8.47316574446259e-11
+   -1.925381659105228e-12
+   -1.155609872488021e-11
+    8.466437540407494e-11
+   -3.469896641439067e-13
+   -1.915265814736538e-12
+   -2.285640759235788e-11
+    8.066945240872356e-11
+ 6.64e+10    
+    8.058732825892214e-11
+   -2.285055050173031e-11
+    8.472837607433983e-11
+   -1.923906499886108e-12
+   -1.156157896144785e-11
+    8.466102052730734e-11
+   -3.426193713815612e-13
+   -1.913795913122767e-12
+   -2.286073966264796e-11
+    8.065799591744378e-11
+ 6.65e+10    
+    8.057607051726247e-11
+   -2.285501512732845e-11
+    8.472507552950404e-11
+   -1.922412413905467e-12
+   -1.156706646325498e-11
+    8.465764647974346e-11
+   -3.382485846402302e-13
+   -1.912307130590868e-12
+    -2.28650634925393e-11
+    8.064650953356516e-11
+ 6.66e+10    
+    8.056478327349095e-11
+     -2.2859471647726e-11
+    8.472175577084579e-11
+   -1.920899406780583e-12
+   -1.157256120060453e-11
+    8.465425322233924e-11
+   -3.338774557602025e-13
+   -1.910799472597761e-12
+   -2.286937900751914e-11
+     8.06349932408453e-11
+ 6.67e+10    
+    8.055346651120512e-11
+   -2.286391998810053e-11
+    8.471841675926266e-11
+   -1.919367484525393e-12
+   -1.157806314363181e-11
+    8.465084071622178e-11
+   -3.295061363604491e-13
+   -1.909272944998476e-12
+   -2.287368613333037e-11
+    8.062344702320678e-11
+ 6.68e+10    
+    8.054212021416344e-11
+   -2.286836007388233e-11
+    8.471505845582277e-11
+      -1.917816653551e-12
+   -1.158357226230463e-11
+    8.464740892269007e-11
+   -3.251347778281395e-13
+   -1.907727554046661e-12
+   -2.287798479597273e-11
+    8.061187086473647e-11
+ 6.69e+10    
+    8.053074436628486e-11
+   -2.287279183075552e-11
+    8.471168082176488e-11
+    -1.91624692066612e-12
+    -1.15890885264234e-11
+    8.464395780321534e-11
+   -3.207635313081899e-13
+   -1.906163306395049e-12
+   -2.288227492170393e-11
+    8.060026474968547e-11
+ 6.7e+10     
+    8.051933895164852e-11
+     -2.2877215184659e-11
+    8.470828381849853e-11
+   -1.914658293077516e-12
+   -1.159461190562107e-11
+    8.464048731943983e-11
+   -3.163925476928626e-13
+   -1.904580209095942e-12
+   -2.288655643704023e-11
+    8.058862866246829e-11
+ 6.71e+10    
+    8.050790395449353e-11
+   -2.288163006178743e-11
+    8.470486740760312e-11
+   -1.913050778390492e-12
+   -1.160014236936319e-11
+    8.463699743317781e-11
+   -3.120219776113682e-13
+    -1.90297826960166e-12
+   -2.289082926875771e-11
+    8.057696258766262e-11
+ 6.72e+10    
+    8.049643935921771e-11
+   -2.288603638859196e-11
+    8.470143155082848e-11
+   -1.911424384609239e-12
+   -1.160567988694799e-11
+    8.463348810641501e-11
+   -3.076519714195525e-13
+   -1.901357495764938e-12
+   -2.289509334389303e-11
+    8.056526651000908e-11
+ 6.73e+10    
+    8.048494515037832e-11
+   -2.289043409178153e-11
+    8.469797621009529e-11
+   -1.909779120137251e-12
+   -1.161122442750658e-11
+    8.462995930130847e-11
+   -3.032826791895872e-13
+    -1.89971789583938e-12
+   -2.289934858974423e-11
+    8.055354041441032e-11
+ 6.74e+10    
+    8.047342131269061e-11
+   -2.289482309832339e-11
+    8.469450134749347e-11
+   -1.908114993777723e-12
+   -1.161677596000277e-11
+    8.462641098018672e-11
+   -2.989142506997243e-13
+   -1.898059478479762e-12
+   -2.290359493387174e-11
+    8.054178428593092e-11
+ 6.75e+10    
+    8.046186783102805e-11
+   -2.289920333544415e-11
+    8.469100692528372e-11
+   -1.906432014733853e-12
+    -1.16223344532335e-11
+    8.462284310554934e-11
+   -2.945468354240863e-13
+   -1.896382252742495e-12
+   -2.290783230409907e-11
+    8.052999810979671e-11
+ 6.76e+10    
+    8.045028469042145e-11
+   -2.290357473063059e-11
+    8.468749290589634e-11
+   -1.904730192609222e-12
+   -1.162789987582866e-11
+    8.461925564006723e-11
+    -2.90180582522489e-13
+   -1.894686228085906e-12
+   -2.291206062851376e-11
+    8.051818187139467e-11
+ 6.77e+10    
+    8.043867187605889e-11
+   -2.290793721163044e-11
+    8.468395925193147e-11
+   -1.903009537408098e-12
+   -1.163347219625137e-11
+    8.461564854658223e-11
+   -2.858156408303385e-13
+   -1.892971414370566e-12
+   -2.291627983546809e-11
+    8.050633555627215e-11
+ 6.78e+10    
+    8.042702937328513e-11
+   -2.291229070645329e-11
+    8.468040592615889e-11
+   -1.901270059535701e-12
+   -1.163905138279802e-11
+     8.46120217881067e-11
+   -2.814521588485544e-13
+   -1.891237821859634e-12
+   -2.292048985357977e-11
+    8.049445915013653e-11
+ 6.79e+10    
+    8.041535716760093e-11
+   -2.291663514337123e-11
+    8.467683289151798e-11
+   -1.899511769798519e-12
+   -1.164463740359851e-11
+    8.460837532782402e-11
+   -2.770902847335361e-13
+   -1.889485461219101e-12
+   -2.292469061173291e-11
+    8.048255263885487e-11
+ 6.8e+10     
+    8.040365524466312e-11
+   -2.292097045091975e-11
+    8.467324011111742e-11
+   -1.897734679404517e-12
+    -1.16502302266163e-11
+    8.460470912908806e-11
+   -2.727301662872166e-13
+   -1.887714343518064e-12
+   -2.292888203907849e-11
+     8.04706160084533e-11
+ 6.81e+10    
+    8.039192359028363e-11
+   -2.292529655789827e-11
+     8.46696275482352e-11
+   -1.895938799963421e-12
+    -1.16558298196486e-11
+    8.460102315542269e-11
+     -2.6837195094711e-13
+   -1.885924480228995e-12
+   -2.293306406503521e-11
+    8.045864924511684e-11
+ 6.82e+10    
+    8.038016219042953e-11
+   -2.292961339337117e-11
+    8.466599516631835e-11
+   -1.894124143486871e-12
+   -1.166143615032664e-11
+    8.459731737052257e-11
+   -2.640157857764656e-13
+   -1.884115883227919e-12
+   -2.293723661929026e-11
+    8.044665233518847e-11
+ 6.83e+10    
+    8.036837103122225e-11
+   -2.293392088666819e-11
+    8.466234292898261e-11
+   -1.892290722388666e-12
+   -1.166704918611568e-11
+    8.459359173825182e-11
+   -2.596618174544483e-13
+   -1.882288564794627e-12
+   -2.294139963179968e-11
+    8.043462526516935e-11
+ 6.84e+10    
+    8.035655009893736e-11
+   -2.293821896738526e-11
+    8.465867080001259e-11
+   -1.890438549484897e-12
+   -1.167266889431529e-11
+    8.458984622264456e-11
+   -2.553101922663806e-13
+   -1.880442537612896e-12
+   -2.294555303278937e-11
+    8.042256802171789e-11
+ 6.85e+10    
+    8.034469938000416e-11
+   -2.294250756538519e-11
+    8.465497874336145e-11
+   -1.888567637994116e-12
+   -1.167829524205962e-11
+    8.458608078790472e-11
+   -2.509610560940418e-13
+   -1.878577814770576e-12
+   -2.294969675275548e-11
+    8.041048059164939e-11
+ 6.86e+10    
+    8.033281886100481e-11
+    -2.29467866107981e-11
+    8.465126672315022e-11
+   -1.886678001537466e-12
+   -1.168392819631745e-11
+    8.458229539840542e-11
+   -2.466145544060243e-13
+   -1.876694409759775e-12
+   -2.295383072246503e-11
+    8.039836296193564e-11
+ 6.87e+10    
+    8.032090852867443e-11
+   -2.295105603402226e-11
+    8.464753470366861e-11
+   -1.884769654138749e-12
+   -1.168956772389258e-11
+     8.45784900186887e-11
+    -2.42270832248151e-13
+   -1.874792336476974e-12
+   -2.295795487295652e-11
+    8.038621511970467e-11
+ 6.88e+10    
+    8.030896836990071e-11
+   -2.295531576572464e-11
+    8.464378264937367e-11
+   -1.882842610224565e-12
+   -1.169521379142397e-11
+    8.457466461346617e-11
+    -2.37930034233962e-13
+   -1.872871609223069e-12
+   -2.296206913554058e-11
+    8.037403705223987e-11
+ 6.89e+10    
+     8.02969983717229e-11
+   -2.295956573684142e-11
+    8.464001052489054e-11
+   -1.880896884624341e-12
+   -1.170086636538601e-11
+    8.457081914761772e-11
+   -2.335923045352301e-13
+   -1.870932242703511e-12
+   -2.296617344180044e-11
+    8.036182874698005e-11
+ 6.9e+10     
+    8.028499852133184e-11
+    -2.29638058785785e-11
+    8.463621829501139e-11
+   -1.878932492570385e-12
+   -1.170652541208875e-11
+    8.456695358619179e-11
+   -2.292577868725894e-13
+   -1.868974252028305e-12
+   -2.297026772359228e-11
+     8.03495901915186e-11
+ 6.91e+10    
+    8.027296880606939e-11
+   -2.296803612241217e-11
+    8.463240592469573e-11
+   -1.876949449697881e-12
+   -1.171219089767823e-11
+    8.456306789440513e-11
+   -2.249266245061908e-13
+    -1.86699765271204e-12
+    -2.29743519130461e-11
+    8.033732137360332e-11
+ 6.92e+10    
+    8.026090921342816e-11
+   -2.297225640008955e-11
+    8.462857337906982e-11
+   -1.874947772044938e-12
+   -1.171786278813661e-11
+    8.455916203764227e-11
+   -2.205989602264383e-13
+   -1.865002460673913e-12
+   -2.297842594256586e-11
+    8.032502228113593e-11
+ 6.93e+10    
+    8.024881973105082e-11
+   -2.297646664362911e-11
+    8.462472062342679e-11
+   -1.872927476052505e-12
+   -1.172354104928271e-11
+    8.455523598145569e-11
+   -2.162749363447762e-13
+   -1.862988692237695e-12
+   -2.298248974483012e-11
+    8.031269290217142e-11
+ 6.94e+10    
+    8.023670034672996e-11
+   -2.298066678532121e-11
+    8.462084762322608e-11
+   -1.870888578564374e-12
+   -1.172922564677207e-11
+    8.455128969156528e-11
+   -2.119546946845689e-13
+   -1.860956364131685e-12
+   -2.298654325279248e-11
+    8.030033322491778e-11
+ 6.95e+10    
+    8.022455104840738e-11
+   -2.298485675772831e-11
+    8.461695434409312e-11
+   -1.868831096827069e-12
+   -1.173491654609732e-11
+    8.454732313385779e-11
+   -2.076383765720476e-13
+   -1.858905493488657e-12
+   -2.299058639968192e-11
+    8.028794323773578e-11
+ 6.96e+10    
+    8.021237182417388e-11
+   -2.298903649368575e-11
+    8.461304075181912e-11
+   -1.866755048489784e-12
+   -1.174061371258856e-11
+    8.454333627438699e-11
+   -2.033261228272878e-13
+   -1.856836097845765e-12
+   -2.299461911900327e-11
+    8.027552292913806e-11
+ 6.97e+10    
+    8.020016266226881e-11
+   -2.299320592630196e-11
+    8.460910681236125e-11
+   -1.864660451604256e-12
+   -1.174631711141367e-11
+    8.453932907937332e-11
+   -1.990180737553153e-13
+   -1.854748195144431e-12
+   -2.299864134453755e-11
+     8.02630722877891e-11
+ 6.98e+10    
+    8.018792355107947e-11
+   -2.299736498895888e-11
+    8.460515249184133e-11
+    -1.86254732462463e-12
+    -1.17520267075786e-11
+    8.453530151520344e-11
+   -1.947143691372381e-13
+   -1.852641803730216e-12
+   -2.300265301034245e-11
+    8.025059130250456e-11
+ 6.99e+10    
+    8.017565447914111e-11
+   -2.300151361531245e-11
+     8.46011777565466e-11
+   -1.860415686407278e-12
+   -1.175774246592774e-11
+    8.453125354842964e-11
+   -1.904151482214885e-13
+   -1.850516942352675e-12
+    -2.30066540507525e-11
+    8.023807996225116e-11
+ 7e+10       
+    8.016335543513601e-11
+   -2.300565173929285e-11
+    8.459718257292866e-11
+   -1.858265556210685e-12
+   -1.176346435114431e-11
+    8.452718514577025e-11
+    -1.86120549715101e-13
+    -1.84837363016514e-12
+   -2.301064440037953e-11
+    8.022553825614561e-11
* NOTE: Solution at 1e+08 Hz used as DC point.

.ends
