* begin ansoft header
* node 1 Diff1
* node 2 Comm1
* node 3 trace_p_1_T1
* node 4 trace_n_1_T1
* node 5 Diff2
* node 6 Comm2
* node 7 trace_p_1_T2
* node 8 trace_n_1_T2
* 
* created by ElectronicsDesktop
* end ansoft header

.subckt m4lines_port_lfws 1 2 3 4 5 6 7 8 
v2_1 2 9 dc 0.0
v2_3 2 10 dc 0.0
v2_4 2 11 dc 0.0
v3_1 3 12 dc 0.0
v3_4 3 13 dc 0.0
v4_1 4 14 dc 0.0
v6_5 6 15 dc 0.0
v6_7 6 16 dc 0.0
v6_8 6 17 dc 0.0
v7_5 7 18 dc 0.0
v7_8 7 19 dc 0.0
v8_5 8 20 dc 0.0
v1_0 1 21 dc 0.0
v2_0 2 22 dc 0.0
v3_0 3 23 dc 0.0
v4_0 4 24 dc 0.0
v5_0 5 25 dc 0.0
v6_0 6 26 dc 0.0
v7_0 7 27 dc 0.0
v8_0 8 28 dc 0.0
rl1_2to1 9 29 63.840555156694
ls1_2to1 29 1 0.0039817286430045n
rl1_2to3 10 30 4.6110165069357
ls1_2to3 30 3 0.010347696898797n
rl1_2to4 11 31 10.980365682825
ls1_2to4 31 4 0.015834478529838n
rl1_3to1 12 32 71.029832734281
ls1_3to1 32 1 0.032344772398123n
rl1_3to4 13 33 21.918881392921
ls1_3to4 33 4 0.047837679150717n
rl1_4to1 14 34 70.245712711744
ls1_4to1 34 1 0.02792988676232n
rl1_6to5 15 35 63.910326686112
ls1_6to5 35 5 0.0046113552910051n
rl1_6to7 16 36 4.6095498034104
ls1_6to7 36 7 0.0104091815262n
rl1_6to8 17 37 10.984660840354
ls1_6to8 37 8 0.01575314083167n
rl1_7to5 18 38 71.066004608921
ls1_7to5 38 5 0.032189049651494n
rl1_7to8 19 39 21.895535092654
ls1_7to8 39 8 0.048261494762328n
rl1_8to5 20 40 70.277075493273
ls1_8to5 40 5 0.027683863205787n
rl1_1to0 21 41 96.70390194301
ls1_1to0 41 0 0.086231140000151n
rl1_2to0 22 42 116.48598502572
ls1_2to0 42 0 0.13977429101775n
rl1_3to0 23 43 96.675385796509
ls1_3to0 43 0 0.086833071581642n
rl1_4to0 24 44 116.56169447299
ls1_4to0 44 0 0.13920231528253n
rl1_5to0 25 45 96.416803617011
ls1_5to0 45 0 0.085231332293128n
rl1_6to0 26 46 116.63154652472
ls1_6to0 46 0 0.14110223216126n
rl1_7to0 27 47 96.690248191268
ls1_7to0 47 0 0.087110252334829n
rl1_8to0 28 48 116.549838167
ls1_8to0 48 0 0.138626684157n
.ends m4lines_port_lfws

