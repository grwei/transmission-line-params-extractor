* BEGIN ANSOFT HEADER
* node 1    1:trace_p_0_T1_A
* node 2    1:trace_n_0_T1_A
* node 3    1:trace_n_1_T1_A
* node 4    1:trace_p_1_T1_A
* node 5    Ground_A
* node 6    1:trace_p_0_T1_B
* node 7    1:trace_n_0_T1_B
* node 8    1:trace_n_1_T1_B
* node 9    1:trace_p_1_T1_B
* node 10   Ground_B
*  Project: 4lines
*   Design: 2-diff-pairs
*   Length: 5
*   Format: HSPICE
*  Creator: Ansoft HFSS
*     Date: Sat Jun 06 10:16:34 2020
* END ANSOFT HEADER

.subckt ckt_m4lines_HFSS_W 1 2 3 4 inref 5 6 7 8 outref length=5.08M

.model m4lines_HFSS_W_1 W MODELTYPE=table N=4 RMODEL=r_m4lines_HFSS_W_1
+ LMODEL=l_m4lines_HFSS_W_1 GMODEL=g_m4lines_HFSS_W_1 CMODEL=c_m4lines_HFSS_W_1

* Example usage:
W1 1 2 3 4 inref 5 6 7 8 outref N=4 L=length TABLEMODEL=m4lines_HFSS_W_1

.model r_m4lines_HFSS_W_1 sp N=4 SPACING=nonuniform VALTYPE=real
+ INTERPOLATION=spline
+ DATA = 700
+ 0           
+        6.906563104539061
+       0.6824161915317021
+        7.004584896377449
+       0.2837910405679777
+       0.9085696485041762
+        7.004887839056049
+       0.1145299239677343
+       0.2838404372629029
+       0.6766741287148066
+        6.856349044729821
+ 2e+08       
+        10.30113018179325
+        1.016369991615166
+        10.42632538041021
+       0.4018314087202817
+        1.334554596554753
+        10.41166364888455
+       0.1591891771844975
+       0.4037052692906891
+       0.9956869977619988
+        10.18231608077756
+ 3e+08       
+        12.64693105855384
+        1.143445082924333
+        12.80083132398006
+       0.4676939192679698
+         1.61106569253252
+         12.7762878231201
+       0.1753503940366344
+       0.4722341824890993
+        1.128844953370267
+        12.46352802132555
+ 4e+08       
+        14.63939197932881
+        1.258953351911071
+        14.82210135968447
+       0.5156127722746302
+        1.846192710895932
+          14.787841859159
+        0.181877090736275
+         0.52253867378994
+        1.249142618813348
+        14.39228693024461
+ 5e+08       
+        16.47200157222983
+        1.384934013041704
+        16.67790545488358
+       0.5602022126706039
+         2.06378850362835
+        16.63424818619715
+       0.1888717287836398
+       0.5693786520762407
+        1.377373107058749
+         16.1634982631831
+ 6e+08       
+        18.17011827891403
+        1.505648952327599
+        18.39373979737844
+       0.6034369240157705
+        2.264998191080702
+        18.34147658651015
+       0.1975974737755371
+       0.6147865607558634
+        1.498931333523312
+        17.80301996088844
+ 7e+08       
+        19.73880326064288
+        1.612446501113803
+        19.97721181134416
+       0.6444640535755874
+        2.449893571943583
+        19.91722839205754
+       0.2069202905547622
+       0.6578909896267338
+         1.60593246301257
+        19.31551094799766
+ 8e+08       
+        21.19426812974825
+        1.706646351512395
+        21.44648842603627
+       0.6826178836295976
+        2.620744225052114
+        21.37958398469257
+        0.215746200272815
+       0.6980109576400029
+        1.700104153249248
+        20.71677202728548
+ 9e+08       
+        22.56356240548607
+        1.795012715869257
+        22.82888586693532
+       0.7179645651863509
+        2.781310092291281
+        22.75579286350476
+       0.2235815349106163
+       0.7352228720687354
+        1.788452779992685
+        22.03380519838202
+ 1e+09       
+         23.8787626072638
+        1.885970198019283
+        24.15519908538059
+       0.7511468146685966
+         2.93583252969783
+        24.07668354204158
+       0.2304596376260809
+       0.7701990279719761
+        1.879579575967833
+        23.29895651296864
+ 1.1e+09     
+        25.13360880680375
+        1.877247010669332
+        25.46015527882673
+       0.7006177817879486
+        3.071174545045083
+        25.37228517375954
+       0.1334815764463078
+       0.7164888255646643
+        1.865935141681817
+        24.48271534323289
+ 1.2e+09     
+          26.413802348726
+        1.917487571151088
+        26.78689155250182
+       0.6668742201136855
+        3.219228316629543
+        26.69002914977433
+      0.04085201756988904
+       0.6794232458096092
+        1.901114284232534
+        25.69262154349731
+ 1.3e+09     
+        27.70271178711088
+        1.995196694252474
+        28.11765985622207
+       0.6471989628528618
+        3.374020354572104
+        28.01229814123893
+     -0.04712763676555201
+       0.6564618393272081
+        1.973735321480377
+         26.9128766354176
+ 1.4e+09     
+         28.9862346561308
+        2.099994894815049
+        29.43766272211967
+       0.6390142536543031
+        3.530819532168033
+        29.32439307246827
+      -0.1301951135517385
+       0.6451561542077671
+        2.073522409669733
+        28.13001365416687
+ 1.5e+09     
+        30.25281907502116
+        2.222936849738949
+        30.73500525899849
+       0.6400050534597476
+        3.685947702940206
+        30.61448642188762
+      -0.2080970837669806
+       0.6432802342447754
+        2.191617934300631
+        29.33293507213535
+ 1.6e+09     
+        31.49334226940813
+        2.356585581118154
+        32.00050606916199
+       0.6481722346137162
+        3.836620953849006
+        31.87343612684141
+      -0.2805803050132432
+       0.6488921226099735
+        2.320654341145846
+        30.51281371744576
+ 1.7e+09     
+        32.70090070723933
+        2.494948083667501
+        33.22742390325894
+       0.6618417113592565
+         3.98081178650944
+        33.09451622322792
+       -0.347394208006092
+       0.6603507341567383
+        2.454689936810639
+        31.66290801824352
+ 1.8e+09     
+        33.87055317896288
+        2.633339875165639
+        34.41114331088961
+       0.6796479618456754
+        4.117127671504956
+        34.27310688523927
+      -0.4082985495883609
+       0.6763058910640306
+        2.589075112619156
+        32.77833036634153
+ 1.9e+09     
+        34.99904663387917
+        2.768219794962333
+        35.54885042424731
+       0.7005042622187286
+        4.244703894688388
+        35.40637455769421
+      -0.4630723215640521
+       0.6956737207681857
+        2.720289554020939
+        33.85579668899106
+ 2e+09       
+        36.08454519537862
+        2.897019330257495
+        36.63921991421584
+       0.7235674603330687
+        4.363109608820293
+        36.49296292595743
+      -0.5115218439454163
+       0.7176053664001651
+         2.84577420083148
+        34.89337662603143
+ 2.1e+09     
+        37.12637543382786
+        3.017979966772407
+        37.68212618130569
+       0.7482020125610711
+        4.472266274306121
+        37.53270761943923
+      -0.5534870826462486
+       0.7414539408031684
+        2.963771138799809
+        35.89025691005155
+ 2.2e+09     
+        38.12479544801801
+         3.13000539082003
+        38.67838583863032
+       0.7739459483816847
+        4.572377642037408
+        38.52638163691456
+      -0.5888459019120804
+       0.7667426039372701
+        3.073178076992598
+        36.84652540924064
+ 2.3e+09     
+        39.08079131014955
+        3.232531338474817
+        39.62953424167434
+       0.8004801076416036
+        4.663870315927253
+        39.47547424693791
+      -0.6175163372374983
+        0.793135298867383
+        3.173420130957934
+        37.76297955121164
+ 2.4e+09     
+        39.99590167191469
+        3.325413525827225
+        40.53763590662891
+       0.8276011782931839
+        4.747343831252056
+        40.38200324586258
+      -0.6394571610084819
+       0.8204108299973468
+        3.264339330800465
+        38.64096023536927
+ 2.5e+09     
+        40.87206953459171
+        3.408832778762414
+        41.40512682560642
+       0.8551985780058389
+        4.823529132741053
+        41.24835864534101
+       -0.654667083635071
+       0.8484404490690942
+        3.346100992980974
+        39.48221061399997
+ 2.6e+09     
+        41.71151911150566
+         3.48321581323818
+        42.23468565434798
+       0.8832349536853334
+        4.893254337556324
+        42.07717483753759
+      -0.6631829362350669
+       0.8771688160199744
+        3.419115445074411
+        40.28875806073339
+ 2.7e+09     
+        42.51665515414317
+        3.549169844048279
+        43.02913028190433
+       0.9117299392270277
+        4.957416713452966
+        42.87122782017345
+      -0.6650771485575796
+       0.9065980446143136
+        3.483973326518623
+        41.06281706712924
+ 2.8e+09     
+        43.28998191204465
+        3.607429160254141
+        43.79133620593243
+       0.9407467611622353
+        5.016959878018944
+        43.63335397228684
+      -0.6604547875686956
+       0.9367744738449049
+        3.541392648696744
+        41.80671056751079
+ 2.9e+09     
+        44.03403892757394
+        3.658811896694104
+        44.52417329034031
+       0.9703812799279194
+        5.072855317999452
+        44.36638701651808
+      -0.6494503698101377
+        0.967777790303923
+        3.592175885383869
+        42.52280717568101
+ 3e+09       
+        44.75135103857981
+        3.704185389183002
+        45.23045777140442
+        1.000753079320065
+        5.126087427739868
+        45.07311008393909
+      -0.6322246109309559
+       0.9997121411823455
+        3.637175517546796
+        43.21347194054515
+ 3.1e+09     
+        45.44439021011045
+        3.744438686742028
+        45.91291673283791
+        1.031998254499914
+        5.177641365007231
+        45.75622014273956
+      -0.6089612319983669
+        1.032698907695593
+        3.677266636471536
+        43.88102843034645
+ 3.2e+09     
+        46.11554709667823
+        3.780460983910714
+        46.57416264244353
+        1.064263591324635
+        5.228493115785835
+        46.41830241591978
+      -0.5798639055774912
+        1.066870845511535
+        3.713325393358125
+        44.52773019529499
+ 3.3e+09     
+        46.76711052050116
+         3.81312491655735
+        47.21667590356453
+        1.097701871889921
+        5.279601244157071
+        47.06181276646844
+       -0.545153395187145
+        1.102367336777762
+        3.746212258896708
+        45.15573990807333
+ 3.4e+09     
+        47.40125332129512
+        3.843273828783185
+        47.84279370684968
+        1.132468080366861
+        5.331899877786682
+        47.68906635469657
+      -0.5050649189939536
+        1.139330534578318
+        3.776759216225821
+        45.76711472363277
+ 3.5e+09     
+        48.02002327994694
+        3.871712263692831
+        48.45470376375133
+        1.168716318266369
+        5.386292543765577
+        48.30223116332631
+      -0.4598457516022048
+        1.177902213573722
+        3.805760152287155
+        46.36379662380951
+ 3.6e+09     
+        48.62533803745464
+        3.899199056594089
+        49.05444176022541
+        1.206597268814421
+        5.443646524334284
+        48.90332523900577
+      -0.4097530655452846
+        1.218221169611476
+        3.833963835491157
+        46.94760671355224
+ 3.7e+09     
+        49.21898312089475
+         3.92644251658192
+        49.64389158826501
+        1.246256076330699
+        5.504787448697839
+        49.49421671499612
+      -0.3550520056299893
+        1.260421036232305
+        3.862068972707726
+        47.52024261224865
+ 3.8e+09     
+        49.80261235098857
+        3.954097273162087
+        50.22478759716299
+         1.28783052882599
+        5.570493877455497
+        50.07662586167979
+      -0.2960139837633213
+        1.304628407572463
+        3.890720927511543
+        48.08327823612194
+ 3.9e+09     
+        50.37775004329847
+        3.982762440583069
+        50.79871825971519
+        1.331449451087649
+        5.641491672195523
+        50.65212856309338
+      -0.2329151785556047
+        1.350961175701608
+        3.920509756254148
+        48.63816539749394
+ 4e+09       
+        50.94579452998509
+        4.012980815928439
+        51.36713077526623
+        1.377231232004953
+        5.718447976872666
+        51.22216074309418
+      -0.1660352222153378
+        1.399527006572316
+        3.951969280885713
+        49.18623675606938
+ 4.1e+09     
+        51.50802262428559
+        4.045238879743968
+        51.93133623586157
+        1.425282424535093
+        5.801964672278301
+        51.78802336821313
+     -0.09565605651215758
+        1.450421893180332
+        3.985576969402753
+        49.72870974872514
+ 4.2e+09     
+        52.06559472829911
+        4.079967411840163
+        52.49251506784654
+        1.475696370276152
+        5.892571203037121
+        52.35088773969727
+     -0.02206093946251131
+        1.503728737959958
+        4.021754438103826
+        50.26669120000732
+ 4.3e+09     
+        52.61956034887759
+        4.117542571540989
+          53.051722532765
+        1.528551813842085
+        5.990716721111709
+        52.91180085833434
+      0.05446641545458153
+          1.5595159295887
+        4.060868426061614
+        50.80118237797789
+ 4.4e+09     
+         53.1708638387851
+        4.158287322454957
+        53.60989413164597
+         1.58391148585273
+        6.096761543847857
+        53.47169070563288
+        0.133642585591065
+         1.61783589295692
+        4.103232122745124
+        51.33308431129314
+ 4.5e+09     
+        53.72035022285134
+        4.202473108051674
+        54.16785080861822
+        1.641820648034076
+        6.210967991137725
+        54.03137133663432
+       0.2151850890365952
+        1.678723605734383
+        4.149106755740776
+        51.86320322531001
+ 4.6e+09     
+        54.26877100336303
+        4.250321706960971
+        54.72630389569141
+        1.702305610251364
+        6.333490747910153
+        54.59154772547262
+       0.2988129566890638
+        1.742195091308372
+        4.198703368032485
+        52.39225598921487
+ 4.7e+09     
+        54.81678986690136
+        4.302007216814584
+        55.28585978244726
+        1.765372247685654
+        6.464366996623367
+        55.15282034668343
+       0.3842472459781272
+        1.808245916285951
+        4.252184734129894
+        52.92087549404097
+ 4.8e+09     
+        55.36498823747494
+        4.357658133263372
+        55.84702433368611
+        1.831004566967411
+        6.603506679992184
+        55.71568951460711
+       0.4712115172093507
+        1.876849741396468
+        4.309667382110382
+        53.44961590412932
+ 4.9e+09     
+        55.91387063912534
+        4.417359506954501
+        56.41020711555567
+        1.899163392662827
+        6.750683384784341
+        56.28055954074964
+       0.5594322954845294
+        1.947956997259803
+        4.371223704779713
+        53.97895774305275
+ 5e+09       
+        56.46386984598216
+        4.481155175932922
+           56.97572552631
+        1.969785269297949
+        6.905526477865711
+        56.84774280465894
+       0.6486395435242955
+        2.021493780326905
+        4.436884157844935
+         54.5093127900176
+ 5.1e+09     
+        57.01535180963184
+        4.549050084065412
+        57.54380896071604
+        2.042781697639141
+        7.067515266223199
+        57.41746386680833
+       0.7385671732287635
+         2.09736108788602
+        4.506639556146861
+        55.04102877484839
+ 5.2e+09     
+        57.56862036305395
+        4.621012707308225
+        58.11460316529986
+        2.118038844946571
+        7.235976078864236
+        57.98986378022911
+       0.8289536260788943
+        2.175434532079142
+        4.580443490251724
+        55.57439386927101
+ 5.3e+09     
+        58.12392170754696
+        4.696977618296096
+        58.68817496214027
+        2.195417884236734
+        7.410083260332271
+        58.56500477821708
+       0.9195425539846749
+        2.255564688241972
+        4.658214894394116
+          56.109640979586
+ 5.4e+09     
+        58.68144869415089
+         4.77684822490769
+        59.26451752787855
+        2.274756123309101
+         7.58886509831535
+        59.14287552447221
+        1.010083632277152
+        2.337578238643423
+        4.739840801978947
+        56.64695185110278
+ 5.5e+09     
+        59.24134491410202
+        4.860499719081026
+        59.84355640753864
+        2.355869076016511
+        7.771215653724818
+        59.72339710501554
+        1.100333534495925
+        2.421280064458819
+        4.825179325509017
+        57.18646099791028
+ 5.6e+09     
+        59.80370861381904
+        4.947782267122491
+        60.42515641519265
+        2.438553601679951
+        7.955913293517154
+         60.3064299137366
+        1.190057093732077
+        2.506456412254103
+        4.914062892817128
+        57.72825947268396
+ 5.7e+09     
+        60.36859644880447
+        5.038524461234284
+        61.00912952199447
+        2.522592190297495
+          8.1416464231296
+        60.89178153196716
+        1.279028666993115
+        2.592879213013484
+        5.006301760001036
+        58.27239849024892
+ 5.8e+09     
+        60.93602708772821
+        5.132537033662937
+        61.59524375529033
+        2.607758399915551
+        8.327046468018747
+        61.47921562571933
+        1.367033707130734
+        2.680311560452954
+        5.101687803178343
+        58.81889291562539
+ 5.9e+09     
+         61.5059846730786
+        5.229616810306308
+        62.18323303243351
+          2.6938233600138
+        8.510727573492941
+        62.06846178420171
+        1.453870531596154
+         2.76851426282041
+        5.199998566647717
+        59.36772462250205
+ 6e+09       
+        62.07842213857897
+        5.329550851489643
+        62.77280773601302
+        2.780563146876943
+         8.69133181547047
+        62.65922610635526
+        1.539352259601943
+        2.857253274469476
+        5.301001515950118
+        59.91884572198492
+ 6.1e+09     
+        62.65326437678969
+        5.432120696843685
+        63.36366571465815
+         2.86776672401219
+        8.867578006538908
+        63.25120221965143
+        1.623308870834883
+        2.946307700538992
+        5.404458413575535
+        60.47218165476411
+ 6.2e+09     
+        63.23041124387496
+        5.537106602789719
+         63.9555032808289
+        2.955244036942165
+        9.038311530779382
+         63.8440823026818
+        1.705589321972236
+        3.035477964304357
+        5.510129706658697
+          61.027634133467
+ 6.3e+09     
+        63.80974038348465
+        5.644291639673813
+        64.54802569185314
+        3.042833773602387
+        9.202552150292171
+        64.43756759795635
+        1.786063644552039
+        3.124593648644296
+        5.617778794565801
+        61.58508391698311
+ 6.4e+09     
+        64.39110984907195
+        5.753465505563049
+        65.14095656018414
+        3.130410265016923
+        9.359536496045065
+         65.0313778610634
+        1.864624941800137
+        3.213520486514052
+        5.727176034263078
+        62.14439339597316
+ 6.5e+09     
+        64.97436050454836
+        5.864427918512837
+        65.73404565643035
+        3.217889017926838
+        9.508752061004916
+        65.62525920993781
+        1.941191204753265
+        3.302165992352966
+         5.83810234616625
+        62.70540896938503
+ 6.6e+09     
+        65.55931818725729
+        5.976991470127565
+        66.32707464948153
+        3.305230446475051
+        9.649959985267046
+        66.21898991876755
+        2.015706880215629
+        3.390483301855109
+        5.950352304193172
+        63.26796319592071
+ 6.7e+09     
+        66.14579562461496
+        6.090983859278855
+        66.91986046727006
+        3.392441499489436
+        9.783204733637856
+        66.81238384027495
+        2.088144144022805
+        3.478472917075141
+         6.06373662978603
+        63.83187671179262
+ 6.8e+09     
+         66.7335941055662
+         6.20624947205278
+        67.51225614431199
+         3.47957504939032
+        9.908809828574579
+        67.40529132271111
+        2.158503860496738
+        3.566182223454015
+        6.178084056876934
+        64.39695991593521
+ 6.9e+09     
+        67.32250491894779
+        6.322650326393272
+        68.10414922490597
+        3.566727096741766
+        10.02735998074077
+        67.99759769061197
+        2.226816239374393
+        3.653702833480851
+        6.293242587156711
+         64.9630144348028
+ 7e+09       
+        67.91231058140002
+        6.440066450472162
+        68.69545798649382
+        3.654032025755576
+         10.1396710977257
+        68.58921955398222
+        2.293141230803429
+        3.741165993126533
+        6.409080205559022
+        65.52983438945579
+ 7.1e+09     
+        68.50278588616652
+        6.558395805852879
+        69.28612591022127
+        3.741656296616448
+        10.24675059806631
+         69.1800993730824
+        2.357568723339221
+        3.828736437848539
+        6.525485167882051
+        66.09720749634049
+ 7.2e+09     
+        69.09369880984426
+        6.677553894919234
+        69.87611493544114
+        3.829791062069507
+          10.349751098004
+        69.77019881568515
+        2.420218626302572
+        3.916605186606772
+         6.64236600084495
+        66.66491603890762
+ 7.3e+09     
+        69.68481131633062
+        6.797473204179948
+         70.4653980815975
+        3.918644238912828
+        10.44992081334903
+        70.35949149035442
+        2.481240924852573
+        4.004981805551772
+        6.759651366972693
+        67.23273774938991
+ 7.4e+09     
+        70.27588009586867
+        6.918102631036625
+        71.05395200506922
+        4.008432550298189
+        10.54855393085806
+        70.94795562342372
+        2.540815793769219
+        4.094086658281377
+        6.877289942624181
+        67.80044663871719
+ 7.5e+09     
+         70.8666572727815
+        7.039407023905529
+        71.64174998984416
+        4.099373991075866
+        10.64694380890907
+        71.53556717864241
+        2.599153845683778
+        4.184143595824546
+        6.995250439716355
+        68.36781380821661
+ 7.6e+09     
+        71.45689110909069
+        7.161366938326259
+        72.22875576529309
+        4.191681070587211
+        10.74634125835885
+        72.12229381284503
+        2.656496573728468
+        4.275373441574557
+        7.113521874358121
+        68.93460827034144
+ 7.7e+09     
+         72.0463267237979
+        7.283978679606379
+        72.81491842020692
+        4.285555072337454
+        10.84791943790803
+        72.70808993688492
+        2.713117030051279
+        4.367988511291768
+        7.232114153429755
+        69.50059779822308
+ 7.8e+09     
+        72.63470684012356
+        7.407254670120267
+        73.40016855698562
+         4.38118145391231
+         10.9527461746304
+        73.29289302578792
+        2.769320762945688
+        4.462188292080153
+        7.351059017604669
+        70.06554981633292
+ 7.9e+09     
+        73.22177256624931
+        7.531224150159904
+        73.98441571720498
+         4.47872640606742
+        11.06176386939348
+        73.87662120939979
+        2.825447018532961
+        4.558156299649294
+        7.470411349965576
+        70.62923233775672
+ 8e+09       
+        73.80726420958982
+        7.655934197535881
+         74.5675470186552
+        4.578334505377751
+         11.1757766205697
+        74.45917208364469
+        2.881870199336718
+        4.656058048467894
+         7.59025083552934
+        71.19141494802284
+ 8.1e+09     
+        74.39092212055897
+        7.781451033999883
+        75.14942687838982
+        4.680127333910271
+        11.29544382116841
+        75.04042261693267
+        2.939001562303194
+        4.756040008319754
+        7.710683939712489
+        71.75186983132244
+ 8.2e+09     
+        74.97248755919527
+        7.907861575992102
+        75.72989765625924
+         4.78420290199026
+        11.42127925385749
+         75.6202299861488
+        2.997291132828575
+        4.858229383202616
+        7.831846163032512
+         72.3103728323028
+ 8.3e+09     
+        75.55170357669934
+        8.035275182441985
+          76.308781035826
+        4.890635693494469
+        11.55365460797918
+        76.19843315903724
+        3.057229808705342
+        4.962734531682152
+        7.953904524374335
+         72.8667045452558
+ 8.4e+09     
+        76.12831590364554
+        8.163825552179752
+        76.88587995986374
+        4.999477152953943
+        11.69280634587727
+        76.77485504005662
+        3.119351627900215
+        5.069645847455179
+          8.0770602247811
+        73.42065142215927
+ 8.5e+09     
+        76.70207383708625
+        8.293672726638803
+        77.46098095069399
+        5.110756445340233
+        11.83884492292312
+        77.34930500977791
+        3.184236175958593
+        5.179036930238052
+        8.201551446624803
+        73.97200689142616
+ 8.6e+09     
+        77.27273111967851
+        8.425005158686325
+        78.03385666657367
+        5.224481338266691
+        11.99176548849131
+        77.92158170879813
+        3.252511111869653
+        5.290965895695326
+        8.327656247933183
+         74.5205724800426
+ 8.7e+09     
+        77.84004680510701
+        8.558041814568346
+        78.60426857012645
+        5.340639078693949
+        12.15145934014154
+        78.49147594186809
+        3.324854794812701
+        5.405476695192314
+        8.455695517539667
+        75.06615893284288
+ 8.8e+09     
+        78.40378610527971
+         8.69303428229002
+        79.17196961030933
+        5.459197159215966
+        12.31772555236504
+        79.05877360335815
+         3.40199899787449
+        5.522600338816494
+        8.586035962784718
+        75.60858732378034
+ 8.9e+09     
+        78.96372121590132
+        8.830268865717168
+        79.73670684346095
+          5.5801038906477
+        12.49028234200656
+         79.6232585491842
+        3.484731698258543
+        5.642355936390698
+         8.71909310716887
+        76.14769015508216
+ 9e+09       
+        79.51963211802493
+        8.970068648952594
+        80.29822394031369
+         5.70328871675104
+         12.6687778573511
+        80.18471536157229
+        3.573899936510043
+        5.764751489910124
+        8.855334280314425
+        76.68331244106648
+ 9.1e+09     
+        80.07130735399349
+        9.112795519937297
+        80.85626354381731
+        5.828662222961936
+        12.85280018324654
+        80.74293197094229
+        3.670412739760577
+        5.889784386410284
+        8.995281586668618
+        77.21531277410226
+ 9.2e+09     
+        80.61854477681395
+        9.258852145735844
+        81.41056945710616
+        5.956115803811822
+        13.04188643972212
+         81.2977021135989
+        3.775244105938817
+        6.017441552607247
+        9.139514842542338
+            77.7435643707
+ 9.3e+09     
+        81.16115227246335
+        9.408683894616557
+        81.96088865211748
+        6.085520963561841
+        13.23553091742649
+         81.8488276150149
+        3.889436047326214
+        6.147699241937942
+        9.288674473379224
+        78.26795609605456
+ 9.4e+09     
+        81.69894845492976
+          9.5627807019412
+        82.50697309759342
+        6.216728231757042
+        13.43319224198906
+        82.39612049665037
+        4.014101692818786
+        6.280522431233059
+        9.443464364682583
+        78.78839346552945
+ 9.5e+09     
+        82.23176333396947
+        9.721678878149929
+         83.0485814109625
+        6.349565680407906
+        13.63429959373998
+        82.93940490992789
+        4.150428448860445
+        6.415863808631421
+         9.60465466091912
+        79.30479962161841
+ 9.6e+09     
+        82.75943895564417
+        9.885962857886437
+        83.58548034232514
+        6.483837032783928
+        13.83825803182647
+        83.47851890464676
+        4.299681219312694
+         6.55366233695756
+        9.773084507089877
+        79.81711628484612
+ 9.7e+09     
+        83.28183001570417
+        10.05626688967877
+         84.1174461009429
+        6.619319355803212
+        14.04445298519778
+        84.01331604120432
+         4.46320568459376
+        6.693841378087971
+         9.94966472763091
+        80.32530467694322
+ 9.8e+09     
+        83.79880444585595
+        10.23327666567078
+         84.6442655356111
+         6.75576032912666
+        14.25225397946364
+        84.54366685691669
+        4.642431640320248
+        6.836306364228728
+        10.13538043698965
+        80.82934641443174
+ 9.9e+09     
+        84.31024397287686
+        10.41773089078248
+        85.16573718044023
+        6.892875084660892
+        14.46101767016425
+        85.06946019678479
+        4.838876395473904
+        6.980942001878422
+         10.3312935757031
+        81.32924437054413
+ 1e+10       
+        84.81604465047202
+        10.61042279043266
+        85.68167217712174
+        7.030342610544302
+        14.67009025108539
+        85.59060441854601
+        5.054148229843528
+        7.127608993862992
+        10.53854536516506
+         81.8250235031658
+ 1.01e+10    
+        84.89643805549137
+        10.48982771951026
+        85.71505501472609
+        6.969545134059105
+        14.50999242878632
+        85.66376329093481
+        5.038011685041097
+        7.066566183012172
+        10.42155914832356
+        81.88322467214805
+ 1.02e+10    
+        84.98949755872313
+        10.37798332289066
+        85.76859018295582
+        6.913419625089061
+        14.36322046457863
+        85.75386228854681
+        5.024131733676015
+        7.010295406597599
+        10.31296951625201
+        81.95431485581983
+ 1.03e+10    
+        85.09506749615508
+        10.27475656076539
+        85.84166262924856
+        6.861910938943441
+        14.22939955524285
+        85.86047190813954
+         5.01249058957216
+        6.958735555742377
+        10.21266395523455
+        82.03813709546317
+ 1.04e+10    
+         85.2129885942288
+        10.18001408873451
+        85.93367116237543
+        6.814963517971915
+        14.10816321314352
+        85.98316736558466
+        5.003069557182215
+        6.911825386174337
+        10.12052864000737
+        82.13453066766667
+ 1.05e+10    
+        85.34309828090429
+        10.09362240217427
+        86.04402841059525
+        6.772521429268772
+        13.99915321612747
+        86.12152895154441
+        4.995849067908524
+          6.8695035446835
+        10.03644862146388
+        82.24333140410499
+ 1.06e+10    
+        85.48523098595176
+         10.0154479720677
+        86.17216075388252
+        6.734528400402042
+        13.90201954444442
+        86.27514234787898
+        4.990808715669071
+        6.831708593958757
+        9.960308004392829
+        82.36437200035182
+ 1.07e+10    
+        85.63921843053666
+        9.945357372705812
+        86.31750823304952
+        6.700927853350858
+        13.81642030623202
+        86.44359890759823
+        4.987927291704778
+        6.798379035980908
+        9.891990115655355
+         82.4974823137791
+ 1.08e+10    
+         85.8048899062039
+        9.883217401650857
+         86.4795244383392
+        6.671662936789882
+        13.74202165296579
+         86.6264959010046
+        4.987182818618761
+        6.769453334117015
+        9.831377663199419
+        82.64248965064495
+ 1.09e+10    
+        85.98207254336289
+        9.828895192331274
+          86.657676379851
+        6.646676556869533
+        13.67849768614762
+        86.82343673049563
+        4.988552583646748
+        6.744869934057661
+        9.778352886289902
+         82.7992190424727
+ 1.1e+10     
+        86.17059156942013
+        9.782258319622754
+        86.85144434195894
+         6.62591140660398
+        13.62553035639061
+        87.03403111637378
+        4.992013171156359
+        6.724567283719677
+         9.73279769733125
+        82.96749351185765
+ 1.11e+10    
+        86.37027055669375
+        9.743174898750413
+        87.06032172368637
+        6.609309993993641
+        13.58280935594708
+        87.25789525582826
+        4.997540494374228
+        6.708483852218041
+        9.694593815634537
+        83.14713432783969
+ 1.12e+10    
+        86.58093166028701
+        9.711513677836097
+         87.2838148668431
+        6.596814668973089
+        13.55003200563364
+        87.49465195714828
+         5.00510982634462
+        6.696558148006126
+         9.66362289348123
+        83.33796125100973
+ 1.13e+10    
+        86.80239584608834
+        9.687144124394004
+        87.52144287355883
+        6.588367649277287
+        13.52690313701128
+        87.74393075107572
+        5.014695830121109
+        6.688728736268455
+         9.63976663481496
+        83.53979276852402
+ 1.14e+10    
+        87.03448310908314
+        9.669936506067245
+        87.77273741470904
+         6.58391104531109
+        13.51313497060107
+         88.0053679810925
+        5.026272588196187
+        6.684934255638638
+        9.622906906885543
+        83.75244631920704
+ 1.15e+10    
+         87.2770126821849
+        9.659761965886485
+        88.03724253059607
+        6.583386884096012
+        13.50844699083776
+        88.27860687431546
+        5.039813631175639
+          6.6851134343129
+        9.612925845157255
+        83.97573850894607
+ 1.16e+10    
+        87.52980323577611
+         9.65649259231315
+        88.31451442511657
+        6.586737132352068
+        13.51256581839604
+        88.56329759457121
+        5.055291965702565
+        6.689205105611332
+        9.609705951782418
+        84.20948531658046
+ 1.17e+10    
+         87.7926730681864
+         9.66000148432528
+        88.60412125454566
+        6.593903718786303
+        13.52522508046086
+        88.85909727910553
+        5.072680101641353
+        6.697148223041051
+        9.613130187929226
+        84.45350229049875
+ 1.18e+10    
+         88.0654402873121
+        9.670162811784881
+        88.90564291195004
+        6.604828555630326
+        13.54616527945657
+        89.16567006029777
+        5.091950078529013
+         6.70888187490587
+        9.623082060243361
+         84.7076047361605
+ 1.19e+10    
+        88.34792298360915
+        9.686851871321704
+        89.21867080815963
+        6.619453559480053
+        13.57513366069556
+        89.48268707365206
+        5.113073491303832
+        6.724345298496829
+        9.639445701712365
+        84.97160789477311
+ 1.2e+10     
+         88.6399393946818
+        9.709945137953683
+        89.54280765012841
+         6.63772067147551
+        13.61188407936118
+        89.80982645325199
+        5.136021515321763
+        6.743477893898316
+        9.662105947191753
+        85.24532711334558
+ 1.21e+10    
+        88.94130806169912
+        9.739320312655757
+        89.87766721744354
+        6.659571876860355
+         13.6561768671955
+        90.14677331578422
+        5.160764930672434
+        6.766219237441803
+         9.69094840384134
+          85.528578006358
+ 1.22e+10    
+        89.25184797786542
+        9.774856366079518
+        90.22287413766149
+        6.684949223959473
+        13.70777869922169
+        90.49321973415798
+        5.187274145806097
+        6.792509094824295
+        9.725859516708951
+        85.82117660927048
+ 1.23e+10    
+        89.57137872918449
+         9.81643357861706
+        90.57806366108311
+        6.713794842587451
+        13.76646246079598
+        90.84886470168532
+        5.215519220481761
+        6.822287433914296
+        9.766726629696713
+        86.12293952412077
+ 1.24e+10    
+        89.89972062774247
+        9.863933576994317
+        90.94288143552387
+        6.746050961939638
+        13.83200711525126
+        91.21341408769943
+        5.245469888053448
+        6.855494437267456
+         9.81343804212365
+        86.43368405743315
+ 1.25e+10    
+        90.23669483774641
+        9.917239367568195
+        91.31698328156405
+        6.781659927960547
+        13.90419757236351
+        91.58658058545699
+          5.2770955771027
+        6.892070514359654
+        9.865883061103487
+        86.75322835068312
+ 1.26e+10    
+        90.58212349455015
+        9.976235366500321
+        91.70003496873105
+        6.820564220238172
+        13.98282455784493
+         91.9680836530694
+        5.310365432434232
+        6.931956313550094
+         9.92395204993524
+        87.08139150354924
+ 1.27e+10    
+        90.93582981689291
+        10.04080742696342
+        92.09171199299787
+        6.862706468414648
+        14.06768448404463
+        92.35764944819819
+        5.345248335445661
+        6.975092733788681
+        9.987536472706138
+        87.41799369018639
+ 1.28e+10    
+        91.29763821258577
+        10.11084286353939
+        92.49169935595393
+        6.908029468152487
+        14.15857932201261
+        92.75501075715808
+        5.381712923886758
+        7.021420936069077
+        10.05652893529119
+        87.76285626875489
+ 1.29e+10    
+        91.66737437786392
+        10.18623047395311
+        92.89969134595808
+        6.956476196656863
+        14.25531647506637
+        93.15990691905289
+        5.419727611020367
+        7.070882354634385
+        10.13082322293122
+        88.11580188443119
+ 1.3e+10     
+        92.04486539063163
+        10.26686055828176
+        93.31539132154107
+        7.007989827766587
+        14.35770865397438
+        93.57208374550007
+        5.459260604199964
+        7.123418707945548
+        10.21031433455837
+        88.47665456612964
+ 1.31e+10    
+        92.42993979782162
+        10.35262493577884
+        93.73851149730663
+          7.0625137466355
+        14.46557375386319
+        93.99129343647679
+        5.500279922877343
+        7.178972009407993
+        10.29489851403714
+        88.84523981716089
+ 1.32e+10    
+        92.82242769707631
+        10.44341695943504
+        94.16877273253371
+        7.119991563997626
+        14.57873473293041
+        94.41729449276845
+        5.542753416053413
+        7.237484577861556
+        10.38447327847603
+        89.22138470004307
+ 1.33e+10    
+        93.22216081297533
+        10.53913152840229
+         94.6059043226644
+        7.180367130037038
+        14.69701949303918
+        94.84985162546712
+        5.586648779186829
+        7.298899047838038
+        10.47893744376182
+        89.60491791568511
+ 1.34e+10    
+        93.62897256800434
+        10.63966509839686
+        95.04964379383377
+         7.24358454786516
+        14.82026076225274
+        95.28873566293559
+        5.631933570573475
+        7.363158379576831
+        10.57819114746142
+        89.99566987715775
+ 1.35e+10    
+         94.0426981484828
+        10.74491569019329
+        95.49973670057527
+        7.309588186612061
+        14.94829597936066
+        95.73372345561387
+        5.678575227211016
+        7.430205868813253
+        10.68213586922864
+        90.39347277825394
+ 1.36e+10    
+        94.46317456563534
+        10.85478289631479
+        95.95593642681463
+        7.378322694133028
+        15.08096718043369
+        96.18459777902299
+        5.726541080159944
+        7.499985156323119
+        10.79067444884765
+        90.79816065704912
+ 1.37e+10    
+        94.89024071201558
+        10.96916788602322
+        96.41800399024285
+        7.449733009347566
+        15.21812088743938
+        96.64114723528498
+        5.775798369417434
+        7.572440237235506
+        10.90371110204117
+        91.20956945465804
+ 1.38e+10    
+        95.32373741346247
+        11.08797340870448
+        96.88570785015075
+        7.523764374201225
+         15.3596079989404
+        97.10316615345918
+        5.826314258313716
+        7.647515470100139
+        11.02115143416305
+        91.62753706938474
+ 1.39e+10    
+        95.76350747678262
+        11.21110379574245
+        97.35882371877733
+        7.600362345262552
+        15.50528368288966
+        97.57045448896206
+        5.878055847445964
+        7.725155585721378
+         11.1429024518888
+        92.05190340645305
+ 1.4e+10     
+         96.2093957333323
+        11.33846496096917
+        97.83713437622534
+        7.679472804958314
+         15.6550072715324
+        98.04281772232585
+        5.930990188161509
+        7.805305695742705
+        11.26887257301915
+        92.48251042350834
+ 1.41e+10    
+        96.66124907867912
+        11.46996439977602
+        98.32042948897454
+        7.761041972446296
+        15.80864215841599
+        98.52006675751979
+        5.985084295602039
+        7.887911300989376
+          11.398971634495
+        92.91920217206174
+ 1.42e+10    
+        97.11891650851257
+        11.60551118696505
+        98.80850543201622
+        7.845016414132463
+        15.96605569750687
+        99.00201782004083
+         6.04030516132191
+        7.972918299564816
+         11.5331108987305
+        93.36182483506528
+ 1.43e+10    
+        97.58224915097331
+        11.74501597341871
+         99.3011651146155
+          7.9313430538363
+        16.12711910440644
+         99.4884923549733
+        6.096619765492029
+        8.060272994696252
+        11.67120305835651
+         93.8102267607742
+ 1.44e+10    
+        98.05110029555468
+        11.88839098165826
+         99.7982178097146
+         8.01996918260104
+        16.29170735965529
+         99.9793169251782
+        6.153995088700261
+         8.14992210233298
+        11.81316223946512
+        94.26425849307404
+ 1.45e+10    
+        98.52532541873875
+         12.0355500003626
+        100.2994789869591
+        8.110842468159166
+        16.45969911411096
+        100.4743231097789
+        6.212398123360179
+        8.241812758488972
+        11.95890400344632
+        94.72377279842425
+ 1.46e+10    
+        99.00478220651642
+        12.18640837791141
+        100.8047701493395
+        8.203910964050138
+        16.63097659638101
+        100.9733474030828
+        6.271795884738901
+        8.335892526331044
+        12.10834534749502
+        95.18862468958093
+ 1.47e+10    
+        99.48933057393789
+        12.34088301501751
+        101.3139186734309
+         8.29912311839443
+        16.80542552229247
+        101.4762311140692
+        6.332155421614915
+         8.43210940301827
+        12.26140470387105
+        95.65867144624016
+ 1.48e+10    
+        99.97883268183229
+         12.4988923565069
+        101.8267576531962
+        8.396427782333133
+        16.98293500637219
+        101.9828202665579
+        6.393443826576178
+        8.530411826273347
+        12.41800193798583
+        96.13377263276018
+ 1.49e+10    
+        100.4731529508403
+        12.66035638230337
+        102.3431257473295
+        8.495774218115724
+        17.16339747531426
+        102.4929655001672
+        6.455628245967597
+        8.630748680706299
+        12.57805834538863
+        96.61379011309083
+ 1.5e+10     
+        100.9721580728817
+        12.82519659767289
+         102.862867030099
+        8.597112106870947
+        17.34670858340866
+         103.006521972148
+        6.518675889500443
+        8.733069303873693
+        12.74149664771891
+         97.0985880630531
+ 1.51e+10    
+        101.4757170201965
+        12.99333602277847
+        103.3858308456514
+        8.700391556030828
+        17.53276712990101
+        103.5233492601941
+        6.582554039529814
+        8.837323492080131
+        12.90824098769313
+        97.58803298010083
+ 1.52e+10    
+        101.9837010520733
+        13.16469918159376
+        103.9118716657311
+        8.805563106429409
+        17.72147497825385
+        104.0433112662809
+        6.647230060011745
+        8.943461505919936
+        13.07821692318412
+        98.08199369068841
+ 1.53e+10    
+         102.495983719388
+        13.33921209022464
+        104.4408489507742
+        8.912577739080238
+        17.91273697728076
+        104.5662761216205
+        6.712671405148971
+        9.051434075559971
+        13.25135142045492
+        98.58034135536455
+ 1.54e+10    
+        103.0124408670677
+        13.51680224467889
+        104.9726270143169
+        9.021386881620074
+        18.10646088411784
+        105.0921160927771
+        6.778845627731471
+        9.161192405757191
+        13.42757284660148
+        99.08294947171896
+ 1.55e+10    
+         103.532950634586
+        13.69739860812968
+        105.5070748906766
+         9.13194241444187
+        18.30255728900492
+        105.6207074890036
+        6.845720387184604
+        9.272688180625511
+        13.60681096125913
+        99.58969387528634
+ 1.56e+10    
+        104.0573934546001
+         13.8809315977107
+        106.0440662058498
+        9.244196676502371
+        18.50093954183887
+        106.1519305708324
+        6.913263457328464
+        9.385873568136303
+        13.78899690762082
+        100.1004527385181
+ 1.57e+10    
+        104.5856520498259
+         14.0673330708819
+        106.5834790515673
+        9.358102470824534
+        18.70152368046947
+        106.6856694599754
+        6.981442733859884
+        9.500701224361364
+        13.97406320281866
+        100.6151065679336
+ 1.58e+10    
+        105.1176114282572
+         14.2565363113999
+        107.1251958624513
+        9.473613069680328
+        18.90422836070152
+        107.2218120505479
+        7.050226241562903
+        9.617124297465114
+         14.1619437277118
+        101.1335381995439
+ 1.59e+10    
+        105.6531588768104
+        14.44847601492995
+        107.6691032962235
+        9.590682219473727
+        19.10897478797088
+        107.7602499216585
+        7.119582141255229
+        9.735096431432089
+        14.35257371612586
+        101.6556327926501
+ 1.6e+10     
+        106.1921839534985
+        14.64308827432919
+        108.2150921168967
+        9.709264145319539
+        19.31568665066063
+        108.3008782513755
+        7.189478736479376
+        9.854571769547421
+         14.5458897435832
+        102.1812778221057
+ 1.61e+10    
+        106.7345784782118
+        14.84031056463257
+        108.7630570808951
+        9.829313555319839
+        19.52429005502167
+        108.8435957320989
+        7.259884479943096
+         9.97550495762037
+        14.74182971556634
+        102.7103630691362
+ 1.62e+10    
+        107.2802365221901
+        15.04008172777248
+         109.312896826048
+        9.950785644549772
+        19.73471346166695
+         109.388304487343
+        7.330767979717862
+        10.09785114695927
+        14.94033285534709
+        103.2427806108014
+ 1.63e+10    
+        107.8290543962691
+        15.24234195705551
+        109.8645137633872
+        10.07363609874901
+        19.94688762360267
+         109.934909989948
+        7.402098005201326
+        10.22156599709947
+        15.14133969142261
+        103.7784248081764
+ 1.64e+10    
+         108.380930637973
+        15.44703278142599
+        110.4178139716979
+          10.197821097732
+        20.16074552576563
+        110.4833209817184
+        7.473843492849161
+        10.34660567828121
+        15.34479204458562
+        104.3171922933414
+ 1.65e+10    
+        108.9357659975278
+        15.65409704953947
+        110.9727070947611
+        10.32329731850794
+        20.37622232603175
+        111.0334493945035
+        7.545973551683881
+        10.47292687368905
+        15.55063301466467
+        104.8589819552455
+ 1.66e+10    
+        109.4934634228695
+        15.86347891366944
+        111.5291062412264
+        10.45002193813027
+        20.59325529766413
+        111.5852102727099
+        7.618457468585204
+        10.60048678144786
+        15.75880696696319
+        105.4036949245207
+ 1.67e+10    
+        110.0539280437019
+         16.0751238134687
+        112.0869278870548
+        10.57795263627003
+        20.81178377316801
+        112.1385216972521
+        7.691264713368831
+        10.72924311638332
+        15.96925951842484
+        105.9512345573174
+ 1.68e+10    
+        110.6170671546852
+        16.28897845960822
+        112.6460917804807
+        10.70704759752078
+        21.03174908952031
+        112.6933047109352
+        7.764364943658244
+        10.85915411154582
+        16.18193752355469
+        106.5015064182269
+ 1.69e+10    
+        111.1827901978004
+        16.50499081731081
+        113.2065208494249
+        10.83726551344062
+         21.2530945347429
+        113.2494832452643
+        7.837728009555033
+        10.99017851950591
+        16.39678906011736
+        107.0544182623483
+ 1.7e+10     
+        111.7510087439585
+        16.72311008979952
+        113.7681411113107
+        10.96856558433287
+        21.47576529578741
+        113.8069840486699
+        7.911323958113853
+        11.12227561341996
+        16.61376341464147
+        107.6098800165694
+ 1.71e+10    
+         112.321636473903
+        16.94328670167762
+        114.3308815852182
+         11.1009075207777
+        21.69970840770257
+        114.3657366161458
+        7.985123037625307
+        11.25540518787362
+        16.83281106774865
+         108.167803760113
+ 1.72e+10    
+        112.8945891584653
+        17.16547228225764
+        114.8946742063276
+        11.23425154491174
+        21.92487270405273
+        114.9256731202817
+        8.059095701713918
+        11.38952755950482
+        17.05388367933141
+        108.7281037044064
+ 1.73e+10    
+        113.4697846382199
+        17.38961964885372
+        115.4594537425944
+        11.36855839146035
+        22.15120876855881
+        115.4867283436865
+        8.133212613253081
+        11.52460356740977
+         17.2769340735997
+        109.2906961723251
+ 1.74e+10    
+        114.0471428025858
+        17.61568279005254
+        116.0251577135973
+        11.50378930854003
+        22.37866888793148
+        116.0488396127773
+        8.207444648104238
+        11.66059457333661
+        17.50191622401395
+        109.8554995768632
+ 1.75e+10    
+        114.6265855684266
+        17.84361684897744
+        116.5917263115136
+        11.63990605821966
+        22.60720700587023
+        116.6119467329313
+        8.281762898683237
+        11.79746246167175
+        17.72878523812481
+        110.4224343992753
+ 1.76e+10    
+        115.2080368581873
+        18.07337810655681
+        117.1591023241637
+        11.77687091685402
+        22.83677867819819
+         117.175991924978
+        8.356138677357876
+          11.935169639222
+        17.95749734233559
+        110.9914231667389
+ 1.77e+10    
+        115.7914225776112
+        18.30492396481138
+        117.7272310600758
+        11.91464667520048
+          23.067341029107
+         117.740919763017
+        8.430543519682288
+        12.07367903479498
+        18.18800986660386
+        111.5623904295768
+ 1.78e+10    
+        116.3766705930797
+        18.53821293016892
+        118.2960602755186
+        12.05319663830814
+        23.29885270848357
+        118.3066771135444
+        8.504949187470425
+         12.2129540985865
+        18.42028122909666
+         112.135262738086
+ 1.79e+10    
+        116.9637107086072
+        18.77320459682023
+        118.8655401034535
+        12.19248462520445
+        23.53127385029416
+        118.8732130758681
+        8.579327671714363
+         12.3529588013756
+        18.65427092081507
+        112.7099686190048
+ 1.8e+10     
+         117.552474642533
+        19.00985963012402
+        119.4356229843579
+        12.33247496836536
+         23.7645660319981
+        119.4404789237991
+        8.653651195349152
+          12.493657633533
+        18.88993949020087
+        113.2864385516666
+ 1.81e+10    
+         118.142896003939
+        19.24813975007159
+        120.0062635988702
+        12.47313251299203
+        23.99869223496817
+        120.0084280485931
+        8.727892215870169
+        12.63501560384714
+        19.12724852773669
+        113.8646049438605
+ 1.82e+10    
+        118.7349102688315
+        19.48800771481925
+        120.5774188022126
+        12.61442261608341
+        24.23361680589138
+        120.5770159031259
+        8.802023427804578
+         12.7769982381726
+        19.36616065055532
+        114.4444021074509
+ 1.83e+10    
+        119.3284547561098
+        19.72942730429735
+        121.1490475603418
+        12.75631114532338
+        24.46930541912681
+        121.1461999472888
+        8.876017765041901
+        12.91957157790647
+        19.60663948706505
+        115.0257662337716
+ 1.84e+10    
+        119.9234686033619
+        19.97236330390315
+        121.7211108877889
+        12.89876447777732
+        24.70572503999733
+        121.7159395945694
+        8.949848403026083
+        13.06270217829455
+        19.84864966160305
+        115.6086353688334
+ 1.85e+10    
+        120.5198927425022
+        20.21678148828559
+        122.2935717871398
+        13.04174949841319
+        24.94284388899246
+         122.286196159818
+        9.023488760813354
+        13.20635710657682
+        20.09215677912963
+        116.1929493883745
+ 1.86e+10    
+        121.1176698752904
+        20.46264860522685
+        122.8663951901157
+        13.18523359844413
+        25.18063140685853
+        122.8569328081601
+        9.096912502997666
+        13.35050393996801
+        20.33712740996724
+        116.7786499727752
+ 1.87e+10    
+        121.7167444487434
+        20.70993235962907
+        123.4395479002096
+        13.32918467349857
+        25.41905822055574
+        123.4281145050501
+        9.170093541508292
+         13.4951107634898
+        20.58352907459744
+        117.3656805818703
+ 1.88e+10    
+        122.3170626304762
+        20.95860139760996
+        124.0129985368444
+        13.47357112163071
+        25.65809611006093
+        123.9997079674342
+        9.243006037282202
+           13.64014616765
+        20.83133022852163
+        117.9539864296767
+ 1.89e+10    
+        122.9185722839862
+        21.20862529071595
+        124.5867174810054
+        13.61836184117053
+        25.89771797599466
+        124.5716816160115
+        9.315624401814144
+        13.78557924597746
+        21.08050024719363
+        118.5435144590621
+ 1.9e+10     
+        123.5212229439014
+        21.45997452025142
+        125.1606768223109
+        13.76352622841491
+        26.13789780805071
+         125.144005528566
+        9.387923298586493
+        13.93137959241423
+        21.33100941103106
+        119.1342133163797
+ 1.91e+10    
+         124.124965791218
+        21.71262046173724
+        125.7348503074882
+        13.90903417517606
+        26.37861065421256
+         125.716651394355
+        9.459877644383871
+         14.0775172985748
+         21.5828288905127
+        119.7260333260854
+ 1.92e+10    
+         124.729753628543
+        21.96653536949524
+        126.3092132902092
+         14.0548560661804
+        26.61983259073229
+        126.2895924695283
+        9.531462610493168
+        14.22396295087331
+        21.83593073136696
+        120.3189264653568
+ 1.93e+10    
+        125.3355408553575
+         22.2216923613662
+        126.8837426822568
+         14.2009627763323
+        26.86154069285704
+        126.8628035335647
+        9.602653623792774
+        14.37068762752164
+        22.09028783985754
+        120.9128463387353
+ 1.94e+10    
+        125.9422834433199
+        22.47806540356502
+        127.4584169059855
+        14.34732566784087
+        27.10371300628242
+        127.4362608466995
+        9.673426367733443
+        14.51766289540718
+        22.34587396817243
+        121.5077481528098
+ 1.95e+10    
+        126.5499389116257
+        22.73562929567413
+        128.0332158480388
+        14.49391658721928
+        27.34632851931576
+        128.0099421083285
+        9.743756783213591
+        14.66486080685313
+        22.60266369991901
+        122.1035886909488
+ 1.96e+10    
+        127.1584663024337
+         22.9943596557801
+        128.6081208142932
+        14.64070786216122
+        27.58936713573176
+        128.5838264163638
+        9.813621069351571
+        14.81225389626436
+        22.86063243573233
+        122.7003262881113
+ 1.97e+10    
+        127.7678261563799
+        23.25423290575533
+        129.1831144859987
+        14.78767229829469
+        27.83280964830375
+         129.157894227531
+        9.882995684157027
+        14.95981517666577
+        23.11975637899881
+        123.2979208057373
+ 1.98e+10    
+        128.3779804881844
+        23.51522625668778
+        129.7581808770781
+        14.93478317582266
+        28.07663771299215
+        129.7321273185784
+          9.9518573451038
+        15.10751813613322
+        23.38001252169959
+        123.8963336067399
+ 1.99e+10    
+        128.9888927623679
+        23.77731769445806
+        130.3333052925577
+         15.0820142460578
+        28.32083382377681
+        130.3065087483832
+        10.02018302960838
+        15.25533673412883
+        23.64137863037789
+        124.4955275306051
+ 2e+10       
+         129.600527869089
+        24.04048596547143
+        130.9084742881032
+        15.22933972784361
+        28.56538128811538
+        130.8810228209441
+        10.08794997541314
+        15.40324539773656
+        23.90383323223244
+        125.0954668686187
+ 2.01e+10    
+          130.21285210011
+        24.30471056253959
+        131.4836756306219
+        15.37673430388412
+        28.81026420301236
+        131.4556550492253
+           10.15513568088
+        15.55121901780824
+        24.16735560134019
+        125.6961173392255
+ 2.02e+10    
+        130.8258331249089
+        24.56997171092051
+        132.0588982599167
+         15.5241731169712
+        29.05546743168542
+        132.0303921198534
+        10.22171790519463
+        15.69923294502022
+         24.4319257450124
+        126.2974460635335
+ 2.03e+10    
+        131.4394399669329
+        24.83625035451092
+        132.6341322513494
+        15.67163176612272
+        29.30097658081233
+        132.6052218586323
+        10.28767466848413
+        15.84726298584941
+        24.69752439028345
+        126.8994215409714
+ 2.04e+10    
+         132.053642980017
+        25.10352814219801
+        133.2093687794981
+        15.81908630263261
+         29.5467779783459
+        133.1801331968698
+        10.35298425185052
+        15.99528539846873
+        24.96413297053729
+        127.5020136251096
+ 2.05e+10    
+        132.6684138249669
+         25.3717874143682
+        133.7846000827761
+        15.96651322603983
+        29.79285865188156
+        133.7551161384946
+        10.41762519732193
+        16.14327688856422
+        25.23173361227321
+        128.1051934996545
+ 2.06e+10    
+        133.2837254463151
+        25.64101118957435
+        134.3598194289904
+         16.1138894800144
+        30.03920630756585
+        134.3301617279454
+        10.48157630772371
+        16.29121460508674
+        25.50030912200989
+        128.7089336546206
+ 2.07e+10    
+        133.8995520492608
+        25.91118315136377
+        134.9350210818131
+        16.26119244817255
+         30.2858093095309
+        134.9052620188189
+         10.5448166464717
+        16.43907613593115
+        25.76984297333333
+        129.3132078626883
+ 2.08e+10    
+        134.5158690767918
+        26.18228763526253
+        135.5102002681414
+        16.40839994982188
+        30.53265665984333
+        135.4804100432606
+        10.60732553728922
+        16.58683950355332
+        26.04031929408652
+        129.9179911557568
+ 2.09e+10    
+        135.1326531870067
+        26.45430961592351
+        136.0853531463253
+        16.55549023563323
+        30.77973797895347
+        136.0555997820741
+        10.66908256385054
+        16.73448316052785
+        26.31172285370401
+         130.523259801696
+ 2.1e+10     
+        135.7498822306282
+        26.72723469443171
+        136.6604767752356
+         16.7024419832594
+        31.02704348663518
+        136.6308261355473
+        10.73006756935234
+        16.88198598504835
+         26.5840390506911
+        131.1289912813004
+ 2.11e+10    
+        136.3675352287251
+        27.00104908577135
+        137.2355690841599
+        16.84923429288602
+        31.27456398340175
+        137.2060848949678
+        10.79026065601445
+        17.02932727637397
+        26.85725390024998
+        131.7351642654576
+ 2.12e+10    
+        136.9855923506408
+        27.27573960645131
+         137.810628843487
+        16.99584668273296
+        31.52229083238754
+        137.7813727148167
+        10.84964218451378
+        17.17648675022978
+        27.13135402205058
+        132.3417585925279
+ 2.13e+10    
+        137.6040348921315
+        27.55129366229255
+        138.3856556361821
+        17.14225908450249
+        31.77021594168532
+        138.3566870856311
+        10.90819277335111
+        17.32344453415715
+        27.40632662815173
+        132.9487552459452
+ 2.14e+10    
+        138.2228452537266
+        27.82769923637244
+         138.960649830012
+        17.28845183877615
+         32.0183317471244
+        138.9320263075058
+        10.96589329815368
+        17.47018116282495
+        27.68215951106528
+        133.5561363320381
+ 2.15e+10    
+        138.8420069192987
+        28.10494487713085
+        139.5356125505122
+        17.43440569037221
+        32.26663119548351
+        139.5073894642423
+         11.0227248909154
+        17.61667757329759
+        27.95884103197298
+        134.1638850580817
+ 2.16e+10    
+        139.4615044348638
+        28.38301968663177
+        140.1105456546724
+        17.58010178365978
+        32.51510772812554
+        140.0827763981094
+        11.07866893917665
+        17.76291510027178
+        28.23636010908622
+        134.7719857105731
+ 2.17e+10    
+        140.0813233876046
+          28.661913308986
+        140.6854517053238
+        17.72552165783202
+        32.76375526504269
+        140.6581876852145
+        11.13370708514432
+        17.90887547127527
+        28.51470620615736
+        135.3804236337442
+ 2.18e+10    
+        140.7014503851178
+        28.94161591892951
+        141.2603339462081
+         17.8706472421494
+        33.01256818930569
+        141.2336246114695
+        11.18782122475552
+        18.05454080183982
+        28.79386932113676
+        135.9891852083069
+ 2.19e+10    
+        141.3218730348931
+        29.22211821055744
+        141.8351962777088
+        18.01546085114802
+        33.26154133190337
+        141.8090891491327
+        11.24099350668513
+        18.19989359064343
+        29.07383997497756
+        136.5982578304354
+ 2.2e+10     
+         141.942579924024
+        29.50341138621649
+        142.4100432332336
+        18.15994517982236
+         33.5106699569669
+         142.384583933927
+        11.29320633130013
+        18.34491671463119
+        29.35460920058787
+        137.2076298909876
+ 2.21e+10    
+        142.5635605991499
+        29.78548714554984
+        142.9848799562272
+        18.30408329877807
+        33.75994974736589
+        142.9601122427031
+        11.34444234956115
+        18.48959342411351
+        29.63616853192924
+        137.8172907549661
+ 2.22e+10    
+        143.1848055466305
+        30.06833767469734
+        143.5597121777928
+        18.44785864936636
+        34.00937679067053
+        143.5356779716534
+         11.3946844618738
+         18.6339073378452
+        29.91850999326195
+        138.4272307412218
+ 2.23e+10    
+        143.8063061729588
+        30.35195563564801
+        144.1345461949215
+        18.59125503879732
+        34.25894756546919
+        144.1112856150508
+        11.44391581689158
+        18.77784243809116
+        30.20162608853543
+        139.0374411023989
+ 2.24e+10    
+        144.4280547854073
+        30.63633415574485
+        144.7093888492958
+        18.73425663523481
+        34.50865892803284
+         144.686940244513
+        11.49211981027043
+        18.92138306567477
+        30.48550979092411
+        139.6479140051252
+ 2.25e+10    
+        145.0500445729092
+        30.92146681734014
+        145.2842475066675
+        18.87684796287755
+        34.75850809931939
+        145.2626474887649
+         11.5392800833783
+        19.06451391501842
+        30.77015453250683
+        140.2586425104445
+ 2.26e+10    
+        145.6722695871793
+        31.20734764760063
+        145.8591300367839
+         19.0190138970314
+        35.00849265230868
+        145.8384135139063
+        11.58538052196048
+        19.20722002917578
+         31.0555541940912
+        140.8696205544949
+ 2.27e+10    
+        146.2947247240705
+        31.49397110846144
+        146.4340447938586
+        19.16073965916505
+        35.25861049966007
+         146.414245004159
+        11.63040525476148
+         19.3494867948559
+         31.3417030951793
+        141.4808429294316
+ 2.28e+10    
+        146.9174057051666
+        31.78133208672687
+         147.009000597563
+        19.30201081196859
+        35.50885988168598
+        146.9901491430873
+        11.67433865210672
+        19.49129993744412
+        31.62859598407526
+        142.0923052645931
+ 2.29e+10    
+        147.5403090596108
+        32.06942588431696
+        147.5840067145349
+        19.44281325439689
+        35.75923935463259
+        147.5661335952868
+        11.71716532444347
+        19.63264551602498
+        31.91622802813575
+        142.7040040079146
+ 2.3e+10     
+        148.1634321061741
+         32.3582482086599
+        148.1590728403782
+        19.58313321672203
+        36.00974777926191
+        148.1422064885205
+        11.75887012084416
+        19.77350991839949
+        32.20459480415725
+        143.3159364075837
+ 2.31e+10    
+        148.7867729355575
+        32.64779516322675
+        148.7342090821591
+         19.7229572555738
+        36.26038430972625
+        148.7183763963033
+        11.79943812747212
+        19.91387985611135
+        32.49369228890517
+        143.9281004939403
+ 2.32e+10    
+        149.4103303929268
+          32.938063238208
+        149.3094259413668
+        19.86227224899237
+        36.51114838272895
+        149.2946523209138
+        11.83885466601224
+        20.05374235947298
+         32.7835168497783
+        144.5404950616197
+ 2.33e+10    
+        150.0341040606889
+        33.22904930133296
+        149.8847342973428
+        20.00106539147924
+         36.7620397069661
+        149.8710436768352
+        11.87710529206744
+        20.19308477260279
+        33.07406523561247
+        145.1531196519384
+ 2.34e+10    
+        150.6580942414958
+        33.52075058882551
+         150.460145391155
+        20.13932418905543
+        37.01305825283875
+        150.4475602746043
+        11.91417579352191
+        20.33189474846694
+        33.36533456761717
+        145.7659745355223
+ 2.35e+10    
+        151.2823019414817
+        33.81316469649914
+        151.0356708099153
+        20.27703645433031
+        37.26420424243441
+        151.0242123050708
+        11.95005218887313
+        20.47016024393518
+        33.65732233044901
+        146.3790606951721
+ 2.36e+10    
+        151.9067288537395
+         34.1062895709902
+        151.6113224715218
+        20.41419030157569
+        37.51547813976522
+        151.6010103240464
+         11.9847207255335
+        20.60786951484477
+        33.95002636341637
+        146.9923798089722
+ 2.37e+10    
+        152.5313773420172
+        34.40012350112222
+        152.1871126098178
+        20.55077414181598
+        37.76688064126351
+        152.1779652373456
+        12.01816787810347
+        20.74501111108412
+        34.24344485181776
+        147.6059342336378
+ 2.38e+10    
+        153.1562504246502
+        34.69466510940741
+         152.763053760159
+        20.68677667792926
+        38.01841266652281
+        152.7550882862008
+        12.05038034661594
+        20.88157387168437
+        34.53757631840917
+        148.2197269880928
+ 2.39e+10    
+        153.7813517587215
+        34.98991334367848
+        153.3391587453756
+        20.82218689976411
+        38.27007534928184
+         153.332391033049
+        12.08134505475556
+        21.01754691993739
+        34.83241961500321
+        148.8337617372932
+ 2.4e+10     
+        154.4066856244471
+        35.28586746885138
+        153.9154406621202
+         20.9569940792729
+        38.52187002864461
+        153.9098853476778
+        12.11104914805123
+        21.15291965852144
+        35.12797391419293
+        149.4480427762734
+ 2.41e+10    
+        155.0322569097844
+        35.58252705881718
+        154.4919128675927
+        21.09118776566418
+        38.77379824053187
+        154.4875833937272
+         12.1394799920461
+        21.28768176465853
+        35.42423870120691
+        150.0625750144368
+ 2.42e+10    
+        155.6580710952703
+        35.87989198846142
+        155.0685889666308
+        21.22475778057403
+         39.0258617093565
+        155.0654976155344
+         12.1666251704432
+        21.42182318528272
+         35.7212137658856
+        150.6773639600652
+ 2.43e+10    
+        156.2841342390749
+        36.17796242581039
+        155.6454827991622
+        21.35769421325654
+           39.27806233992
+        155.6436407253152
+         12.1924724832302
+        21.55533413223952
+        36.01889919478451
+        151.2924157050671
+ 2.44e+10    
+        156.9104529622797
+         36.4767388243006
+        156.2226084279992
+        21.48998741580192
+        39.53040220952337
+        156.2220256906784
+        12.21700994478322
+         21.6882050775039
+        36.31729536339983
+        151.9077369099485
+ 2.45e+10    
+        157.5370344343703
+        36.77622191517288
+         156.799980126982
+        21.62162799837368
+        39.78288356028796
+        156.8006657224613
+        12.24022578195125
+        21.82042674842692
+        36.61640292851455
+          152.52333478901
+ 2.46e+10    
+        158.1638863589523
+        37.07641269998663
+        157.3776123694425
+        21.75260682447129
+        40.03550879167998
+        157.3795742628771
+        12.26210843212142
+         21.9519901230065
+        36.91622282066572
+        153.1392170957672
+ 2.47e+10    
+        158.7910169596723
+        37.37731244325513
+        157.9555198170036
+         21.8829150062221
+        40.28828045323646
+        157.9587649739776
+        12.28264654126783
+        22.08288642518788
+        37.21675623672988
+        153.7553921085956
+ 2.48e+10    
+        159.4184349663643
+        37.67892266519943
+         158.533717308683
+        22.01254389969812
+        40.54120123748525
+        158.5382517264098
+        12.30182896198317
+        22.21310712019154
+        37.51800463262564
+        154.3718686165905
+ 2.49e+10    
+        160.0461496013944
+        37.98124513461855
+        159.1122198503129
+        22.14148510026007
+        40.79427397305637
+        159.1180485884714
+        12.31964475149531
+        22.34264390987152
+        37.81996971613334
+        154.9886559056503
+ 2.5e+10     
+        160.6741705662255
+        38.28428186187632
+        159.6910426042544
+        22.26973043793533
+        41.04750161797865
+        159.6981698154523
+        12.33608316966957
+        22.47148872810394
+        38.12265343982739
+        155.6057637447691
+ 2.51e+10    
+        161.3025080281794
+        38.58803509200091
+        160.2702008794048
+        22.39727197282164
+        41.30088725315892
+        160.2786298392592
+        12.35113367699731
+        22.59963373620752
+        38.42605799412399
+        156.2232023725504
+ 2.52e+10    
+         161.931172607415
+        38.89250729789872
+        160.8497101214927
+        22.52410199052563
+        41.55443407603832
+        160.8594432583139
+        12.36478593257213
+        22.72707131839634
+        38.73018580043833
+        156.8409824839252
+ 2.53e+10    
+        162.5601753640964
+        39.19770117367649
+        161.4295859036488
+        22.65021299763051
+        41.80814539442164
+        161.4406248277187
+        12.37702979205468
+        22.85379407726732
+         39.0350395044542
+        157.4591152170844
+ 2.54e+10    
+        163.1895277857763
+        39.50361962807693
+        162.0098439172466
+        22.77559771719955
+        42.06202462047574
+        162.0221894496901
+        12.38785530562672
+        22.97979482931927
+        39.34062196950116
+        158.0776121406176
+ 2.55e+10    
+        163.8192417749648
+        39.81026577801948
+        162.5904999630133
+        22.90024908431434
+        42.31607526489444
+        162.6041521642443
+        12.39725271593558
+        23.10506660050909
+        39.64693627003989
+        158.6964852408537
+ 2.56e+10    
+        164.4493296369059
+        40.11764294224819
+          163.17156994239
+        23.02416024164403
+        42.57030093122277
+        163.1865281401359
+        12.40521245602969
+        23.22960262184409
+        39.95398568525433
+        159.3157469094103
+ 2.57e+10    
+        165.0798040675413
+        40.42575463508553
+        163.7530698491518
+        23.14732453505199
+        42.82470531034024
+        163.7693326660417
+        12.41172514728591
+        23.35339632500829
+        40.26177369274684
+        159.9354099309384
+ 2.58e+10    
+        165.7106781416718
+        40.73460456028985
+        164.3350157612686
+        23.26973550923994
+          43.079292175097
+        164.3525811419856
+        12.41678159733008
+        23.47644133802704
+        40.57030396233906
+        160.5554874710686
+ 2.59e+10    
+        166.3419653013053
+        41.04419660501451
+        164.9174238330031
+         23.3913869034277
+         43.3340653751008
+        164.9362890709968
+        12.42037279795098
+        23.59873148096912
+         40.8795803499729
+        161.1759930645524
+ 2.6e+10     
+        166.9736793441951
+        41.35453483386789
+         165.500310287249
+        23.51227264706874
+        43.58902883165054
+         165.520472050998
+        12.42248992300896
+        23.72026076168881
+        41.18960689171391
+        161.7969406035999
+ 2.61e+10    
+        167.6058344125658
+         41.6656234830742
+        166.0836914080908
+        23.63238685560737
+        43.84418653281191
+        166.1051457669163
+        12.42312432633932
+        23.84102337160096
+         41.5003877978525
+        162.4183443264051
+ 2.62e+10    
+        168.2384449820193
+         41.9774669547304
+        166.6675835335886
+        23.75172382627102
+        44.09954252863486
+        166.6903259830172
+        12.42226753965249
+        23.96101368150362
+        41.81192744710388
+        163.0402188058633
+ 2.63e+10    
+         168.871525850627
+        42.29006981116027
+        167.2520030487755
+        23.87027803390291
+        44.35510092650564
+         167.276028535447
+        12.41991127043033
+        24.08022623743302
+         42.1242303809052
+        163.6625789384784
+ 2.64e+10    
+        169.5050921281967
+        42.60343676936529
+        167.8369663788729
+        23.98804412683407
+        44.61086588663314
+          167.86226932499
+        12.41604739981978
+        24.19865575656078
+        42.43730129780682
+        164.2854399334504
+ 2.65e+10    
+        170.1391592257243
+        42.91757269556706
+        168.4224899827057
+        24.10501692279622
+        44.86684161766538
+        168.4490643100258
+        12.41066798052569
+        24.31629712313543
+        42.75114504795813
+        164.9088173019483
+ 2.66e+10    
+        170.7737428450125
+        43.23248259984357
+        169.0085903463202
+        24.22119140487201
+        45.12303237243261
+        169.0364294996926
+        12.40376523470089
+        24.43314538445685
+        43.06576662768659
+        165.5327268465652
+ 2.67e+10    
+        171.4088589684697
+        43.54817163085637
+        169.5952839767987
+         24.3365627174895
+        45.37944244381448
+        169.6243809472358
+         12.3953315518375
+        24.54919574689931
+        43.38117117416675
+        166.1571846509466
+ 2.68e+10    
+        172.0445238490762
+        43.86464507066738
+        170.1825873962656
+         24.4511261624553
+        45.63607616072925
+         170.212934743559
+        12.38535948665752
+        24.66444357197337
+        43.69736396018134
+        166.7822070696036
+ 2.69e+10    
+        172.6807540005217
+        44.18190832964418
+        170.7705171360764
+        24.56487719502951
+        45.89293788423991
+        170.8021070109548
+        12.37384175700426
+        24.77888437242677
+        44.01435038896892
+        167.4078107178912
+ 2.7e+10     
+        173.3175661875067
+        44.49996694145327
+        171.3590897311948
+        24.67781142004306
+        46.15003200377742
+        171.3919138970211
+        12.36077124173549
+        24.89251380839144
+        44.33213598916063
+        168.0340124621621
+ 2.71e+10    
+        173.9549774162132
+        44.81882655813712
+        171.9483217147383
+        24.78992458805438
+        46.40736293347442
+        171.9823715687519
+         12.3461409786186
+        25.00532768356991
+        44.65072640980287
+         168.660829410094
+ 2.72e+10    
+        174.5930049249326
+        45.13849294527848
+        172.5382296127068
+        24.90121259155246
+        46.66493510861178
+        172.5734962068078
+        12.32994416222851
+         25.1173219414658
+        44.97012741546401
+        169.2882789011753
+ 2.73e+10    
+        175.2316661748597
+        45.45897197724562
+        173.1288299388721
+        25.01167146119787
+        46.92275298217032
+        173.1653039999523
+        12.31217414184883
+        25.22849266165574
+        45.29034488142636
+        169.9163784973649
+ 2.74e+10    
+        175.8709788410419
+        45.78026963252169
+        173.7201391898329
+        25.12129736210802
+        47.18082102148877
+         173.757811139657
+         12.2928244193763
+        25.33883605610343
+        45.61138478895968
+        170.5451459739119
+ 2.75e+10    
+        176.5109608034841
+        46.10239198911262
+        174.3121738402353
+        25.23008659018569
+        47.43914370502358
+        174.3510338148708
+        12.27188864723063
+        25.44834846551903
+         45.9332532206764
+        171.1745993103337
+ 2.76e+10    
+        177.1516301384134
+         46.4253452200374
+         174.904950338145
+        25.33803556848852
+        47.69772551920876
+        174.9449882069409
+         12.2493606262683
+        25.55702635575929
+        46.25595635596591
+        171.8047566815554
+ 2.77e+10    
+         177.793005109689
+        46.74913558889377
+        175.4984851005711
+        25.44514084364278
+        47.95657095541384
+        175.5396904847003
+        12.22523430370187
+        25.66486631426961
+        46.57950046651001
+        172.4356364492071
+ 2.78e+10    
+        178.4351041603663
+        47.07376944550351
+        176.0927945091446
+         25.5513990823005
+        48.21568450699667
+        176.1351567996965
+         12.1995037710262
+        25.77186504657419
+        46.90389191187384
+         173.067257153074
+ 2.79e+10    
+        179.0779459044113
+        47.39925322163158
+        176.6878949059344
+        25.65680706763562
+        48.47507066644921
+        176.7314032815763
+        12.17216326194928
+        25.87801937280347
+        47.22913713517445
+         173.699637502698
+ 2.8e+10     
+        179.7215491185574
+          47.725593426783
+        177.2838025894133
+        25.76136169589078
+        48.73473392263426
+        177.3284460336089
+        12.14320715033177
+        25.98332622426692
+        47.55524265882448
+        174.3327963691327
+ 2.81e+10    
+        180.3659327343072
+        48.05279664406997
+        177.8805338105537
+        25.86505997295731
+        48.99467875811125
+        177.9263011283576
+        12.11262994813246
+        26.08778264007201
+        47.88221508035113
+        174.9667527768454
+ 2.82e+10    
+        181.0111158300806
+        48.38086952615348
+         178.478104769062
+        25.96789901100763
+        49.25490964654786
+        178.5249846034835
+        12.08042630336229
+        26.19138576378077
+        48.21006106828623
+        175.6015258957628
+ 2.83e+10    
+        181.6571176234995
+        48.70981879125719
+        179.0765316097459
+         26.0698760251654
+        49.51543105021683
+        179.1245124576891
+        12.04659099804642
+        26.29413284011352
+        48.53878735813038
+        176.2371350334679
+ 2.84e+10    
+        182.3039574638114
+         49.0396512192485
+        179.6758304190066
+        26.17098833021811
+        49.77624741757423
+        179.7249006467893
+        12.01111894619441
+        26.39602121169487
+         48.8684007483872
+        176.8735996275316
+ 2.85e+10    
+         182.951654824452
+        49.37037364779274
+        180.2760172214556
+        26.27123333737734
+        50.03736318091956
+        180.3261650799165
+        11.97400519178048
+         26.4970483158421
+        49.19890809666701
+         177.510939237989
+ 2.86e+10    
+        183.6002292957415
+        49.70199296857159
+        180.8771079766545
+        26.37060855107674
+        50.29878275413293
+        180.9283216158461
+        11.93524490673197
+        26.59721168139652
+        49.53031631586105
+        178.1491735399543
+ 2.87e+10    
+        184.2497005777108
+        50.03451612357235
+        181.4791185759767
+        26.46911156581666
+        50.56051053049057
+        181.5313860594518
+        11.89483338892846
+        26.69650892559837
+        49.86263237038027
+        178.7883223163696
+ 2.88e+10    
+        184.9000884730663
+        50.36795010143992
+        182.0820648395763
+        26.56674006304971
+        50.82255088055339
+         182.135374158275
+        11.85276606021091
+        26.79493775100484
+        50.19586327246545
+        179.4284054508939
+ 2.89e+10    
+        185.5514128802746
+        50.70230193389565
+        182.6859625134769
+        26.66349180810851
+        51.08490815012964
+        182.7403015992136
+        11.80903846440052
+        26.89249594244712
+        50.53001607855762
+        180.0694429209139
+ 2.9e+10     
+         186.203693786784
+        51.03757869221916
+        183.2908272667682
+        26.75936464717903
+        51.34758665830892
+        183.3461840053275
+         11.7636462653302
+         26.9891813640381
+        50.86509788573807
+        180.7114547906995
+ 2.91e+10    
+         186.856951262362
+         51.3737874837953
+        183.8966746889114
+        26.85435650431215
+        51.61059069556509
+        183.9530369327522
+        11.71658524488512
+        27.08499195621253
+        51.20111582822862
+        181.3544612046773
+ 2.92e+10    
+        187.5112054525689
+        51.71093544871896
+        184.5035202871424
+        26.94846537848237
+        51.87392452192768
+        184.5608758677271
+        11.66785130105665
+        27.17992573281679
+        51.53807707395629
+         181.998482380837
+ 2.93e+10    
+        188.1664765723395
+        52.04902975646531
+        185.1113794839881
+        27.04168934068245
+        52.13759236521881
+        185.1697162237248
+        11.61744044600655
+        27.27398077823761
+        51.87598882117947
+        182.6435386042625
+ 2.94e+10    
+        188.8227848996964
+         52.3880776026166
+        185.7202676148695
+        27.13402653106763
+        52.40159841935542
+        185.7795733386887
+        11.56534880414473
+        27.36715524457387
+        52.21485829517392
+        183.2896502207825
+ 2.95e+10    
+        189.4801507695785
+        52.72808620565005
+        186.3301999258115
+        27.22547515613632
+         52.6659468427146
+        186.3904624723708
+        11.51157261021852
+        27.45944734884919
+        52.55469274498053
+        183.9368376307507
+ 2.96e+10    
+        190.1385945677831
+        53.06906280378376
+        186.9411915712426
+         27.3160334859525
+         52.9306417565595
+        187.0023988037698
+        11.45610820741458
+        27.55085537026734
+        52.89549944020873
+         184.585121282935
+ 2.97e+10    
+        190.7981367250299
+        53.41101465187821
+        187.5532576118849
+        27.40569985141402
+        53.19568724352597
+        187.6153974286645
+        11.39895204547459
+        27.64137764750752
+        53.23728566790211
+         185.234521668539
+ 2.98e+10    
+        191.4587977111348
+        53.75394901839608
+        188.1664130127391
+        27.49447264155809
+         53.4610873461687
+        188.2294733572454
+        11.34010067882339
+         27.7310125760628
+        53.58005872945741
+        185.8850593153259
+ 2.99e+10    
+        192.1205980292925
+        54.09787318241616
+        188.7806726411489
+        27.58235030090771
+        53.72684606556218
+        188.8446415118346
+        11.27955076471077
+        27.81975860561791
+        53.92382593760138
+        186.5367547818691
+ 3e+10       
+        192.7835582104816
+        54.44279443070302
+        189.3960512649599
+        27.66933132686549
+        53.99296735995984
+        189.4609167247001
+        11.21729906136759
+        27.90761423746855
+        54.26859461342319
+         187.189628651907
+ 3.01e+10    
+        193.4476988079631
+        54.78872005482839
+        190.0125635507514
+        27.75541426713748
+        54.25945514350549
+        190.0783137359542
+        11.15334242617465
+        27.99457802198127
+        54.61437208345964
+        187.8437015288159
+ 3.02e+10    
+        194.1130403918984
+        55.13565734834781
+        190.6302240621582
+        27.84059771720743
+        54.52631328499959
+        190.6968471915415
+        11.08767781384702
+         28.0806485560926
+         54.9611656768369
+        188.4989940301897
+ 3.03e+10    
+        194.7796035440672
+        55.48361360402724
+        191.2490472582628
+        27.92488031784566
+        54.79354560671617
+        191.3165316413093
+        11.02030227463194
+        28.16582448085169
+        55.30898272246106
+         189.155526782529
+ 3.04e+10    
+        195.4474088526929
+         55.8325961111218
+        191.8690474920713
+         28.0082607526592
+        55.06115588327039
+        191.9373815371598
+        10.95121295252131
+        28.25010447899725
+        55.65783054626414
+        189.8133204160364
+ 3.05e+10    
+        196.1164769073682
+        56.18261215270533
+        192.4902390090588
+        28.09073774568467
+        55.32914784053592
+         192.559411231281
+        10.88040708347998
+        28.33348727258047
+         56.0077164684994
+        190.4723955595191
+ 3.06e+10    
+        196.7868282940811
+        56.53366900304802
+        193.1126359457887
+        28.17231005901477
+        55.59752515460949
+        193.1826349744628
+        10.80788199368714
+        28.41597162062026
+        56.35864780108741
+        191.1327728353925
+ 3.07e+10    
+        197.4584835903498
+        56.88577392504462
+        193.7362523286056
+        28.25297649047005
+        55.86629145082265
+        193.8070669144757
+          10.733635097795
+        28.49755631680631
+        56.71063184501123
+        191.7944728547858
+ 3.08e+10    
+        198.1314633604415
+        57.23893416768879
+        194.3611020723934
+        28.33273587130646
+        56.13545030279968
+        194.4327210945375
+        10.65766389720107
+        28.57824018723161
+        57.06367588776087
+         192.457516212755
+ 3.09e+10    
+        198.8057881507017
+        57.59315696359667
+        194.9871989794018
+        28.41158706396277
+          56.405005231559
+        195.0596114518447
+        10.57996597833687
+        28.65802208817043
+        57.41778720082539
+        193.1219234835829
+ 3.1e+10     
+        199.4814784849713
+        57.94844952657563
+         195.614556738139
+        28.48952895984589
+        56.67495970465929
+        195.6877518161781
+        10.50053901097217
+        28.73690090389236
+        57.77297303723306
+        193.7877152161914
+ 3.11e+10    
+        200.1585548601011
+        58.30481904923926
+         196.243188922329
+        28.56656047715521
+        56.94531713538682
+        196.3171559085728
+        10.41938074653481
+        28.81487554451461
+        58.12924062913658
+        194.4549119296379
+ 3.12e+10    
+         200.837037741557
+        58.66227270066641
+        196.8731089899255
+        28.64268055874518
+         57.2160808819846
+        196.9478373400623
+        10.33648901644621
+        28.89194494388897
+        58.48659718544504
+        195.1235341087144
+ 3.13e+10    
+        201.5169475591215
+        59.02081762410722
+        197.5043302821947
+        28.71788817002354
+        57.48725424692184
+        197.5798096104803
+        10.25186173047399
+        28.96810805753395
+        58.84504988950093
+        195.7936021996371
+ 3.14e+10    
+         202.198304702679
+        59.38046093472988
+        198.1368660228456
+        28.79218229689064
+        57.75884047620261
+        198.2130861073355
+        10.16549687509947
+        29.04336386059557
+         59.2046058968011
+        196.4651366058271
+ 3.15e+10    
+        202.8811295180955
+         59.7412097174121
+        198.7707293172316
+        28.86556194371395
+        58.03084275871284
+        198.8476801047413
+        10.07739251190268
+         29.1177113458504
+         59.5652723327625
+        197.1381576837882
+ 3.16e+10    
+        203.5654423031843
+        60.10307102457411
+        199.4059331515941
+        28.93802613133614
+        58.30326422560402
+        199.4836047624054
+        9.987546775962613
+        29.19114952174403
+        59.92705629052835
+        197.8126857390639
+ 3.17e+10    
+        204.2512633037556
+        60.46605187405366
+        200.0424903923671
+        29.00957389512766
+        58.57610794971416
+        200.1208731246891
+        9.895957874275476
+        29.26367741046522
+        60.28996482882061
+        198.4887410222932
+ 3.18e+10    
+        204.9386127097559
+        60.83015924702273
+         200.680413785537
+        29.08020428306943
+        58.84937694502424
+        200.7594981197117
+        9.802624084188295
+         29.3352940460569
+        60.65400496982956
+        199.1663437253465
+ 3.19e+10    
+        205.6275106514859
+        61.19540008594241
+        201.3197159560456
+        29.14991635387223
+        59.12307416614812
+        201.3994925585211
+        9.707543751849878
+        29.40599847256242
+        61.01918369714903
+         199.845513977551
+ 3.2e+10     
+        206.3179771959102
+        61.56178129256028
+        201.9604094072479
+        29.21870917513522
+        59.39720250785692
+        202.0408691343113
+        9.610715290678833
+        29.47578974220794
+        61.38550795374805
+        200.5262718419979
+ 3.21e+10    
+        207.0100323430344
+        61.92930972594466
+        202.6025065204207
+        29.28658182153568
+         59.6717648046363
+        202.6836404216991
+        9.512137179847926
+        29.54466691362036
+        61.75298463998476
+        201.2086373119344
+ 3.22e+10    
+        207.7036960223793
+        62.29799220056002
+        203.2460195543129
+        29.35353337305814
+        59.94676383027569
+        203.3278188760526
+        9.411807962786021
+        29.61262905007797
+        62.12162061165893
+        201.8926303072364
+ 3.23e+10    
+        208.3989880895201
+        62.66783548437583
+        203.8909606447451
+        29.41956291325509
+         60.2222022974881
+        203.9734168328647
+        9.309726245696918
+        29.67967521779929
+        62.49142267810259
+        202.5782706709657
+ 3.24e+10    
+        209.0959283227114
+        63.03884629701903
+        204.5373418042538
+        29.48466952754404
+        60.49808285756134
+        204.6204465071848
+        9.205890696094968
+        29.74580448426275
+        62.86239760030886
+        203.2655781660002
+ 3.25e+10    
+         209.794536419587
+        63.41103130795647
+        205.1851749217731
+        29.54885230153969
+        60.77440810003773
+        205.2689199930915
+        9.100300041359072
+        29.81101591656367
+        63.23455208909875
+         203.954572471749
+ 3.26e+10    
+        210.4948319939388
+        63.78439713472022
+         205.834471762372
+        29.61211031941648
+        61.05118055242327
+        205.9188492632145
+        8.992953067302368
+        29.87530857980202
+         63.6078928033243
+        204.6452731809432
+ 3.27e+10    
+        211.1968345725624
+        64.15895034116262
+        206.4852439670147
+         29.6744426623098
+        61.32840267992506
+        206.5702461683053
+        8.883848616760702
+        29.93868153550636
+        63.98242634810804
+        205.3376997964991
+ 3.28e+10    
+        211.9005635921863
+        64.53469743575134
+        207.1375030523775
+        29.73584840674807
+        61.60607688521554
+        207.2231224368454
+        8.772985588197738
+        30.00113384008808
+        64.35815927311782
+        206.0318717284613
+ 3.29e+10    
+         212.606038396468
+        64.91164486989526
+        207.7912604106927
+        29.79632662311756
+        61.88420550822414
+        207.8774896747082
+        8.660362934327699
+        30.06266454333172
+        64.73509807087807
+        206.7278082910166
+ 3.3e+10     
+        213.3132782330623
+        65.28979903630778
+        208.4465273096349
+        29.85587637416107
+        62.16279082595341
+        208.5333593648494
+        8.545979660755961
+        30.12327268691632
+        65.11324917511513
+         207.425528699586
+ 3.31e+10    
+        214.0223022507605
+        65.66916626740017
+        209.1033148922425
+         29.9144967135099
+        62.44183505232268
+        209.1907428670526
+        8.429834824636457
+        30.18295730296757
+        65.49261895913543
+        208.1250520679789
+ 3.32e+10    
+        214.7331294967022
+        66.04975283371189
+        209.7616341768788
+         29.9721866842457
+        62.72134033803437
+        209.8496514177035
+        8.311927533347458
+        30.24171741264519
+        65.87321373423984
+        208.8263974056288
+ 3.33e+10    
+        215.4457789136495
+        66.43156494237022
+        210.4214960572195
+        30.02894531749835
+        63.00130877046539
+        210.5100961296126
+        8.192256943184704
+        30.29955202476024
+        66.25503974816924
+        209.5295836148913
+ 3.34e+10    
+        216.1602693373378
+        66.81460873558366
+        211.0829113022802
+         30.0847716310705
+        63.28174237358141
+        211.1720879918656
+         8.07082225807164
+        30.35646013442244
+        66.63810318358401
+        210.2346294884164
+ 3.35e+10    
+         216.876619493882
+        67.19889028916747
+        211.7458905564747
+        30.13966462809823
+        63.56264310787388
+        211.8356378697204
+        7.947622728288433
+        30.41244072172298
+        67.02241015657424
+        210.9415537065833
+ 3.36e+10    
+        217.5948479972608
+        67.58441561109801
+        212.4104443397016
+        30.19362329574072
+         63.8440128703198
+        212.5007565045321
+         7.82265764921787
+        30.46749275044301
+        67.40796671520397
+        211.6503748350062
+ 3.37e+10    
+        218.3149733468535
+        67.97119064010101
+        213.0765830474679
+        30.24664660389992
+        64.12585349436191
+        213.1674545137168
+        7.695926360108906
+        30.52161516679713
+        67.79477883808332
+        212.3611113221032
+ 3.38e+10    
+        219.0370139250537
+        68.35922124426833
+         213.744316951036
+        30.29873350397276
+        64.40816674991106
+        213.8357423907503
+         7.56742824285875
+        30.57480689820378
+        68.18285243297623
+        213.0737814967339
+ 3.39e+10    
+         219.760987994934
+        68.74851321970409
+        214.4136561976025
+        30.34988292763341
+        64.69095434336835
+        214.5056305051962
+        7.437162720811934
+        30.62706685208861
+        68.57219333543324
+        213.7884035658959
+ 3.4e+10     
+        220.4869136979803
+        69.13907228920162
+        215.0846108105039
+        30.40009378564426
+        64.97421791766746
+        215.1771291027684
+        7.305129257577441
+        30.67839391471475
+        68.96280730745829
+        214.5049956124875
+ 3.41e+10    
+         221.214809051886
+        69.53090410094872
+        215.7571906894522
+        30.44936496669739
+        65.25795905233556
+        215.8502483054227
+        7.171327355863708
+        30.72878695004535
+         69.3547000362037
+        215.2235755931353
+ 3.42e+10    
+        221.9446919484046
+        69.92401422726161
+          216.43140561079
+        30.49769533628626
+        65.54217926357414
+         216.524998111481
+        7.035756556331192
+        30.77824479863245
+        69.74787713269259
+        215.9441613360747
+ 3.43e+10    
+        222.6765801512631
+        70.31840816334692
+        217.1072652277795
+        30.54508373560505
+         65.8268800043581
+        217.2013883957863
+        6.898416436463044
+        30.82676627653789
+        70.14234413057412
+        216.6667705391017
+ 3.44e+10    
+        223.4104912941377
+        70.71409132609284
+        217.7847790709101
+        30.59152898047947
+        66.11206266455086
+        217.8794289098769
+        6.759306609453219
+        30.87435017427972
+        70.53810648490185
+        217.3914207675752
+ 3.45e+10    
+        224.1464428786778
+        71.11106905288476
+        218.4639565482319
+        30.63702986032209
+        66.39772857104008
+        218.5591292822029
+        6.618426723112457
+        30.92099525580923
+        70.93516957094488
+        218.1181294524825
+ 3.46e+10    
+        224.8844522726021
+        71.50934660045155
+        219.1448069457128
+        30.68158513712091
+        66.68387898788654
+        219.2404990183566
+         6.47577645879236
+        30.96670025751498
+        71.33353868302237
+        218.8469138885617
+ 3.47e+10    
+        225.6245367078327
+        71.90892914373563
+        219.8273394276149
+        30.72519354445307
+        66.97051511649232
+        219.9235475013343
+        6.331355530326903
+        31.01146388725543
+        71.73321903336826
+        219.5777912324828
+ 3.48e+10    
+        226.3667132787031
+         72.3098217747912
+        220.5115630369012
+        30.76785378652555
+        67.25763809578417
+        220.6082839918259
+        6.185163682991618
+        31.05528482341781
+         72.1342157510214
+        220.3107785010815
+ 3.49e+10    
+         227.110998940208
+         72.7120295017082
+        221.1974866956509
+        30.80956453724695
+        67.54524900241128
+        221.2947176285259
+        6.037200692481067
+        31.09816171400564
+        72.53653388074262
+        221.0458925696518
+ 3.5e+10     
+        227.8574105063128
+        73.11555724756039
+         221.885119205503
+        30.85032443932327
+        67.83334885095914
+        221.9828574284662
+        5.887466363903556
+         31.1400931757528
+        72.94017838195681
+        221.7831501702944
+ 3.51e+10    
+        228.6059646483157
+        73.52040984938024
+        222.5744692481194
+        30.89013210338298
+        68.12193859417872
+        222.6727122873783
+        5.735960530793745
+        31.18107779326356
+         73.3451541277224
+        222.5225678903126
+ 3.52e+10    
+        229.3566778932624
+         73.9265920571596
+        223.2655453856662
+        30.92898610712702
+        68.41101912322861
+        223.3642909800706
+        5.582683054143004
+        31.22111411818084
+        73.75146590372412
+        223.2641621706676
+ 3.53e+10    
+        230.1095666224115
+        74.33410853287278
+        223.9583560613096
+         30.9668849945067
+        68.70059126793136
+         224.057602160835
+        5.427633821447614
+        31.26020066837924
+        74.15911840729356
+        224.0079493044869
+ 3.54e+10    
+        230.8646470697534
+        74.74296384952407
+        224.6529095997341
+        31.00382727492702
+        68.99065579704404
+        224.7526543638676
+        5.270812745773995
+        31.29833592718328
+        74.56811624645131
+        224.7539454356174
+ 3.55e+10    
+        231.6219353205771
+        75.15316249022314
+        225.3492142076795
+        31.03981142247664
+        69.28121341854131
+        225.4494560037142
+        5.112219764842708
+         31.3355183426146
+        74.97846393897619
+        225.5021665572401
+ 3.56e+10    
+        232.3814473100892
+         75.5647088472774
+        226.0472779744844
+        31.07483587518377
+        69.57226477991092
+        226.1480153757363
+        4.951854840128963
+        31.37174632666074
+        75.39016591149669
+        226.2526285105224
+ 3.57e+10    
+        233.1431988220817
+        75.97760722131535
+        226.7471088726613
+        31.10889903429602
+        69.86381046846309
+        226.8483406565905
+        4.789717955981516
+        31.40701825457263
+        75.80322649860778
+        227.0053469833312
+ 3.58e+10    
+        233.9072054876459
+        76.39186182042687
+         227.448714758473
+        31.14199926358765
+        70.15585101164898
+        227.5504399047323
+        4.625809118758688
+        31.44133246418325
+        76.21764994200957
+        227.7603375089914
+ 3.59e+10    
+        234.6734827839371
+        76.80747675932943
+        228.1521033725303
+         31.1741348886902
+        70.44838687739505
+        228.2543210609381
+        4.460128355982157
+        31.47468725525512
+        76.63344038967007
+        228.5176154650877
+ 3.6e+10     
+        235.4420460329871
+        77.22445605855663
+        228.8572823404062
+        31.20530419644832
+        70.74141847444456
+         228.959991948839
+        4.292675715508253
+          31.507080888849
+        77.05060189501117
+        229.2771960723209
+ 3.61e+10    
+        236.2129104005575
+        77.64280364366807
+        229.5642591732588
+        31.23550543430058
+        71.03494615271322
+        229.6674602754761
+         4.12345126471676
+        31.53851158671841
+        77.46913841611665
+        230.0390943934108
+ 3.62e+10    
+        236.9860908950478
+        78.06252334448179
+        230.2730412684696
+        31.26473680968406
+        71.32897020365334
+        230.3767336318721
+         3.95245508971696
+        31.56897753072745
+        77.88905381496249
+         230.803325332038
+ 3.63e+10    
+        237.7616023664414
+        78.48361889432961
+        230.9836359102993
+        31.29299648946316
+         71.6234908606304
+        231.0878194936167
+        3.779687294571591
+        31.59847686229315
+        78.31035185666991
+        231.5699036318409
+ 3.64e+10    
+        238.5394595053014
+        78.90609392933085
+        231.6960502705458
+        31.32028259938195
+        71.91850829930785
+        231.8007252214662
+        3.605148000537669
+        31.62700768185076
+          78.733036208779
+        232.3388438754509
+ 3.65e+10    
+        239.3196768418056
+        79.32995198769071
+        232.4102914092249
+        31.34659322354034
+        72.21402263804298
+        232.5154580619632
+        3.428837345324997
+        31.65456804834186
+        79.15711044054562
+        233.1101604835772
+ 3.66e+10    
+        240.1022687448329
+        79.75519650901818
+        233.1263662752577
+        31.37192640389313
+        72.51003393829217
+        233.2320251480627
+        3.250755482372011
+        31.68115597872668
+        79.58257802225847
+        233.8838677141306
+ 3.67e+10    
+        240.8872494210829
+        80.18183083366431
+        233.8442817071661
+        31.39628013977311
+        72.80654220502413
+        233.9504334997805
+        3.070902580138563
+        31.70676944751755
+        80.00944232457681
+        234.6599796613951
+ 3.68e+10    
+        241.6746329142463
+        80.60985820208116
+         234.564044433786
+        31.41965238743606
+         73.1035473871442
+        234.6706900248458
+         2.88927882141661
+        31.73140638633717
+        80.43770661789071
+        235.4385102552385
+ 3.69e+10    
+        242.4644331042133
+        81.03928175420262
+        235.2856610749839
+        31.44204105962805
+        73.40104937792563
+        235.3928015193758
+        2.705884402657297
+          31.755064683497
+        80.86737407169963
+        236.2194732603685
+ 3.7e+10     
+        243.2566637063258
+        81.47010452884314
+        236.0091381423898
+        31.46344402517735
+        73.69904801544982
+         236.116774668554
+        2.520719533316168
+        31.77774218359955
+        81.29844775401406
+        237.0028822756276
+ 3.71e+10    
+        244.0513382706654
+        81.90232946311727
+         236.734482040132
+        31.48385910860471
+        73.99754308305549
+        236.8426160473282
+         2.33378443521439
+        31.79943668716038
+        81.73093063077384
+        237.7887507333303
+ 3.72e+10    
+          244.84847018139
+        82.33595939187951
+        237.4616990655893
+        31.50328408975961
+        74.29653430979428
+        237.5703321211135
+        2.145079341918176
+        31.82014595025496
+         82.1648255652904
+        238.5770918986425
+ 3.73e+10    
+        245.6480726561009
+        82.77099704718239
+        238.1907954101441
+        31.52171670347551
+        74.59602137089524
+         238.299929246509
+        1.954604498134518
+        31.83986768418337
+        82.60013531770581
+        239.3679188689977
+ 3.74e+10    
+        246.4501587452587
+        83.20744505775443
+          238.92177715995
+        31.53915463924785
+        74.89600388823673
+        239.0314136720267
+        1.762360159124209
+        31.85859955515915
+        83.03686254447122
+         240.161244573553
+ 3.75e+10    
+        247.2547413316319
+        83.64530594849819
+        239.6546502967032
+        31.55559554093258
+          75.196481430825
+        239.7647915388299
+        1.568346590131861
+        31.87633918401769
+        83.47500979784772
+        240.9570817726898
+ 3.76e+10    
+        248.0618331297828
+        84.08458214000427
+        240.3894206984245
+         31.5710370064664
+        75.49745351527969
+        240.5000688814761
+        1.372564065832714
+        31.89308414594576
+        83.91457952542217
+        241.7554430575424
+ 3.77e+10    
+        248.8714466855994
+        84.52527594808801
+        241.1260941402486
+        31.58547658760765
+        75.79891960632737
+        241.2372516286789
+         1.17501286979635
+        31.90883197023105
+        84.35557406964467
+        242.5563408495746
+ 3.78e+10    
+        249.6835943758527
+        84.96738958334016
+        241.8646762952128
+        31.59891178969739
+        76.10087911729974
+        241.9763456040706
+       0.9756932939672804
+        31.92358014003348
+        84.79799566738394
+        243.3597874001902
+ 3.79e+10    
+         250.498288407804
+        85.41092515070039
+         242.605172735066
+         31.6113400714417
+        76.40333141063984
+        242.7173565269792
+       0.7746056381624582
+        31.93732609217536
+        85.24184644950195
+         244.165794790377
+ 3.8e+10     
+        251.3155408188392
+        85.85588464904571
+        243.3475889310732
+        31.62275884471384
+        76.70627579841366
+        243.4602900132089
+       0.5717502095851001
+        31.95006721695206
+         85.6871284404443
+         244.974374930391
+ 3.81e+10    
+        252.1353634761424
+        86.30226997079774
+        244.0919302548291
+        31.63316547437595
+        77.00971154282854
+        244.2051515758329
+       0.3671273223558682
+        31.96180085796269
+        86.13384355785324
+        245.7855395594799
+ 3.82e+10    
+        252.9577680764049
+        86.75008290154834
+        244.8382019790788
+        31.64255727812153
+        77.31363785675498
+        244.9519466259916
+       0.1607372970598284
+        31.97252431195924
+        86.58199361219344
+        246.5993002456323
+ 3.83e+10    
+         253.782766145572
+        87.19932511970315
+        245.5864092785432
+        31.65093152633643
+        77.61805390425798
+         245.700680473699
+     -0.04741953968916768
+        31.98223482871644
+        87.03158030640064
+        247.4156683853725
+ 3.84e+10    
+        254.6103690386192
+        87.64999819614039
+         246.336557230749
+        31.65828544198008
+        77.92295880112954
+        246.4513583286534
+       -0.257342855668111
+        31.99092961091979
+         87.4826052355433
+        248.2346552035838
+ 3.85e+10    
+        255.4405879393668
+        88.10210359389015
+        247.0886508168637
+        31.66461620048559
+        78.22835161543051
+        247.2039853010634
+      -0.4690323134477241
+        31.99860581407339
+        87.93506988650657
+        249.0562717533671
+ 3.86e+10    
+        256.2734338603293
+        88.55564266782841
+        247.8426949225356
+        31.66992092967927
+        78.53423136803312
+        247.9585664024627
+      -0.6824875707788358
+        32.00526054642538
+        88.38897563768832
+        249.8805289159361
+ 3.87e+10    
+         257.108917642592
+        89.01061666438909
+        248.5986943387396
+        31.67419670971774
+        78.84059703317291
+        248.7151065465573
+      -0.8977082809627612
+        32.01089086891319
+        88.84432375871778
+        250.7074374005414
+ 3.88e+10    
+        257.9470499557304
+        89.46702672129287
+        249.3566537626239
+        31.67744057304544
+        79.14744753900221
+        249.4736105500513
+       -1.114694093204893
+        32.01549379512588
+        89.30111541018601
+        251.5370077444317
+ 3.89e+10    
+        258.7878412977533
+        89.92487386729331
+        250.1165777983636
+        31.67964950436871
+        79.45478176814873
+        250.2340831334973
+       -1.333444652952274
+        32.01906629128616
+        89.75935164339738
+        252.3692503128431
+ 3.9e+10     
+        259.6313019950822
+        90.38415902193779
+        250.8784709580171
+        31.68082044064982
+        79.76259855828033
+        250.9965289221419
+       -1.553959602214698
+        32.02160527624895
+        90.21903340013625
+        253.2041752990302
+ 3.91e+10    
+        260.4774422025652
+         90.8448829953477
+         251.642337662385
+        31.68095027111813
+        80.07089670267152
+        251.7609524467829
+       -1.776238579870012
+        32.02310762151814
+        90.68016151244908
+         254.041792724311
+ 3.92e+10    
+        261.3262719035181
+        91.30704648801225
+        252.4081822418736
+        31.68003583729809
+        80.37967495077643
+        252.5273581446271
+       -2.000281221952922
+        32.02357015128203
+        91.14273670244593
+        254.8821124381659
+ 3.93e+10    
+        262.1778009097974
+        91.77065009060048
+        253.1760089373626
+        31.67807393305777
+        80.68893200880385
+         253.295750360152
+       -2.226087161927938
+         32.0229896424643
+        91.60675958211398
+        255.7251441183453
+ 3.94e+10    
+        263.0320388619062
+        92.23569428378774
+        253.9458219010681
+        31.67506130467182
+        80.99866654029734
+        254.0661333459758
+       -2.453656030946143
+        32.02136282479416
+        92.07223065315291
+         256.570897271029
+ 3.95e+10    
+        263.8889952291289
+        92.70217943809942
+        254.7176251974216
+        31.67099465090288
+        81.30887716671883
+        254.8385112637285
+       -2.682987458086386
+        32.01868638089183
+        92.53915030682106
+        257.4193812309968
+ 3.96e+10    
+         264.748679309699
+        93.17010581377151
+        255.4914228039399
+        31.66587062310124
+        81.61956246803473
+        255.6128881849261
+       -2.914081070579773
+        32.01495694637203
+        93.00751882380104
+        258.2706051618437
+ 3.97e+10    
+        265.6111002309901
+        93.63947356062258
+        256.2672186121013
+        31.65968582531985
+        81.93072098330782
+        256.3892680918535
+         -3.1469364940194
+        32.01017110996391
+        93.47733637407859
+        259.1245780562118
+ 3.98e+10    
+         266.476266949745
+        94.11028271794746
+        257.0450164282245
+        31.65243681444607
+         82.2423512112893
+        257.1676548784424
+       -3.381553352553289
+        32.00432541364705
+        93.94860301684091
+        259.9813087360671
+ 3.99e+10    
+        267.3441882523271
+        94.58253321442157
+        257.8248199743502
+        31.64412010035154
+         82.5544516110171
+        257.9480523511594
+       -3.617931269062182
+        31.99741635280478
+        94.42131870038607
+        260.8408058529865
+ 4e+10       
+         268.214872755001
+        95.05622486802264
+        258.6066328891186
+        31.63473214605654
+         82.8670206024149
+        258.7304642298955
+       -3.856069865321685
+        31.98944037639193
+        94.89548326205087
+        261.7030778884899
+ 4.01e+10    
+        269.0883289042485
+        95.53135738596836
+        259.3904587286601
+        31.62426936791189
+         83.1800565668961
+         259.514894148857
+       -4.095968762148269
+        31.98039388712075
+        95.37109642815456
+        262.5681331543911
+ 4.02e+10    
+        269.9645649771057
+         96.0079303646683
+        260.1763009674734
+        31.61272813579651
+        83.49355784796855
+        260.3013456574595
+       -4.337627579530216
+        31.97027324166114
+        95.84815781395521
+        263.4359797931775
+ 4.03e+10    
+        270.8435890815276
+        96.48594328969074
+         260.964162999316
+        31.60010477333065
+        83.80752275184393
+        261.0898222212229
+       -4.581045936743139
+        31.95907475085598
+        96.32666692362351
+        264.3066257784193
+ 4.04e+10    
+        271.7254091567834
+        96.96539553574539
+        261.7540481380869
+        31.58639555810437
+        84.12194954804811
+        261.8803272226738
+       -4.826223452449427
+        31.94679467995497
+        96.80662315023123
+        265.1800789152065
+ 4.05e+10    
+        272.6100329738813
+        97.44628636668044
+        262.5459596187212
+        31.57159672192306
+        84.43683647003537
+        262.6728639622406
+       -5.073159744783115
+         31.9334292488593
+        97.28802577575384
+        266.0563468406086
+ 4.06e+10    
+        273.4974681360147
+        97.92861493549546
+        263.3399005980748
+        31.55570445106659
+        84.75218171580478
+        263.4674356591635
+       -5.321854431418986
+        31.91897463238532
+         97.7708739710891
+        266.9354370241648
+ 4.07e+10    
+        274.3877220790358
+        98.41238028436783
+        264.1358741558155
+        31.53871488656469
+        85.06798344851789
+         264.264045452393
+       -5.572307129626338
+        31.90342696054113
+        98.25516679609068
+        267.8173567684007
+ 4.08e+10    
+          275.28080207196
+        98.89758134469371
+        264.9338832953115
+        31.52062412448682
+        85.38423979711935
+        265.0626964014969
+       -5.824517456307977
+         31.8867823188182
+        98.74090319961455
+        268.7021132093666
+ 4.09e+10    
+         276.176715217491
+        99.38421693714605
+        265.7339309445263
+        31.50142821624739
+        85.70094885696093
+        265.8633914875714
+       -6.078485028023684
+         31.8690367484987
+         99.2280820195832
+        269.5897133172043
+ 4.1e+10     
+        277.0754684525758
+         99.8722857717442
+         266.536019956905
+        31.48112316892492
+        86.01810869042453
+        266.6661336141431
+       -6.334209460998863
+        31.85018624697559
+        99.71670198306111
+        270.4801638967413
+ 4.11e+10    
+        277.9770685489809
+        100.3617864479391
+        267.3401531122683
+        31.45970494559631
+        86.33571732754973
+        267.4709256080843
+       -6.591690371118277
+        31.83022676808799
+        100.2067617063472
+        271.3734715881044
+ 4.12e+10    
+        278.8815221138992
+        100.8527174547135
+        268.1463331177039
+        31.43716946568507
+        86.65377276666301
+        268.2777702205209
+       -6.850927373904442
+        31.80915422247131
+        100.6982596950812
+        272.2696428673655
+ 4.13e+10    
+        279.7888355905736
+        101.3450771706961
+        268.9545626084572
+        31.41351260532441
+        86.97227297500727
+        269.0866701277443
+       -7.111920084481751
+        31.78696447792003
+         101.191194344362
+        273.1686840472003
+ 4.14e+10    
+        280.6990152589572
+          101.83886386429
+        269.7648441488224
+         31.3887301977331
+        87.29121588937394
+        269.8976279321229
+        -7.37466811752537
+        31.76365335976435
+        101.6855639388852
+        274.0706012775874
+ 4.15e+10    
+        281.6120672363834
+        102.3340756938139
+        270.5771802330333
+        31.36281803360631
+        87.61059941673696
+        270.7106461630179
+       -7.639171087195512
+        31.73921665126225
+        102.1813666530903
+        274.9754005465165
+ 4.16e+10    
+        282.5279974782744
+        102.8307107076608
+        271.3915732861554
+         31.3357718615201
+        87.93042143488803
+        271.5257272776904
+       -7.905428607057079
+        31.71365009400311
+        102.6786005513232
+        275.8830876807259
+ 4.17e+10    
+        283.4468117788596
+         103.328766844466
+        272.2080256649731
+        31.30758738834813
+        88.25067979307288
+        272.3428736622202
+       -8.173440289984983
+        31.68694938832486
+        103.1772635880141
+        276.7936683464656
+ 4.18e+10    
+        284.3685157719326
+        103.8282419332949
+        273.0265396588832
+        31.27826027969362
+        88.57137231262958
+        273.1620876324163
+       -8.443205748054522
+        31.65911019374576
+        103.6773536078686
+         277.707148050281
+ 4.19e+10    
+        285.2931149316146
+        104.3291336938389
+         273.847117490781
+        31.24778616033305
+         88.8924967876281
+        273.9833714347334
+       -8.714724592417507
+        31.63012812940759
+        104.1788683460729
+        278.6235321398188
+ 4.2e+10     
+        286.2206145731562
+        104.8314397366293
+          274.66976131795
+        31.21616061467342
+        89.21405098550993
+        274.8067272471807
+       -8.987996433164218
+        31.59999877453237
+        104.6818054285116
+         279.542825804655
+ 4.21e+10    
+        287.1510198537555
+        105.3351575632632
+        275.4944732329491
+        31.18337918722305
+        89.53603264773122
+        275.6321571802429
+       -9.263020879170671
+        31.56871766889202
+        105.1861623720021
+        280.4650340771518
+ 4.22e+10    
+        288.0843357733957
+        105.8402845666442
+        276.3212552645002
+        31.14943738307359
+        89.85843949040473
+         276.459663277785
+       -9.539797537932017
+        31.53628031329031
+        105.6919365845392
+        281.3901618333241
+ 4.23e+10    
+        289.0205671757079
+         106.346818031235
+        277.1501093783729
+        31.11433066839605
+        90.18126920494369
+        277.2892475179718
+         -9.8183260153818
+        31.50268217005631
+        106.1991253655569
+        282.3182137937393
+ 4.24e+10    
+        289.9597187488623
+        106.8547551333257
+        277.9810374782689
+        31.07805447094863
+        90.50451945870687
+        278.1209118141762
+       -10.09860591569666
+        31.46791866355226
+        106.7077259062014
+        283.2491945244346
+ 4.25e+10    
+        290.9017950264669
+        107.3640929413152
+        278.8140414067088
+        31.04060418059718
+        90.82818789564459
+        278.9546580158952
+        -10.3806368410877
+         31.4319851806913
+        107.2177352896193
+        284.1831084378533
+ 4.26e+10    
+        291.8468003885029
+         107.874828416005
+        279.6491229459123
+        31.00197514984677
+        91.15227213694484
+        279.7904879096583
+        -10.6644183915777
+        31.39487707146832
+        107.7291504912578
+         285.119959793805
+ 4.27e+10    
+        292.7947390622725
+        108.3869584109084
+        280.4862838186796
+        30.96216269438668
+         91.4767697816812
+        280.6284032199383
+       -10.94995016476413
+        31.35658964950249
+        108.2419683791799
+        286.0597527004481
+ 4.28e+10    
+          293.74561512337
+         108.900479672571
+        281.3255256892732
+        30.92116209364632
+        91.80167840746057
+        281.4684056100635
+       -11.23723175556908
+        31.31711819259055
+        108.7561857143916
+        287.0024911152846
+ 4.29e+10    
+        294.6994324966741
+        109.4153888409074
+        282.1668501642944
+        30.87896859136244
+        92.12699557107153
+        282.3104966831251
+       -11.52626275597497
+         31.2764579432733
+        109.2717991511848
+        287.9481788461893
+ 4.3e+10     
+         295.656194957362
+        109.9316824495478
+        283.0102587935654
+        30.83557739615894
+        92.45271880913548
+        283.1546779828866
+       -11.81704275474698
+        31.23460410941176
+        109.7888052374904
+        288.8968195524452
+ 4.31e+10    
+        296.6159061319416
+        110.4493569262013
+        283.8557530709985
+         30.7909836821375
+        92.77884563875463
+        284.0009509946906
+       -12.10957133714174
+        31.19155186477499
+        110.3072004152475
+        289.8484167458085
+ 4.32e+10    
+        297.5785694993084
+        110.9684085930312
+        284.7033344354803
+        30.74518258947882
+        93.10537355816358
+        284.8493171463634
+       -12.40384808460295
+         31.1472963496397
+        110.8269810207845
+         290.802973791588
+ 4.33e+10    
+        298.5441883918157
+        111.4888336670427
+        285.5530042717353
+        30.69816922505612
+        93.43230004738025
+        285.6997778091234
+       -12.69987257444312
+        31.10183267139955
+        111.3481432852138
+        291.7604939097459
+ 4.34e+10    
+        299.5127659963723
+         112.010628260485
+        286.4047639112049
+        30.64993866305825
+        93.75962256885721
+         286.552334298485
+       -12.99764437951282
+        31.05515590518617
+        111.8706833348393
+        292.7209801760175
+ 4.35e+10    
+        300.4843053555537
+        112.5337883812657
+        287.2586146329115
+        30.60048594562454
+        94.08733856813295
+        287.4069878751567
+       -13.29716306785601
+        31.00726109449991
+        112.3945971915781
+        293.6844355230525
+ 4.36e+10    
+        301.4588093687383
+        113.0583099333806
+        288.1145576643348
+        30.54980608348992
+        94.41544547448497
+        288.2637397459483
+       -13.59842820235272
+        30.95814325185223
+        112.9198807733942
+        294.6508627415709
+ 4.37e+10    
+        302.4362807932561
+        113.5841887173528
+        288.9725941822694
+        30.49789405664016
+        94.74394070158083
+        289.1225910646673
+       -13.90143934034868
+        30.90779735941668
+        113.4465298947456
+        295.6202644815385
+ 4.38e+10    
+        303.4167222455648
+        114.1114204306889
+        289.8327253136985
+        30.44474481497838
+        95.07282164813215
+        289.9835429330193
+       -14.20619603327204
+        30.85621836969175
+        113.9745402670453
+        296.5926432533658
+ 4.39e+10    
+        304.4001362024359
+        114.6400006683451
+        290.6949521366501
+        30.39035327900003
+        95.40208569854597
+        290.8465964015047
+       -14.51269782623734
+        30.80340120617257
+        114.5039074991337
+        297.5680014291189
+ 4.4e+10     
+        305.3865250021697
+        115.1699249232092
+        291.5592756810652
+        30.33471434047997
+        95.73173022357916
+        291.7117524703157
+       -14.82094425763669
+        30.74934076403277
+        115.0346270977658
+         298.546341243749
+ 4.41e+10    
+        306.3758908458191
+        115.7011885865924
+         292.425696929652
+         30.2778228631674
+        96.06175258098955
+        292.5790120902271
+       -15.13093485871824
+        30.69403191081645
+        115.5666944681102
+         299.527664796349
+ 4.42e+10    
+        307.3682357984357
+        116.2337869487376
+        293.2942168187478
+        30.21967368349222
+        96.39215011619105
+        293.4483761634955
+       -15.44266915315264
+        30.63746948713878
+        116.1001049142615
+        300.5119740514119
+ 4.43e+10    
+        308.3635617903397
+        116.7677151993384
+         294.164836239175
+        30.16026161127975
+        96.72292016290531
+        294.3198455447429
+       -15.75614665658631
+        30.57964830739736
+        116.6348536397648
+         301.499270840121
+ 4.44e+10    
+        309.3618706183941
+        117.3029684280705
+        295.0375560370916
+        30.09958143047513
+          97.054060043815
+        295.1934210418507
+       -16.07136687618327
+        30.52056316049141
+        117.1709357481549
+        302.4895568616502
+ 4.45e+10    
+        310.3631639473138
+        117.8395416251383
+        295.9123770148486
+        30.03762789987776
+        97.38556707121735
+        296.0691034168469
+       -16.38832931015383
+          30.460208810551
+        117.7083462435065
+        303.4828336844836
+ 4.46e+10    
+        311.3674433109774
+        118.3774296818335
+        296.7892999318385
+         29.9743957538838
+        97.71743854767668
+        296.9468933867921
+       -16.70703344727207
+        30.39857999767523
+        118.2470800309978
+        304.4791027477518
+ 4.47e+10    
+        312.3747101137631
+        118.9166273911049
+        297.6683255053426
+        29.90987970323802
+        98.04967176667674
+        297.8267916246609
+       -17.02747876638056
+        30.33567143867864
+        118.7871319174876
+        305.4783653625827
+ 4.48e+10    
+        313.3849656319102
+        119.4571294481446
+        298.5494544113807
+        29.84407443579508
+        98.38226401327465
+          298.70879876023
+       -17.34966473588389
+        30.27147782784688
+        119.3284966121039
+        306.4806227134723
+ 4.49e+10    
+        314.3982110148737
+        119.9989304509823
+        299.4326872855534
+        29.77697461728858
+        98.71521256475161
+        299.5929153809535
+       -17.67359081322959
+        30.20599383770087
+        119.8711687268476
+        307.4858758596739
+ 4.5e+10     
+        315.4144472867251
+        120.5420249010975
+        300.3180247238852
+        29.70857489210883
+        99.04851469126596
+        300.4791420328426
+       -17.99925644437807
+        30.13921411976907
+        120.4151427772048
+        308.4941257365928
+ 4.51e+10    
+        316.4336753475482
+        121.0864072040399
+        301.2054672836673
+        29.63886988409024
+         99.3821676565055
+        301.3674792213464
+       -18.32666106326072
+        30.07113330536828
+        120.9604131827775
+        309.5053731572146
+ 4.52e+10    
+         317.455895974861
+        121.6320716700668
+        302.0950154842932
+         29.5678541973047
+          99.716168718338
+         302.257927412224
+       -18.65580409122641
+        30.00174600639226
+        121.5069742679205
+        310.5196188135271
+ 4.53e+10    
+         318.481109825057
+        122.1790125147891
+         302.986669808099
+        29.49552241686528
+        100.0505151294633
+        303.1504870324171
+       -18.98668493647684
+        29.93104681610885
+        122.0548202623975
+         311.536863277982
+ 4.54e+10    
+        319.5093174348496
+        122.7272238598339
+        303.8804307011952
+         29.4218691097365
+        100.3852041380633
+        304.0451584709214
+       -19.31930299349047
+        29.85903030996425
+        122.6039453020442
+        312.5571070049526
+ 4.55e+10    
+        320.5405192227492
+        123.2766997335172
+         304.776298574303
+        29.34688882555305
+        100.7202329884538
+        304.9419420796577
+       -19.65365764243571
+        29.78569104639568
+        123.1543434294485
+        313.5803503322174
+ 4.56e+10    
+        321.5747154905433
+        123.8274340715298
+        305.6742738035801
+        29.27057609744574
+        101.0555989217331
+        305.8408381743387
+        -19.9897482485724
+        29.71102356765083
+        123.7060085946399
+        314.6065934824566
+ 4.57e+10    
+        322.6119064247995
+        124.3794207176376
+        306.5743567314531
+        29.19292544287554
+         101.391299176432
+        306.7418470353318
+       -20.32757416164319
+        29.63502240061534
+        124.2589346557947
+        315.6358365647631
+ 4.58e+10    
+        323.6520920983833
+        124.9326534243913
+        307.4765476674455
+        29.11393136447456
+        101.7273309891636
+         307.644968908525
+       -20.66713471525355
+        29.55768205764746
+        124.8131153799492
+        316.6680795761679
+ 4.59e+10    
+        324.6952724719854
+         125.487125853853
+        308.3808468889981
+        29.03358835089447
+         102.063691595271
+        308.5502040061888
+       -21.00842922624151
+        29.47899703741921
+         125.368544443732
+        317.7033224031796
+ 4.6e+10     
+        325.7414473956748
+        126.0428315783311
+        309.2872546422955
+        28.95189087766159
+        102.4003782294759
+        309.4575525078333
+       -21.35145699403666
+        29.39896182576562
+        125.9252154341029
+        318.7415648233466
+ 4.61e+10    
+         326.790616610458
+        126.5997640811318
+        310.1957711430852
+         28.8688334080398
+        102.7373881265256
+        310.3670145610675
+       -21.69621730000897
+        29.31757089653952
+        126.4831218491069
+        319.7828065068175
+ 4.62e+10    
+        327.8427797498564
+        127.1579167573195
+        311.1063965774939
+        28.78441039389932
+        103.0747185218396
+         311.278590282452
+       -22.04270940680692
+        29.23481871247376
+        127.0422570986409
+        320.8270470179303
+ 4.63e+10    
+        328.8979363415019
+        127.7172829144933
+        312.0191311028514
+        28.69861627659297
+         103.412366652157
+        312.1922797583558
+       -22.39093255768611
+        29.15069972605077
+        127.6026145052336
+        321.8742858168158
+ 4.64e+10    
+        329.9560858087402
+        128.2778557735738
+        312.9339748484952
+        28.61144548783798
+        103.7503297561804
+        313.1080830458031
+       -22.74088597582724
+        29.06520838037606
+        128.1641873048342
+        322.9245222609994
+ 4.65e+10    
+        331.0172274722551
+         128.839628469603
+        313.8509279165927
+        28.52289245060527
+        104.0886050752225
+        314.0260001733283
+       -23.09256886364471
+        28.97833911006114
+        128.7269686476193
+        323.9777556070365
+ 4.66e+10    
+        332.0813605517047
+        129.4025940525576
+        314.7699903829451
+        28.43295158001418
+        104.4271898538487
+         314.946031141816
+       -23.44598040208514
+        28.89008634210976
+        129.2909515988069
+        325.0339850121487
+ 4.67e+10    
+         333.148484167371
+        129.9667454881731
+        315.6911622977981
+        28.34161728423351
+        104.7660813405214
+        315.8681759253542
+       -23.80111974991664
+        28.80044449681182
+        129.8561291394867
+        326.0932095358761
+ 4.68e+10    
+        334.2185973418264
+        130.5320756587841
+        316.6144436866516
+        28.24888396538849
+        105.1052767882424
+        316.7924344720686
+       -24.15798604300788
+        28.70940798864299
+        130.4224941674604
+        327.1554281417477
+ 4.69e+10    
+        335.2916990016088
+        131.0985773641714
+        317.5398345510589
+        28.15474602047371
+        105.4447734551952
+        317.7188067049709
+       -24.51657839359891
+        28.61697122716908
+        130.9900394980967
+        328.2206396989621
+ 4.7e+10     
+        336.3677879789195
+        131.6662433224276
+        318.4673348694329
+        28.05919784227171
+        105.7845686053853
+        318.6472925227947
+       -24.87689588956179
+        28.52312861795678
+        131.5587578651959
+        329.2888429840751
+ 4.71e+10    
+        337.4468630133262
+        132.2350661708313
+        319.3969445978465
+         27.9622338202761
+        106.1246595092808
+        319.5778918008297
+       -25.23893759365291
+        28.42787456348954
+        132.1286419218692
+        330.3600366827135
+ 4.72e+10    
+        338.5289227534832
+        132.8050384667354
+        320.3286636708306
+        27.86384834162218
+        106.4650434444522
+        320.5106043917639
+       -25.60270254275591
+        28.33120346408883
+        132.6996842414309
+        331.4342193912899
+ 4.73e+10    
+        339.6139657588661
+        133.3761526884684
+        321.2624920021719
+        27.76403579202029
+        106.8057176962106
+        321.4454301265073
+       -25.96818974711604
+        28.23310971884057
+        133.2718773182999
+        332.5113896187368
+ 4.74e+10    
+        340.7019905015192
+        133.9484012362455
+        322.1984294857059
+        27.66279055669614
+        107.1466795582446
+        322.3823688150302
+       -26.33539818956594
+        28.13358772652622
+        133.8452135689171
+        333.5915457882521
+ 4.75e+10    
+        341.7929953678135
+        134.5217764330968
+         323.136475996112
+        27.56010702133505
+        107.4879263332582
+        323.3214202471876
+       -26.70432682474291
+          28.032631886559
+        134.4196853326728
+        334.6746862390517
+ 4.76e+10    
+        342.8869786602222
+        135.0962705258035
+         324.076631389706
+        27.45597957303155
+        107.8294553336063
+          324.26258419355
+       -27.07497457829815
+        27.93023659992463
+        134.9952848728479
+        335.7608092281458
+ 4.77e+10    
+        343.9839385991045
+        135.6718756858488
+        325.0188955052225
+        27.35040260124293
+        108.1712638819283
+        325.2058604062208
+       -27.44734034609717
+        27.82639627012698
+        135.5720043775668
+        336.8499129321153
+ 4.78e+10    
+         345.083873324506
+        136.2485840103819
+        325.9632681646126
+        27.24337049874795
+        108.5133493117836
+        326.1512486196694
+       -27.82142299341294
+        27.72110530413775
+        136.1498359607627
+        337.9419954489086
+ 4.79e+10    
+        346.1867808979718
+        136.8263875231921
+        326.9097491738181
+        27.13487766261003
+        108.8557089682826
+        327.0987485515417
+       -28.19722135411075
+        27.61435811335048
+        136.7287716631555
+        339.0370547996454
+ 4.8e+10     
+        347.2926593043677
+        137.4052781756985
+        327.8583383235668
+        27.02491849514382
+        109.1983402087203
+         328.048359903487
+       -28.57473422982578
+        27.50614911453888
+        137.3088034532422
+        340.1350889304348
+ 4.81e+10    
+        348.4015064537188
+        137.9852478479489
+        328.8090353901438
+        26.91348740488632
+        109.5412404032054
+        329.0000823619691
+       -28.95396038913264
+        27.39647273081917
+        137.8899232282987
+        341.2360957142072
+ 4.82e+10    
+        349.5133201830577
+        138.5662883496338
+        329.7618401361786
+        26.80057880757238
+         109.884406935291
+        329.9539155990866
+       -29.33489856670811
+        27.28532339261586
+        138.4721228153956
+        342.3400729525507
+ 4.83e+10    
+        350.6280982582867
+        139.1483914211116
+        330.7167523114214
+        26.68618712711305
+        110.2278372026022
+         330.909859273378
+       -29.71754746248607
+         27.1726955386319
+         139.055393972425
+        343.4470183775674
+ 4.84e+10    
+        351.7458383760501
+        139.7315487344463
+        331.6737716535192
+        26.57030679657843
+        110.5715286174643
+        331.8679130306434
+       -30.10190574080625
+        27.05858361682174
+        139.6397283891399
+        344.5569296537336
+ 4.85e+10    
+        352.8665381656188
+        140.3157518944581
+        332.6328978887902
+        26.45293225918343
+        110.9154786075287
+        332.8280765047438
+       -30.48797202955517
+        26.94298208536827
+         140.225117688206
+        345.6698043797775
+ 4.86e+10    
+        353.9901951907893
+        140.9009924397851
+        333.5941307329975
+        26.33405796927718
+        111.2596846163976
+        333.7903493184141
+       -30.87574491930133
+        26.82588541366267
+        140.8115534262668
+        346.7856400905641
+ 4.87e+10    
+        355.1168069517924
+        141.4872618439611
+        334.5574698921217
+        26.21367839333552
+        111.6041441042492
+        334.7547310840661
+       -31.26522296242297
+        26.70728808328808
+        141.3990270950189
+        347.9044342589918
+ 4.88e+10    
+        356.2463708872089
+        142.0745515164995
+        335.5229150631289
+        26.09178801095658
+        111.9488545484588
+        335.7212214045925
+       -31.65640467223049
+        26.58718458900523
+        141.9875301223013
+        349.0261842978996
+ 4.89e+10    
+         357.378884375908
+        142.6628528039964
+        336.4904659347384
+        25.96838131585957
+        112.2938134442216
+         336.689819874169
+       -32.04928852208165
+        26.46556943974188
+        142.5770538731966
+         350.150887561987
+ 4.9e+10     
+        358.5143447389872
+        143.2521569912424
+        337.4601221881927
+        25.84345281688554
+        112.6390183051719
+        337.6605260790545
+       -32.44387294449184
+        26.34243715958461
+        143.1675896511452
+        351.2785413497421
+ 4.91e+10    
+        359.6527492417259
+         143.842455302346
+        338.4318834980166
+        25.71699703900213
+        112.9844666640035
+        338.6333395983879
+       -32.84015633023763
+        26.21778228877292
+        143.7591286990692
+        352.4091429053809
+ 4.92e+10    
+        360.7940950955518
+        144.4337389018726
+        339.4057495327866
+        25.58900852430902
+        113.3301560730861
+        339.6082600049841
+       -33.23813702745542
+        26.09159938469643
+        144.3516622005118
+        353.5426894207989
+ 4.93e+10    
+        361.9383794600177
+        145.0259988959933
+        340.3817199558849
+        25.45948183304763
+        113.6760841050824
+        340.5852868661307
+       -33.63781334073417
+        25.96388302289357
+        144.9451812807876
+        354.6791780375277
+ 4.94e+10    
+          363.08559944479
+        145.6192263336472
+        341.3597944262696
+        25.32841154461142
+        114.0222483535628
+        341.5644197443779
+       -34.03918353020322
+         25.8346277980533
+         145.539677008145
+         355.818605848713
+ 4.95e+10    
+        364.2357521116423
+        146.2134122077154
+        342.3399725992239
+        25.19579225855954
+        114.3686464336204
+        342.5456581983327
+       -34.44224581061474
+        25.70382832501756
+        146.1351403949394
+        356.9609699010825
+ 4.96e+10    
+         365.388834476472
+        146.8085474562094
+        343.3222541271195
+        25.06161859563136
+        114.7152759824819
+        343.5290017834456
+       -34.84699835042155
+        25.57147923978774
+        146.7315623988241
+        358.1062671969502
+ 4.97e+10    
+        366.5448435113112
+        147.4046229634675
+        344.3066386601657
+        24.92588519876327
+         115.062134660119
+        344.5144500527965
+       -35.25343927085022
+        25.43757520053003
+         147.328933923945
+        359.2544946962054
+ 4.98e+10    
+        367.7037761463621
+        148.0016295613698
+         345.293125847174
+        24.78858673410742
+        115.4092201498598
+        345.5020025578867
+       -35.66156664496955
+        25.30211088858514
+        147.9272458221559
+        360.4056493183305
+ 4.99e+10    
+        368.8656292720356
+        148.5995580305592
+         346.281715336298
+        24.64971789205119
+        115.7565301589944
+        346.4916588494171
+       -36.07137849675475
+        25.16508100947766
+        148.5264888942413
+        361.5597279444164
+ 5e+10       
+        370.0303997410026
+        149.1983991016791
+        347.2724067757939
+        24.50927338823869
+        116.1040624193835
+        347.4834184780744
+         -36.482872800148
+        25.02648029392691
+          149.12665389115
+        362.7167274191886
+ 5.01e+10    
+          371.19808437025
+        149.7981434566223
+        348.2651998147702
+        24.36724796459299
+        116.4518146880638
+          348.47728099531
+        -36.8960474781142
+        24.88630349886047
+        149.7277315152488
+         363.876644553057
+ 5.02e+10    
+        372.3686799431603
+        150.3987817297911
+        349.2600941039277
+        24.22363639034011
+        116.7997847478511
+        349.4732459541212
+       -37.31090040169385
+         24.7445454084263
+         150.329712421577
+        365.0394761241485
+ 5.03e+10    
+        373.5421832115824
+        151.0003045093714
+        350.2570892963179
+        24.07843346303271
+        117.1479704079434
+        350.4713129098283
+        -37.7274293890521
+        24.60120083500803
+        150.9325872191239
+        366.2052188803756
+ 5.04e+10    
+        374.7185908979278
+        151.6027023386182
+         351.256185048083
+        23.93163400957587
+        117.4963695045217
+        351.4714814208496
+       -38.14563220452435
+        24.45626462023964
+        151.5363464721113
+        367.3738695414975
+ 5.05e+10    
+        375.8978996972685
+        152.2059657171529
+        352.2573810191973
+         23.7832328872529
+        117.8449799013489
+        352.4737510494784
+       -38.56550655765914
+        24.30973163602098
+        152.1409807012905
+        368.5454248011948
+ 5.06e+10    
+        377.0801062794477
+         152.810085102275
+        353.2606768742207
+        23.63322498475148
+         118.193799490369
+        353.4781213626562
+        -38.9870501022578
+        24.16159678553439
+        152.7464803852543
+        369.7198813291558
+ 5.07e+10    
+         378.265207291196
+        153.4150509102837
+        354.2660722830311
+        23.48160522319041
+        118.5428261923022
+        354.4845919327423
+        -39.4102604354115
+        24.01185500426079
+        153.3528359617553
+        370.8972357731668
+ 5.08e+10    
+        379.4531993582642
+        154.0208535178124
+        355.2735669215703
+        23.32836855714691
+        118.8920579572406
+        355.4931623382881
+       -39.83513509653594
+        23.86050126099678
+        153.9600378290422
+        372.0774847612163
+ 5.09e+10    
+        380.6440790875574
+         154.627483263178
+        356.2831604725812
+        23.17350997568319
+          119.24149276524
+        356.5038321648009
+        -40.2616715664037
+        23.70753055887065
+        154.5680763472044
+        373.2606249035995
+ 5.1e+10     
+        381.8378430692834
+         155.234930447738
+        357.2948526263512
+        23.01702450337339
+        119.5911286269136
+        357.5166010055171
+       -40.68986726617484
+        23.55293793635989
+        155.1769418395306
+        374.4466527950439
+ 5.11e+10    
+         383.034487879109
+        155.8431853372639
+        358.3086430814433
+        22.85890720133079
+        119.9409635840197
+        358.5314684621634
+       -41.11971955642468
+        23.39671846830699
+        155.7866245938786
+        375.6355650168304
+ 5.12e+10    
+        384.2340100803237
+        156.4522381633246
+        359.3245315454365
+        22.69915316823385
+        120.2909957100516
+        359.5484341457267
+       -41.55122573617139
+        23.23886726693587
+        156.3971148640591
+        376.8273581389323
+ 5.13e+10    
+        385.4364062260143
+        157.0620791246831
+        360.3425177356629
+         22.5377575413521
+        120.6412231108242
+        360.5674976772131
+       -41.98438304190091
+        23.07937948286752
+        157.0084028712291
+        378.0220287221551
+ 5.14e+10    
+        386.6416728612495
+        157.6726983887053
+        361.3626013799353
+        22.37471549757171
+        120.9916439250571
+        361.5886586884128
+       -42.41918864659151
+        22.91825030613432
+        157.6204788052988
+        379.2195733202912
+ 5.15e+10    
+        387.8498065252685
+        158.2840860927798
+         362.384782217288
+        22.21002225441983
+        121.3422563249609
+        362.6119168226626
+       -42.85563965873711
+        22.75547496719522
+         158.233332826351
+        380.4199884822785
+ 5.16e+10    
+          389.06080375368
+        158.8962323457522
+        363.4090599987037
+        22.04367307108789
+        121.6930585168152
+        363.6372717356002
+        -43.2937331213695
+        22.59104873794804
+        158.8469550660721
+        381.6232707543643
+ 5.17e+10    
+        390.2746610806749
+        159.5091272293702
+        364.4354344878487
+         21.8756632494552
+        122.0440487415522
+        364.6647230959288
+        -43.7334660110807
+        22.42496693274215
+         159.461335629194
+        382.8294166822863
+ 5.18e+10    
+        391.4913750412395
+        160.1227607997408
+        365.4639054618018
+        21.70598813510911
+        122.3952252753316
+         365.694270586171
+        -44.1748352370445
+        22.25722490938968
+        160.0764645949515
+         384.038422813451
+ 5.19e+10    
+        392.7109421733844
+        160.7371230888004
+        366.4944727117817
+        21.53464311836607
+        122.7465864301185
+        366.7259139034272
+        -44.6178376400382
+        22.08781807017461
+        160.6923320185481
+        385.2502856991277
+ 5.2e+10     
+        393.9333590203719
+        161.3522041057965
+        367.5271360438794
+        21.36162363528987
+        123.0981305542576
+        367.7596527601277
+       -45.06246999146413
+        21.91674186286195
+        161.3089279326358
+        386.4650018966426
+ 5.21e+10    
+        395.1586221329649
+        161.9679938387824
+        368.5618952797834
+        21.18692516870848
+        123.4498560330455
+        368.7954868847889
+       -45.50872899237213
+        21.74399178170346
+        161.9262423488067
+        387.6825679715889
+ 5.22e+10    
+        396.3867280716691
+         162.584482256123
+         369.598750257508
+        21.01054324922993
+        123.8017612893026
+        369.8334160227685
+       -45.95661127248218
+        21.56956336844344
+        162.5442652590974
+        388.9029805000363
+ 5.23e+10    
+        397.6176734089988
+        163.2016593080138
+        370.6377008321177
+        20.83247345625534
+        124.1538447839408
+        370.8734399370122
+       -46.40611338920805
+        21.39345221332083
+        163.1629866375028
+        390.1262360707518
+ 5.24e+10    
+        398.8514547317336
+        163.8195149280107
+        371.6787468764548
+        20.65271141899047
+        124.5061050165315
+        371.9155584088063
+       -46.85723182668147
+        21.21565395607163
+        163.7823964415059
+        391.3523312874302
+ 5.25e+10    
+        400.0880686431977
+         164.438039034575
+        372.7218882818633
+         20.4712528174555
+        124.8585405258714
+        372.9597712385307
+       -47.30996299477903
+        21.03616428692681
+         164.402484613616
+        392.5812627709262
+ 5.26e+10    
+        401.3275117655384
+        165.0572215326254
+        373.7671249589114
+        20.28809338349082
+         125.211149890544
+        374.0060782464036
+       -47.76430322814867
+        20.85497894760925
+        165.0232410829215
+        393.8130271614934
+ 5.27e+10    
+        402.5697807420158
+        165.6770523151082
+        374.8144568381151
+        20.10322890176349
+        125.5639317294837
+        375.0544792732318
+       -48.22024878523939
+        20.67209373232853
+        165.6446557666531
+        395.0476211210383
+ 5.28e+10    
+        403.8148722392954
+        166.2975212645736
+        375.8638838706622
+        19.91665521076769
+        125.9168847025329
+         376.104974181157
+       -48.67779584733253
+         20.4875044887723
+        166.2667185717607
+        396.2850413353744
+ 5.29e+10    
+        405.0627829497552
+        166.9186182547699
+        376.9154060291351
+        19.72836820382539
+         126.270007511002
+        377.1575628544012
+       -49.13694051757466
+        20.30120711909557
+        166.8894193964992
+        397.5252845164803
+ 5.3e+10     
+        406.3135095937967
+        167.5403331522448
+        377.9690233082286
+        19.53836383008233
+        126.6232988982231
+        378.2122452000127
+       -49.59767882001414
+        20.11319758090708
+        167.5127481320304
+        398.7683474047732
+ 5.31e+10    
+        407.5670489221558
+        168.1626558179612
+          379.02473572547
+        19.34663809550132
+        126.9767576501039
+        379.2690211486089
+       -50.06000669863929
+        19.92347188825279
+        168.1366946640337
+        400.0142267713837
+ 5.32e+10    
+        408.8233977182394
+         168.785576108927
+        380.0825433219464
+        19.15318706385435
+        127.3303825956819
+        380.3278906551245
+       -50.52392001642008
+        19.73202611259618
+        168.7612488743304
+        401.2629194204345
+ 5.33e+10    
+        410.0825528004461
+        169.4090838798317
+        381.1424461630167
+        18.95800685770844
+        127.6841726076704
+        381.3888536995489
+       -50.98941455435263
+        19.53885638379572
+        169.3864006425189
+        402.5144221913355
+ 5.34e+10    
+        411.3445110245128
+        170.0331689846993
+        382.2044443390318
+        18.76109365941065
+        128.0381266030091
+        382.4519102876699
+       -51.45648601050739
+        19.34395889107851
+        170.0121398476224
+        403.7687319610703
+ 5.35e+10    
+        412.6092692858581
+        170.6578212785528
+        383.2685379660575
+        18.56244371206813
+        128.3922435434073
+        383.5170604518141
+       -51.92512999908107
+          19.147329884011
+        170.6384563697485
+        405.0258456465036
+ 5.36e+10    
+        413.8768245219325
+        171.2830306190893
+        384.3347271865907
+        18.36205332052572
+        128.7465224358903
+        384.5843042515909
+       -52.39534204945203
+        18.94896567346583
+        171.2653400917618
+        406.2857602066893
+ 5.37e+10    
+        415.1471737145847
+        171.9087868683671
+        385.4030121702713
+        18.15991885233914
+        129.1009623333382
+        385.6536417746279
+       -52.86711760524003
+        18.74886263258509
+        171.8927809009647
+        407.5484726451763
+ 5.38e+10    
+        416.4203138924191
+        172.5350798945069
+        386.4733931146104
+        17.95603673874411
+        129.4555623350272
+        386.7250731373151
+       -53.34045202337049
+        18.54701719773994
+        172.5207686907958
+        408.8139800123387
+ 5.39e+10    
+        417.6962421331769
+        173.1618995734014
+        387.5458702456968
+        17.75040347562206
+        129.8103215871654
+        387.7985984855358
+       -53.81534057314325
+        18.34342586948571
+        173.1492933625339
+        410.0822794076925
+ 5.4e+10     
+        418.9749555661094
+        173.7892357904403
+        388.6204438189203
+        17.54301562446167
+         130.165239283429
+        388.8742179954118
+       -54.29177843530595
+        18.13808521351365
+        173.7783448270195
+        411.3533679822334
+ 5.41e+10    
+        420.2564513743654
+        174.4170784422466
+        389.6971141196856
+        17.33386981331606
+        130.5203146654952
+        389.9519318740394
+       -54.76976070113269
+        17.93099186159841
+        174.4079130063843
+        412.6272429407682
+ 5.42e+10    
+        421.5407267973854
+        175.0454174384214
+        390.7758814641276
+         17.1229627377552
+        130.8755470235724
+        391.0317403602223
+       -55.24928237150834
+         17.7221425125402
+        175.0379878357936
+         413.903901544263
+ 5.43e+10    
+        422.8277791332947
+         175.674242703306
+        391.8567461998284
+        16.91029116181461
+        131.2309356969293
+        392.1136437252117
+       -55.73033835601767
+        17.51153393310435
+        175.6685592652016
+         415.183341112191
+ 5.44e+10    
+        424.1176057413143
+        176.3035441777514
+          392.93970870653
+        16.69585191893895
+        131.5864800744214
+        393.1976422734404
+       -56.21292347204118
+        17.29916295895413
+         176.299617261117
+        416.4655590248848
+ 5.45e+10    
+        425.4102040441655
+        176.9333118209018
+        394.0247693968545
+        16.47964191292104
+        131.9421795950152
+        394.2837363432589
+       -56.69703244385605
+        17.08502649558102
+        176.9311518083808
+         417.750552725897
+ 5.46e+10    
+        426.7055715304897
+        177.5635356119899
+        395.1119287170148
+         16.2616581188362
+        132.2980337483102
+        395.3719263076686
+        -57.1826599017442
+        16.86912151922853
+        177.5631529119569
+        419.0383197243672
+ 5.47e+10    
+        428.0037057572703
+         178.194205552144
+        396.2011871475289
+        16.04189758397093
+        132.6540420750582
+        396.4622125750588
+       -57.66980038110653
+        16.65144507781205
+        178.1956105987319
+        420.3288575973918
+ 5.48e+10    
+        429.3046043522601
+        178.8253116662042
+        397.2925452039379
+        15.82035742874765
+         133.010204167682
+         397.554595589938
+       -58.15844832158376
+        16.43199429183338
+        178.8285149193304
+        421.6221639923985
+ 5.49e+10    
+        430.6082650164163
+        179.4568440045566
+         398.386003437521
+        15.59703484764306
+        133.3665196707895
+        398.6490758336699
+       -58.64859806618462
+        16.21076635528976
+        179.4618559499374
+        422.9182366295302
+ 5.5e+10     
+        431.9146855263381
+        180.0887926449705
+        399.4815624360015
+        15.37192711010211
+        133.7229882816872
+        399.7456538252055
+       -59.14024386042119
+        15.98775853657851
+        180.0956237941377
+        424.2170733040313
+ 5.51e+10    
+        433.2238637367178
+        180.7211476944576
+        400.5792228242735
+        15.14503156144568
+        134.0796097508905
+        400.8443301218144
+       -59.63337985145161
+         15.7629681793953
+        180.7298085847606
+         425.518671888637
+ 5.52e+10    
+        434.5357975827852
+        181.3538992911335
+        401.6789852651071
+        14.91634562377344
+        134.4363838826326
+         401.945105319821
+       -60.12800008723091
+        15.53639270362745
+        181.3644004857427
+         426.823030335973
+ 5.53e+10    
+        435.8504850827663
+        181.9870376060967
+         402.780850459865
+        14.68586679686058
+        134.7933105353698
+        403.0479800553354
+       -60.62409851566915
+        15.30802960624154
+        181.9993896939981
+        428.1301466809538
+ 5.54e+10    
+        437.1679243403472
+        182.6205528453164
+        403.8848191492178
+        14.45359265904883
+        135.1503896222853
+        404.1529550049817
+       -61.12166898379831
+        15.07787646216546
+        182.6347664413011
+         429.440019043194
+ 5.55e+10    
+        438.4881135471403
+        183.2544352515349
+         404.990892113858
+        14.21952086813187
+        135.5076211117912
+        405.2600308866379
+       -61.62070523694781
+        14.84593092516384
+        183.2705209961811
+        430.7526456294138
+ 5.56e+10    
+        439.8110509851551
+        183.8886751061774
+        406.0990701752131
+        13.98364916223412
+        135.8650050280259
+         406.369208460159
+       -62.12120091792787
+        14.61219072870885
+        183.9066436658285
+        432.0680247358619
+ 5.57e+10    
+        441.1367350292761
+         184.523262731279
+        407.2093541961616
+        13.74597536068393
+        136.2225414513523
+        407.4804885281158
+       -62.62314956622298
+        14.37665368684356
+        184.5431247980137
+        433.3861547507294
+ 5.58e+10    
+         442.465164149751
+        185.1581884914163
+        408.3217450817434
+        13.50649736488028
+        136.5802305188498
+        408.5938719365207
+       -63.12654461719314
+        14.13931769504012
+        185.1799547830137
+        434.7070341565823
+ 5.59e+10    
+        443.7963369146701
+        185.7934427956576
+        409.4362437798822
+        13.26521315915307
+        136.9380724248081
+        409.7093595755598
+       -63.63137940128604
+        13.90018073105106
+        185.8171240555548
+        436.0306615327861
+ 5.6e+10     
+        445.1302519924661
+        186.4290160995187
+         410.552851282089
+        13.02212081161733
+        137.2960674212145
+        410.8269523803306
+       -64.13764714325752
+        13.65924085575453
+        186.4546230967645
+        437.3570355579424
+ 5.61e+10    
+        446.4669081544075
+        187.0648989069364
+        411.6715686241895
+        12.77721847502018
+        137.6542158182419
+        411.9466513315626
+       -64.64534096140304
+        13.41649621399285
+        187.0924424361336
+        438.6861550123306
+ 5.62e+10    
+        447.8063042771071
+        187.7010817722455
+        412.7923968870261
+        12.53050438758179
+        138.0125179847321
+        413.0684574563547
+       -65.15445386679794
+         13.1719450354047
+        187.7305726534931
+        440.0180187803464
+ 5.63e+10    
+          449.14843934502
+        188.3375553021755
+        413.9153371971832
+         12.2819768738291
+        138.3709743486783
+        414.1923718289069
+       -65.66497876254948
+        12.92558563525008
+        188.3690043809987
+        441.3526258529535
+ 5.64e+10    
+        450.4933124529671
+        188.9743101578532
+        415.0403907276997
+        12.03163434542285
+        138.7295853977035
+        415.3183955712464
+       -66.17690844305885
+         12.6774164152291
+        189.0077283051298
+        442.6899753301366
+ 5.65e+10    
+        451.8409228086445
+        189.6113370568191
+        416.1675586987789
+        11.77947530197758
+        139.0883516795378
+        416.4465298539636
+       -66.69023559329281
+        12.42743586429363
+        189.6467351686979
+         444.030066423353
+ 5.66e+10    
+        453.1912697351455
+        190.2486267750541
+        417.2968423785141
+        11.52549833187458
+        139.4472738024927
+        417.5767758969394
+       -67.20495278806881
+        12.17564255945167
+        190.2860157728672
+        445.3728984579977
+ 5.67e+10    
+        454.5443526734884
+        190.8861701490179
+        418.4282430835974
+        11.26970211306717
+        139.8063524359318
+        418.7091349700785
+        -67.7210524913491
+        11.92203516656468
+        190.9255609791857
+        446.7184708758662
+ 5.68e+10    
+        455.9001711851515
+        191.5239580776996
+        419.5617621800346
+        11.01208541387979
+        140.1655883107404
+        419.8436083940373
+       -68.23852705554751
+        11.66661244113802
+        191.5653617116283
+        448.0667832376215
+ 5.69e+10    
+        457.2587249545969
+        192.1619815246779
+        420.6974010838726
+        10.75264709379845
+        140.5249822197927
+        420.9801975409612
+       -68.75736872084754
+        11.40937322910404
+         192.205408958651
+        449.4178352252706
+ 5.7e+10     
+        458.6200137918191
+        192.8002315201949
+        421.8351612619036
+        10.49138610425434
+        140.8845350184142
+        422.1189038352069
+        -69.2775696145323
+         11.1503164675972
+        192.8456937752564
+        450.7716266446376
+ 5.71e+10    
+        459.9840376348852
+        193.4386991632377
+        422.9750442323927
+        10.22830148939964
+        141.2442476248439
+         423.259728754083
+       -69.79912175032703
+        10.88944118572257
+          193.48620728507
+        452.1281574278461
+ 5.72e+10    
+        461.3507965524852
+        194.0773756236347
+        424.1170515657859
+        9.963392386876016
+        141.6041210206925
+         424.402673828577
+       -70.32201702775338
+        10.62674650531531
+        194.1269406824264
+        453.4874276358022
+ 5.73e+10    
+        462.7202907464773
+        194.7162521441607
+         425.261184885438
+         9.69665802857463
+        141.9641562513987
+        425.5477406440843
+       -70.84624723149693
+         10.3622316416947
+        194.7678852344707
+        454.8494374606836
+ 5.74e+10    
+         464.092520554453
+        195.3553200426551
+        426.4074458683239
+         9.42809774138914
+        142.3243544266825
+        426.6949308411471
+       -71.37180403078661
+        10.09589590440805
+        195.4090322832657
+        456.2141872284294
+ 5.75e+10    
+        465.4674864522898
+        195.9945707141499
+        427.5558362457629
+        9.157710947959947
+         142.684716720996
+        427.8442461161812
+       -71.89867897878811
+        9.827738697968236
+        196.0503732479142
+        457.5816774012385
+ 5.76e+10    
+        466.8451890567178
+        196.6339956330064
+        428.7063578041328
+        8.885497167410819
+        143.0452443739709
+        428.9956882222106
+       -72.42686351200987
+        9.557759522582582
+          196.69189962669
+         458.951908580063
+ 5.77e+10    
+        468.2256291278886
+        197.2735863550704
+        429.8590123855944
+        8.611456016077081
+        143.4059386908642
+        430.1492589695985
+       -72.95634894972237
+        9.285957974874258
+        197.3336029991812
+        460.3248815071195
+ 5.78e+10    
+        469.6088075719458
+        197.9133345198287
+        431.0138018888092
+          8.3355872082261
+        143.7668010430005
+        431.3049602267831
+       -73.48712649339178
+        9.012333748594894
+        197.9754750284441
+        461.7005970683846
+ 5.79e+10    
+        470.9947254436019
+        198.5532318525854
+        432.1707282696628
+        8.057890556768895
+         144.127832868213
+        432.4627939210083
+       -74.01918722612703
+        8.736886635329427
+        198.6175074631673
+        463.0790562961129
+ 5.8e+10     
+        472.3833839487148
+        199.1932701666417
+        433.3297935419828
+          7.7783659739637
+        144.4890356712793
+         433.622762039058
+       -74.55252211214024
+        8.459616525192498
+        199.2596921398475
+        464.4602603713436
+ 5.81e+10    
+        473.7747844468734
+        199.8334413654928
+         434.490999778263
+        7.497013472110428
+        144.8504110243556
+        434.7848666279893
+       -75.08712199622289
+        8.180523407516251
+        199.9020209849753
+        465.8442106264192
+ 5.82e+10    
+        475.1689284539854
+        200.4737374450316
+        435.6543491103874
+         7.21383316423789
+         145.211960567411
+        435.9491097958719
+         -75.622977603235
+        7.899607371530511
+        200.5444860172341
+        467.2309085475058
+ 5.83e+10    
+        476.5658176448604
+        201.1141504957639
+        436.8198437303481
+         6.92882526478054
+        145.5736860086526
+        437.1154937125116
+       -76.16007953760933
+        7.616868607033091
+        201.1870793497065
+        468.6203557771137
+ 5.84e+10    
+        477.9654538558138
+         201.754672705037
+        437.9874858909744
+        6.641990090248434
+        145.9355891249553
+        438.2840206102003
+       -76.69841828287147
+        7.332307405052735
+        201.8297931920936
+        470.0125541166233
+ 5.85e+10    
+        479.3678390872558
+         202.395296359276
+        439.1572779066573
+        6.353328059886495
+        146.2976717622829
+        439.4546927844372
+       -77.23798420117315
+        7.045924158502494
+        202.4726198529444
+        471.4075055288135
+ 5.86e+10    
+        480.7729755062954
+        203.0360138462314
+        440.3292221540675
+        6.062839696326408
+        146.6599358361085
+        440.6275125946739
+       -77.77876753284197
+        6.757719362824837
+        203.1155517418964
+        472.8052121403967
+ 5.87e+10    
+        482.1808654493453
+        203.6768176572381
+        441.5033210728866
+        5.770525626228821
+        147.0223833318342
+        441.8024824650457
+       -78.32075839594617
+         6.46769361662766
+        203.7585813719248
+        474.2056762445499
+ 5.88e+10    
+         483.591511424723
+         204.317700389486
+        442.6795771665357
+        5.476386580916502
+        147.3850163052043
+        442.9796048851126
+       -78.86394678587524
+        6.175847622311501
+         204.401701361606
+        475.6089003034513
+ 5.89e+10    
+        485.0049161152722
+        204.9586547482994
+        443.8579930028959
+        5.180423396998931
+        147.7478368827178
+        444.1588824105931
+       -79.40832257493582
+        5.882182186687658
+        205.0449044373881
+        477.0148869508282
+ 5.9e+10     
+        486.4210823809655
+        205.5996735494266
+        445.0385712150376
+        4.882637016986955
+        148.1108472620384
+        445.3403176641049
+        -79.9538755119633
+         5.58669822158766
+        205.6881834358742
+        478.4236389944925
+ 5.91e+10    
+        487.8400132615245
+        206.2407497213425
+        446.2213145019518
+        4.583028489898863
+        148.4740497123997
+         446.523913335899
+       -80.50059522195076
+        5.289396744462557
+        206.3315313061136
+        479.8351594188928
+ 5.92e+10    
+        489.2617119790442
+        206.8818763075588
+        447.4062256292758
+        4.281598971856663
+        148.8374465750097
+        447.7096721846026
+       -81.04847120569281
+        4.990278878974571
+        206.9749411119078
+        481.2494513876603
+ 5.93e+10    
+        490.6861819406088
+        207.5230464689477
+        448.5933074300253
+        3.978349726673704
+        149.2010402634512
+        448.8975970379575
+        -81.5974928394465
+        4.689345855578154
+        207.6184060341221
+        482.6665182461635
+ 5.94e+10    
+        492.1134267409238
+        208.1642534860732
+        449.7825628053225
+         3.67328212643171
+        149.5648332640795
+        450.0876907935577
+       -82.14764937460897
+        4.386599012092386
+        208.2619193730108
+        484.0863635240598
+ 5.95e+10    
+        493.5434501649387
+         208.805490761534
+        450.9739947251272
+        3.366397652049505
+         149.928828136417
+         451.279956419593
+       -82.69892993741122
+        4.082039794264091
+         208.905474550551
+        485.5089909378562
+ 5.96e+10    
+        494.9762561904827
+        209.4467518223162
+        452.1676062289739
+        3.057697893841503
+        150.2930275135458
+        452.4743969555864
+       -83.25132352862931
+         3.77566975632077
+        209.5490651127879
+         486.934404393467
+ 5.97e+10    
+        496.4118489909004
+        210.0880303221578
+        453.3634004266918
+        2.747184552066843
+        150.6574341024963
+        453.6710155131414
+       -83.80481902331312
+        3.467490561514765
+        210.1926847321892
+         488.362607988775
+ 5.98e+10    
+        497.8502329376832
+        210.7293200439226
+        454.5613804991588
+        2.434859437468589
+        151.0220506846343
+        454.8698152766801
+       -84.35940517053092
+        3.157503982658092
+        210.8363272100106
+        489.7936060162014
+ 5.99e+10    
+         499.291412603115
+         211.370614901981
+        455.7615496990124
+        2.120724471803678
+         151.386880116042
+        456.0707995041839
+       -84.91507059313223
+        2.845711902646897
+        211.4799864786715
+        491.2274029652699
+ 6e+10       
+        500.7353927629113
+         212.011908944607
+        456.9639113514019
+        1.804781688362443
+        151.7519253279008
+        457.2739715279411
+       -85.47180378752836
+        2.532116314976342
+        212.1236566041388
+        492.6640035251748
+ 6.01e+10    
+        502.1821783988652
+        212.6531963563808
+        458.1684688547157
+        1.487033232478895
+        152.1171893268671
+        458.4793347552915
+        -86.0295931234904
+        2.216719324246501
+        212.7673317883244
+        494.1034125873578
+ 6.02e+10    
+         503.631774701498
+        213.2944714606031
+        459.3752256813237
+        1.167481362031017
+        152.4826751954479
+        459.6868926693709
+       -86.58842684396475
+         1.89952314665776
+        213.4110063714884
+        495.5456352480797
+ 6.03e+10    
+        505.0841870727036
+        213.9357287217191
+        460.5841853783083
+       0.8461284479305053
+        152.8483860923704
+        460.8966488298508
+       -87.14829306490644
+        1.580530110496905
+        214.0546748346573
+        496.9906768109987
+ 6.04e+10    
+        506.5394211284095
+        214.5769627477523
+        461.7953515682084
+       0.5229769746034556
+        153.2143252529519
+        462.1086068736934
+        -87.7091797751311
+        1.259742656613039
+        214.6983318020468
+        498.4385427897483
+ 6.05e+10    
+        507.9974827012213
+        215.2181682927475
+        463.0087279497557
+       0.1980295404607038
+        153.5804959894654
+        463.3227705158928
+       -88.27107483618505
+       0.9371633388836855
+        215.3419720434975
+        499.8892389105196
+ 6.06e+10    
+        509.4583778430949
+        215.8593402592271
+        464.2243182986158
+      -0.1287111416424125
+        153.9469016915006
+        464.5391435502243
+       -88.83396598223278
+        0.612794824670992
+        215.9855904769207
+        501.3427711146453
+ 6.07e+10    
+         510.922112827979
+        216.5004737006504
+        465.4421264681276
+      -0.4572422439559922
+        154.3135458263248
+        465.7577298499929
+       -89.39784081996414
+       0.2866398952678466
+        216.6291821707531
+        502.7991455611858
+ 6.08e+10    
+        512.3886941544948
+        217.1415638238907
+        466.6621563900492
+      -0.7875608233950189
+         154.680431939239
+        466.9785333687841
+       -89.96268682851877
+      -0.0412985536653494
+        217.2727423464213
+         504.258368629515
+ 6.09e+10    
+        513.8581285485882
+        217.7826059917154
+        467.8844120752951
+       -1.119663821110599
+        155.0475636539306
+        468.2015581412064
+       -90.52849135943048
+      -0.3710175116755678
+        217.9162663808141
+        505.7204469219135
+ 6.1e+10     
+           515.3304229662
+        218.4235957252802
+        469.1088976146855
+       -1.453548062069581
+        155.4149446728252
+        469.4268082836542
+       -91.09524163658948
+      -0.7025138531002622
+        218.5597498087689
+         507.185387266157
+ 6.11e+10    
+        516.8055845959406
+        219.0645287066306
+        470.3356171796858
+       -1.789210254645884
+        155.7825787774327
+        470.6542879950481
+       -91.66292475622332
+       -1.035784336661834
+         219.203188325564
+        508.6531967181135
+ 6.12e+10    
+        518.2836208617521
+        219.7054007812123
+        471.5645750231546
+        -2.12664699022119
+        156.1504698286928
+        471.8840015575927
+       -92.23152768689749
+       -1.370825605071508
+        219.8465777894213
+        510.1238825643393
+ 6.13e+10    
+        519.7645394255869
+        220.3462079603949
+        472.7957754800934
+       -2.465854742796591
+        156.5186217673156
+        473.1159533375276
+        -92.8010372695347
+       -1.707634184644672
+        220.4899142240182
+          511.59745232467
+ 6.14e+10    
+        521.2483481900831
+        220.9869464239996
+        474.0292229683852
+       -2.806829868614061
+        156.8870386141199
+         474.350147785882
+       -93.37144021745323
+       -2.046206484924227
+        221.1331938210104
+        513.0739137548337
+ 6.15e+10    
+        522.7350553012391
+        221.6276125228409
+        475.2649219895523
+       -3.149568605788867
+        157.2557244703696
+        475.5865894392293
+       -93.94272311642459
+       -2.386538798316735
+        221.7764129425623
+        514.5532748490368
+ 6.16e+10    
+         524.224669151097
+         222.268202781275
+         476.502877129498
+       -3.494067073951884
+        157.6246835181037
+        476.8252829204401
+       -94.51487242475029
+       -2.728627299736839
+        222.4195681238872
+          516.03554384258
+ 6.17e+10    
+        525.7171983804171
+        222.9087138997579
+        477.7430930592642
+       -3.840321273902184
+        157.9939200204687
+        478.0662329394441
+       -95.08787447335801
+       -3.072468046262857
+        223.0626560757981
+        517.5207292144594
+ 6.18e+10    
+        527.2126518813677
+        223.5491427574138
+        478.9855745357749
+       -4.188327087271405
+        158.3634383220409
+        479.3094442939782
+       -95.66171546591791
+       -3.418056976802797
+        223.7056736872651
+        519.0088396899695
+ 6.19e+10    
+        528.7110388002059
+        224.1894864146113
+         480.230326402594
+        -4.53808027619665
+        158.7332428491529
+        480.5549218703528
+       -96.23638147897731
+       -3.765389911770688
+        224.3486180279835
+        520.4998842433162
+ 6.2e+10     
+        530.2123685399682
+        224.8297421155499
+        481.4773535906756
+        -4.88957648300523
+        159.1033381102115
+        481.8026706442068
+       -96.81185846211545
+       -4.114462552772292
+        224.9914863509523
+        521.9938721002259
+ 6.21e+10    
+        531.7166507631523
+        225.4699072908531
+        482.7266611191181
+       -5.242811229909476
+         159.473728696015
+        483.0526956812649
+       -97.38813223811815
+       -4.465270482302817
+        225.6342760950582
+        523.4908127405573
+ 6.22e+10    
+        533.2238953944142
+        226.1099795601739
+         483.978254095922
+        -5.59777991871246
+        159.8444192800682
+        484.3050021381019
+         -97.965188503172
+       -4.817809163453679
+        226.2769848876726
+        524.9907159009161
+ 6.23e+10    
+        534.7341126232558
+        226.7499567348072
+        485.2321377187407
+       -5.954477830523514
+        160.2154146188911
+        485.5595952629026
+       -98.54301282707806
+       -5.172073939630597
+        226.9196105472541
+        526.4935915772679
+ 6.24e+10    
+        536.2473129067203
+          227.38983682031
+        486.4883172756415
+       -6.312900125484864
+         160.586719552328
+        486.8164803962211
+       -99.12159065348534
+       -5.528060034281333
+        227.5621510859607
+        527.9994500275542
+ 6.25e+10    
+        537.7635069720875
+        228.0296180191334
+        487.7467981458652
+       -6.673041842508438
+        160.9583390038527
+        488.0756629717491
+       -99.70090730014414
+       -5.885762550634093
+        228.2046047122739
+        529.5083017743146
+ 6.26e+10    
+        539.2827058195655
+        228.6692987332614
+        489.0075858005798
+       -7.034897899024491
+        161.3302779808677
+        489.3371485170734
+         -100.28094795918
+       -6.245176471447071
+        228.8469698336265
+        531.0201576073031
+ 6.27e+10    
+        540.8049207249976
+        229.3088775668566
+        490.2706858036429
+       -7.398463090738288
+        161.7025415750047
+        490.6009426544452
+       -100.8616976973861
+       -6.606296658767405
+        229.4892450590421
+        532.5350285861067
+ 6.28e+10    
+        542.3301632425556
+        229.9483533289183
+        491.5361038123643
+       -7.763732091399984
+        162.0751349624198
+        491.8670511015447
+        -101.443141456537
+       -6.969117853701015
+        230.1314292017833
+        534.0529260427761
+ 6.29e+10    
+        543.8584452074418
+        230.5877250359477
+        492.8038455782656
+       -8.130699452583604
+        162.4480634040841
+        493.1354796722454
+       -102.0252640537208
+       -7.333634676193038
+        230.7735212820068
+        535.5738615844388
+ 6.3e+10     
+        545.3897787385899
+        231.2269919146176
+        494.0739169478428
+        -8.49935960347737
+        162.8213322460739
+        494.4062342773819
+       -102.6080501816928
+       -7.699841624818397
+        231.4155205294284
+        537.0978470959319
+ 6.31e+10    
+        546.9241762413761
+        231.8661534044588
+        495.3463238633317
+       -8.869706850683428
+         163.194946919858
+        495.6793209255222
+       -103.1914844092484
+       -8.067733076583345
+        232.0574263859955
+        538.6248947424239
+ 6.32e+10    
+        548.4616504103152
+        232.5052091605477
+        496.6210723634771
+       -9.241735378029801
+        163.5689129425784
+        496.9547457237294
+        -103.775551181616
+       -8.437303286736709
+         232.699238508569
+        540.1550169720482
+ 6.33e+10    
+        550.0022142317724
+        233.1441590562019
+        497.8981685842854
+       -9.615439246391423
+        163.9432359173314
+        498.2325148783378
+       -104.3602348208688
+       -8.808546388591948
+        233.3409567716121
+        541.6882265185233
+ 6.34e+10    
+        551.5458809866685
+        233.7830031856914
+         499.177618759806
+       -9.990812393523235
+        164.3179215334438
+         499.512634695721
+       -104.9455195263599
+       -9.181456393360151
+        233.9825812698879
+        543.2245364037897
+ 6.35e+10    
+        553.0926642531909
+        234.4217418669499
+        500.4594292228915
+       -10.36784863390207
+        164.6929755667475
+        500.7951115830638
+       -105.5313893751726
+       -9.556027189992394
+        234.6241123211658
+        544.7639599406366
+ 6.36e+10    
+        554.6425779095048
+        235.0603756442972
+        501.7436064059672
+       -10.74654165858058
+        165.0684038798487
+        502.0799520491345
+       -106.1178283225944
+       -9.932252545033576
+        235.2655504689344
+        546.3065107353382
+ 6.37e+10    
+        556.1956361364565
+         235.698905291171
+         503.030156841803
+       -11.12688503505098
+        165.4442124223967
+        503.3671627050583
+       -106.7048202026103
+       -10.31012610248555
+        235.9068964851247
+        547.8522026902867
+ 6.38e+10    
+        557.7518534202995
+         236.337331812866
+        504.3190871642851
+       -11.50887220711974
+        165.8204072313474
+        504.6567502650942
+       -107.2923487284141
+       -10.68964138368221
+        236.5481513728389
+        549.4010500066195
+ 6.39e+10    
+        559.3112445553932
+        236.9756564492756
+        505.6104041091792
+       -11.89249649479234
+        166.1969944312245
+        505.9487215474048
+       -107.8803974929414
+       -11.07079178717295
+        237.1893163690883
+        550.9530671868665
+ 6.4e+10     
+         560.873824646928
+        237.6138806776517
+         506.904114514918
+       -12.27775109416865
+        166.5739802343785
+        507.2430834748386
+       -108.4689499694223
+       -11.45357058861856
+        237.8303929475381
+        552.5082690375776
+ 6.41e+10    
+        562.4396091136343
+        238.2520062153622
+         508.200225323361
+        -12.6646290773489
+        166.9513709412411
+         508.539843075701
+       -109.0579895119531
+       -11.83797094069566
+        238.4713828212618
+         554.066670671962
+ 6.42e+10    
+        564.0086136905057
+        238.8900350226624
+         509.498743580577
+       -13.05312339235074
+         167.329172940577
+        509.8390074845367
+       -109.6474993560886
+       -12.22398587301287
+        239.1122879455008
+        555.6282875125318
+ 6.43e+10    
+        565.5808544315108
+        239.5279693054704
+        510.7996764376168
+       -13.44322686303482
+        167.7073927097336
+        511.1405839429068
+       -110.2374626194532
+       -12.61160829203606
+        239.7531105204337
+        557.1931352937343
+ 6.44e+10    
+        567.1563477123098
+        240.1658115181515
+         512.103031151293
+       -13.83493218904318
+        168.0860368148864
+        512.4445798001683
+       -110.8278623023733
+       -13.00083098102536
+        240.3938529939506
+        558.7612300645943
+ 6.45e+10    
+         568.735110232982
+        240.8035643663115
+        513.4088150849524
+       -14.22823194574611
+        168.4651119112812
+        513.7510025142541
+       -111.4186812885269
+       -13.39164659998027
+        241.0345180644386
+        560.3325881913596
+ 6.46e+10    
+        570.3171590207364
+        241.4412308095924
+         514.717035709259
+       -14.62311858420081
+         168.844624743475
+        515.0598596524542
+       -112.0099023456158
+       -13.78404768559776
+        241.6751086835694
+        561.9072263601373
+ 6.47e+10    
+        571.9025114326411
+        242.0788140644823
+        516.0277006029726
+       -15.01958443111921
+        169.2245821455716
+        516.3711588922008
+       -112.6015081260544
+       -14.17802665123803
+        242.3156280591001
+        563.4851615795395
+ 6.48e+10    
+        573.4911851583345
+        242.7163176071249
+        517.3408174537277
+       -15.41762168884686
+        169.6049910414548
+        517.6849080218441
+       -113.1934811676794
+       -14.57357578690178
+        242.9560796576756
+        565.0664111833252
+ 6.49e+10    
+        575.0831982227608
+         243.353745176143
+        518.6563940588146
+       -15.81722243535152
+        169.9858584450201
+        519.0011149414479
+       -113.7858038944794
+       -14.97068725921751
+        243.5964672076423
+        566.6509928330476
+ 6.5e+10     
+        576.6785689888782
+        243.9911007754637
+        519.9744383259659
+       -16.21837862422285
+        170.3671914604009
+        520.3197876635602
+       -114.3784586173421
+       -15.36935311143835
+        244.2367947018675
+         568.238924520694
+ 6.51e+10    
+         578.277316160396
+        244.6283886771535
+        521.2949582741339
+       -16.62108208468086
+        170.7489972821938
+        521.6409343140131
+       -114.9714275348224
+       -15.76956526344995
+        244.8770664005635
+        569.8302245713371
+ 6.52e+10    
+        579.8794587844902
+        245.2656134242599
+        522.6179620342784
+       -17.02532452159679
+        171.1312831956783
+        522.9645631326953
+       -115.5646927339287
+       -16.17131551178714
+        245.5172868341221
+         571.424911645777
+ 6.53e+10    
+        581.4850162545303
+        245.9027798336574
+        523.9434578501493
+       -17.43109751552112
+        171.5140565770371
+        524.2906824743512
+       -116.1582361909277
+       -16.57459552966175
+        246.1574608059543
+        573.0230047431894
+ 6.54e+10    
+        583.0940083128053
+        246.5398929989043
+         525.271454079077
+       -17.83839252272413
+        171.8973248935694
+        525.6193008093621
+         -116.75203977217
+        -16.9793968669994
+        246.7975933953359
+        574.6245232037744
+ 6.55e+10    
+        584.7064550532494
+        247.1769582931011
+        526.6019591927524
+       -18.24720087524558
+         172.281095703904
+        526.9504267245352
+       -117.3460852349322
+       -17.38571095048701
+        247.4376899602607
+        576.2294867114027
+ 6.56e+10    
+        586.3223769241704
+        247.8139813717609
+        527.9349817780225
+       -18.65751378095445
+        172.6653766582083
+        528.2840689238994
+       -117.9403542282793
+       -17.79352908362961
+        248.0777561403011
+        577.8379152962663
+ 6.57e+10    
+        587.9417947309711
+        248.4509681756809
+        529.2705305376707
+       -19.06932232361858
+        173.0501754983938
+        529.6202362294855
+       -118.5348282939458
+       -18.20284244681776
+        248.7177978594716
+        579.4498293375249
+ 6.58e+10    
+        589.5647296388837
+        249.0879249338235
+        530.6086142912127
+       -19.48261746298402
+        173.4355000583193
+        530.9589375821264
+       -119.1294888672332
+       -18.61364209740296
+        249.3578213291042
+        581.0652495659574
+ 6.59e+10    
+        591.1912031756887
+        249.7248581662028
+        531.9492419756816
+       -19.89739003486439
+        173.8213582639919
+        532.3001820422469
+       -119.7243172779285
+       -19.02591896978521
+        249.9978330507251
+         582.684197066611
+ 6.6e+10     
+        592.8212372344516
+        250.3617746867774
+        533.2924226464239
+       -20.31363075124081
+         174.207758133762
+        533.6439787906518
+         -120.31929475124
+       -19.43966387550858
+        250.6378398189387
+        584.3066932814527
+ 6.61e+10    
+        594.4548540762462
+        250.9986816063486
+        534.6381654778876
+       -20.73133020037023
+        174.5947077785194
+        534.9903371293258
+       -120.9144024087496
+       -19.85486750336657
+        251.2778487243213
+        585.9327600120189
+ 6.62e+10    
+        596.0920763328843
+        251.6355863354654
+         535.986479764419
+       -21.15047884690414
+        174.9822154018831
+        536.3392664822262
+       -121.5096212693864
+       -20.27152041951772
+        251.9178671563163
+         587.562419422067
+ 6.63e+10    
+        597.7329270096428
+        252.2724965873344
+        537.3373749210486
+       -21.57106703201721
+        175.3702893003886
+        537.6907763960726
+       -122.1049322504137
+       -20.68961306761025
+        252.5579028061346
+        589.1956940402245
+ 6.64e+10    
+        599.3774294879946
+        252.9094203807359
+         538.690860484291
+       -21.99308497354488
+        175.7589378636749
+        539.0448765411506
+       -122.7003161684389
+         -21.109135768916
+        253.1979636696696
+        590.8326067626506
+ 6.65e+10    
+        601.0256075283403
+        253.5463660429471
+        540.0469461129431
+       -22.41652276613098
+        176.1481695746656
+        540.4015767121033
+        -123.295753740436
+       -21.53007872247442
+        253.8380580504044
+        592.4731808556728
+ 6.66e+10    
+        602.6774852727301
+        254.1833422126684
+        541.4056415888726
+       -22.84137038138498
+        176.5379930097464
+        541.7608868287278
+       -123.8912255847886
+        -21.9524320052451
+        254.4781945623371
+        594.1174399584507
+ 6.67e+10    
+        604.3330872476004
+        254.8203578429572
+        542.7669568178188
+       -23.26761766804713
+        176.9284168389446
+        543.1228169367787
+        -124.486712222349
+       -22.37618557227061
+        255.1183821329028
+         595.765408085624
+ 6.68e+10    
+        605.9924383664999
+         255.457422204165
+        544.1309018301864
+       -23.69525435216562
+        177.3194498260982
+        544.4873772087587
+       -125.0821940775148
+       -22.80132925684698
+        255.7586300059079
+        597.4171096299693
+ 6.69e+10    
+          607.65556393282
+        256.0945448868822
+        545.4974867818486
+       -24.12427003728041
+        177.7111008290305
+        545.8545779447256
+        -125.677651479322
+       -23.22785277070532
+        256.3989477444632
+         599.072569365044
+ 6.7e+10     
+        609.3224896425232
+        256.7317358048875
+        546.8667219549411
+       -24.55465420461791
+        178.1033787997135
+        547.2244295730845
+       -126.2730646625541
+       -23.65574570420063
+        257.0393452339283
+        600.7318124478514
+ 6.71e+10    
+         610.993241586875
+        257.3690051981013
+        548.2386177586656
+       -24.98639621329387
+        178.4962927844349
+        548.5969426513942
+       -126.8684137688701
+       -24.08499752651142
+         257.679832684856
+        602.3948644214806
+ 6.72e+10    
+        612.6678462551705
+        258.0063636355427
+         549.613184730083
+       -25.41948530052661
+         178.889851923958
+        549.9721278671661
+       -127.4636788479468
+       -24.51559758584685
+         258.320420635947
+        604.0617512177716
+ 6.73e+10    
+        614.3463305374646
+        258.6438220182979
+        550.9904335349225
+       -25.85391058185732
+        179.2840654536819
+        551.3499960386662
+       -128.0588398586375
+       -24.94753510966312
+         258.961119957004
+        605.7324991599604
+ 6.74e+10    
+        616.0287217273036
+        259.2813915824851
+        552.3703749683776
+        -26.2896610513811
+        179.6789427037951
+        552.7305581157153
+       -128.6538766701468
+       -25.38079920488938
+        259.6019418518949
+        607.4071349653358
+ 6.75e+10    
+        617.7150475244509
+        259.9190839022291
+        553.7530199559069
+       -26.72672558198579
+        180.0744930994306
+         554.113825180497
+       -129.2487690632227
+       -25.81537885816162
+        260.2428978615192
+        609.0856857478891
+ 6.76e+10    
+        619.4053360376191
+        260.5569108926406
+        555.1383795540413
+       -27.16509292560055
+        180.4707261608139
+        555.4998084483533
+       -129.8434967313622
+       -26.25126293606557
+        260.8839998667794
+        610.7681790209724
+ 6.77e+10    
+        621.0996157871915
+        261.1948848127972
+        556.5264649511845
+       -27.60475171345193
+        180.8676515034115
+        556.8885192685951
+       -130.4380392820338
+        -26.6884401853886
+        261.5252600915546
+        612.4546426999444
+ 6.78e+10    
+        622.7979157079653
+        261.8330182687313
+        557.9172874684137
+        -28.0456904563294
+        181.2652788380742
+        558.2799691253053
+       -131.0323762379134
+       -27.12689923337826
+        262.1666911056856
+        614.1451051048309
+ 6.79e+10    
+        624.5002651518596
+        262.4713242164211
+        559.3108585602902
+       -28.48789754485943
+        181.6636179711795
+        559.6741696381417
+       -131.6264870381384
+       -27.56662858801262
+        262.8083058279536
+        615.8395949629711
+ 6.8e+10     
+        626.2066938906604
+        263.1098159647854
+        560.7071898156565
+       -28.93136124978802
+        182.0626788047687
+        561.0711325631414
+       -132.2203510395726
+       -28.00761663827577
+        263.4501175290727
+        617.5381414116704
+ 6.81e+10    
+        627.9172321187385
+        263.7485071786844
+        562.1062929584497
+       -29.37606972227135
+        182.4624713366851
+        562.4708697935322
+       -132.8139475180898
+       -28.44985165444328
+        264.0921398346827
+        619.2407740008598
+ 6.82e+10    
+        629.6319104557792
+        264.3874118819239
+        563.5081798485006
+       -29.82201099417477
+        182.8630056607044
+        563.8733933605325
+       -133.4072556698686
+       -28.89332178837576
+        264.7343867283445
+        620.9475226957362
+ 6.83e+10    
+        631.3507599495065
+        265.0265444602584
+        564.9128624823386
+       -30.26917297838042
+        183.2642919666664
+         565.278715434162
+       -134.0002546127017
+       -29.33801507381979
+        265.3768725545427
+         622.658417879425
+ 6.84e+10    
+        633.0738120784166
+        265.6659196644086
+        566.3203529940062
+         -30.717543469103
+        183.6663405406027
+        566.6868483240499
+       -134.5929233873221
+       -29.78391942671846
+          266.01961202169
+        624.3734903556253
+ 6.85e+10    
+        634.8010987544932
+        266.3055526130721
+        567.7306636558606
+       -31.16711014221267
+        184.0691617648606
+        568.0978044802367
+       -135.1852409587384
+       -30.23102264552718
+        266.6626202051345
+        626.0927713512577
+ 6.86e+10    
+        636.5326523259359
+        266.9454587959418
+        569.1438068793773
+       -31.61786055556791
+        184.4727661182251
+        569.5115964939869
+       -135.7771862175886
+       -30.67931241154094
+        267.3059125501741
+        627.8162925191253
+ 6.87e+10    
+        638.2685055798892
+        267.5856540767294
+        570.5597952159665
+       -32.06978214935381
+        184.8771641760392
+        570.9282370985974
+       -136.3687379815021
+       -31.12877628922621
+        267.9495048750705
+        629.5440859405535
+ 6.88e+10    
+        640.0086917451625
+        268.2261546961903
+        571.9786413577751
+        -32.5228622464304
+        185.2823666103186
+        572.3477391701998
+       -136.9598749964783
+       -31.57940172656213
+        268.5934133740682
+        631.2761841280451
+ 6.89e+10    
+        641.7532444949487
+        268.8669772751504
+        573.4003581384959
+       -32.97708805268693
+         185.688384189868
+        573.7701157285795
+       -137.5505759382769
+       -32.03117605538937
+        269.2376546204186
+        633.0126200279282
+ 6.9e+10     
+        643.5021979495552
+        269.5081388175394
+        574.8249585341772
+       -33.43244665740526
+        186.0952277803897
+        575.1953799379773
+       -138.1408194138212
+       -32.48408649176595
+        269.8822455694037
+        634.7534270230035
+ 6.91e+10    
+        645.2555866791193
+        270.1496567134241
+        576.2524556640303
+       -33.88892503362967
+         186.502908344594
+        576.6235451078978
+        -138.730583962611
+       -32.93812013633047
+        270.5272035613642
+        636.4986389351922
+ 6.92e+10    
+        647.0134457063306
+        270.7915487420461
+        577.6828627912416
+       -34.34651003854552
+        186.9114369423041
+        578.0546246939259
+       -139.3198480581522
+       -33.39326397467349
+        271.1725463247346
+        638.2482900281894
+ 6.93e+10    
+        648.7758105091524
+        271.4338330748607
+        579.1161933237763
+       -34.80518841386262
+        187.3208247305594
+        579.4886322985282
+        -139.908590109394
+        -33.8495048777155
+         271.818291979072
+         640.002415010101
+ 6.94e+10    
+        650.5427170235372
+        272.0765282785831
+        580.5524608151946
+       -35.26494678620945
+        187.7310829637163
+        580.9255816718709
+         -140.49678846218
+       -34.30682960209207
+        272.4644590380984
+        641.7610490360978
+ 6.95e+10    
+        652.3142016461516
+        272.7196533182275
+         581.991678965457
+       -35.72577166753182
+        188.1422229935465
+        582.3654867126231
+       -141.0844214007092
+       -34.76522479054617
+        273.1110664127372
+        643.5242277110582
+ 6.96e+10    
+        654.0903012370842
+        273.3632275601611
+        583.4338616217369
+       -36.18764945549948
+        188.5542562693314
+        583.8083614687721
+         -141.67146714901
+       -35.22467697232808
+         273.758133414156
+        645.2919870922108
+ 6.97e+10    
+        655.8710531225677
+        274.0072707751492
+        584.8790227792254
+       -36.65056643391985
+        188.9671943379559
+        585.2542201384299
+       -142.2579038724209
+       -35.68517256360109
+        274.4056797568108
+        647.0643636917815
+ 6.98e+10    
+        657.6564950976986
+        274.6518031414097
+        586.3271765819491
+       -37.11450877315879
+         189.381048843998
+         586.703077070646
+       -142.8437096790881
+        -36.1466978678549
+        275.0537255614945
+        648.8413944796386
+ 6.99e+10    
+        659.4466654291384
+        275.2968452476656
+        587.7783373235729
+        -37.5794625305678
+        189.7958315298166
+        588.1549467662171
+        -143.428862621466
+       -36.60923907632507
+        275.7022913583829
+        650.6231168859276
+ 7e+10       
+        661.2416028578411
+         275.942418096203
+        589.2325194482166
+       -38.04541365091759
+        190.2115542356375
+        589.6098438784957
+       -144.0133406978339
+       -37.07278226841991
+        276.3513980900868
+        652.4095688037188
* NOTE: Solution at 1e+08 Hz used as DC point.

.model l_m4lines_HFSS_W_1 sp N=4 SPACING=nonuniform VALTYPE=real
+ INTERPOLATION=spline
+ INFINITY =
+    4.771275496612187e-07
+    1.992620892018445e-07
+    4.599493106995181e-07
+    6.333700301101069e-08
+    1.283548577953231e-07
+    4.599264508819013e-07
+    2.830257265266555e-08
+    6.339692795622215e-08
+    1.993667267423742e-07
+    4.775330895971331e-07
+ DATA = 700
+ 0           
+    4.187375639716964e-07
+    1.499780296080442e-07
+    4.160104447847029e-07
+    4.559175281127766e-08
+      9.3362516970571e-08
+    4.159107655224221e-07
+    2.474797370846747e-08
+    4.559883258452768e-08
+    1.500178654245671e-07
+     4.18915896522694e-07
+ 2e+08       
+    4.152409295458201e-07
+    1.496357305871249e-07
+    4.124619577225161e-07
+    4.548151148332848e-08
+      9.2913481972087e-08
+    4.123676835644636e-07
+    2.471316967566081e-08
+    4.548809260884237e-08
+    1.496823467245008e-07
+    4.154633204210293e-07
+ 3e+08       
+    4.136486656757639e-07
+    1.495163480809376e-07
+    4.108544222836318e-07
+    4.542229773637365e-08
+    9.271611584391797e-08
+    4.107642254925401e-07
+    2.469173623432938e-08
+    4.542794895367581e-08
+    1.495623570531414e-07
+    4.138979002356905e-07
+ 4e+08       
+    4.127491121110181e-07
+    1.494674564879319e-07
+    4.099434383939512e-07
+    4.539229528127803e-08
+    9.260776279126221e-08
+    4.098566144861343e-07
+    2.468312840559359e-08
+    4.539725852963568e-08
+    1.495126419631506e-07
+    4.130184879975287e-07
+ 5e+08       
+    4.121313746128284e-07
+    1.494315581240394e-07
+    4.093168219391762e-07
+    4.537387643230625e-08
+    9.253361250161293e-08
+    4.092328666957902e-07
+    2.467882915622239e-08
+    4.537829677420827e-08
+    1.494763879888115e-07
+    4.124167743840308e-07
+ 6e+08       
+    4.116606371114502e-07
+    1.493998803351824e-07
+    4.088397915546797e-07
+     4.53606269268681e-08
+    9.247712803445569e-08
+    4.087582166247306e-07
+    2.467580053249492e-08
+    4.536458521887698e-08
+    1.494446090073347e-07
+     4.11959011756301e-07
+ 7e+08       
+    4.112849431016661e-07
+    1.493727465672836e-07
+    4.084597465168611e-07
+    4.535032585077475e-08
+    9.243225166966005e-08
+    4.083801157525448e-07
+    2.467331398647141e-08
+    4.535388116828527e-08
+    1.494174616029349e-07
+    4.115940282130534e-07
+ 8e+08       
+    4.109786239826518e-07
+     1.49350648695808e-07
+    4.081501796886804e-07
+    4.534212976387202e-08
+    9.239595057502099e-08
+    4.080721446939833e-07
+    2.467133421986299e-08
+    4.534533432088021e-08
+    1.493953604773808e-07
+    4.112967749299486e-07
+ 9e+08       
+    4.107254835411902e-07
+    1.493331689259142e-07
+    4.078942439898151e-07
+    4.533562699302215e-08
+    9.236622925020992e-08
+    4.078175450740826e-07
+    2.466995580577002e-08
+     4.53385281155439e-08
+    1.493778561619893e-07
+    4.110514931708178e-07
+ 1e+09       
+    4.105136024924595e-07
+    1.493193440705552e-07
+    4.076796662179595e-07
+    4.533053841996527e-08
+    9.234158265688879e-08
+    4.076041127226923e-07
+     2.46692448524731e-08
+    4.533317717036472e-08
+    1.493639705729949e-07
+    4.108465377447294e-07
+ 1.1e+09     
+    4.104202826859234e-07
+    1.493538769171751e-07
+    4.075820137037365e-07
+    4.531579175664737e-08
+    9.234113385434064e-08
+    4.075073361738556e-07
+    2.466258577860408e-08
+    4.531862601988128e-08
+    1.493987214278646e-07
+    4.107588020961512e-07
+ 1.2e+09     
+    4.103238980288448e-07
+    1.493785811622875e-07
+    4.074810590166204e-07
+    4.530205008188562e-08
+    9.233653225599419e-08
+    4.074072430350871e-07
+    2.465589816739153e-08
+    4.530497437721173e-08
+    1.494236503247642e-07
+    4.106678947755146e-07
+ 1.3e+09     
+    4.102259598345665e-07
+    1.493951101007474e-07
+    4.073785504595165e-07
+    4.528950340605285e-08
+    9.232912804855798e-08
+    4.073055678820231e-07
+    2.464936279794644e-08
+    4.529244045001071e-08
+    1.494404081271479e-07
+    4.105752602259324e-07
+ 1.4e+09     
+    4.101277841760492e-07
+    1.494050094749475e-07
+    4.072759723649872e-07
+    4.527826320559618e-08
+    9.231992394244825e-08
+    4.072037841359851e-07
+    2.464313904757545e-08
+    4.528115806342246e-08
+    1.494505361749364e-07
+    4.104821632982791e-07
+ 1.5e+09     
+    4.100304824083551e-07
+    1.494096589630412e-07
+    4.071745509299042e-07
+    4.526838848027486e-08
+    9.230967142774388e-08
+     4.07103109924019e-07
+     2.46373647754362e-08
+    4.527120323443528e-08
+    1.494554090837679e-07
+    4.103896787362664e-07
+ 1.6e+09     
+    4.099349669312446e-07
+    1.494102535558261e-07
+    4.070752719102485e-07
+    4.525990342525768e-08
+    9.229893704502655e-08
+    4.070045255850295e-07
+    2.463215732993045e-08
+    4.526261274670229e-08
+    1.494562169800732e-07
+    4.102986953523529e-07
+ 1.7e+09     
+    4.098419660795698e-07
+    1.494078070818759e-07
+    4.069789050511995e-07
+    4.525280929947188e-08
+    9.228814900220803e-08
+    4.069087977833684e-07
+    2.462761510928252e-08
+    4.525539696795348e-08
+     1.49453969510951e-07
+    4.102099290325914e-07
+ 1.8e+09     
+    4.097520438277476e-07
+    1.494031668981093e-07
+    4.068860315224332e-07
+    4.524709238233046e-08
+    9.227763073114043e-08
+    4.068165065683095e-07
+    2.462381935860325e-08
+     4.52495486502576e-08
+    1.494495107504464e-07
+    4.101239404646812e-07
+ 1.9e+09     
+    4.096656213733883e-07
+    1.493970332557593e-07
+    4.067970717828267e-07
+    4.524272933089763e-08
+    9.226762557850397e-08
+     4.06728072852418e-07
+    2.462083602864691e-08
+    4.524504897610135e-08
+    1.494435386060059e-07
+    4.100411548074913e-07
+ 2e+09       
+    4.095829986845196e-07
+    1.493899796828038e-07
+    4.067123122019413e-07
+    4.523969081685297e-08
+    9.225831532476957e-08
+    4.066437846677075e-07
+    2.461871759883096e-08
+    4.524187173044978e-08
+    1.494366251384291e-07
+    4.099618814864822e-07
+ 2.1e+09     
+    4.095043748311024e-07
+    1.493824724444589e-07
+    4.066319294440564e-07
+    4.523794402081901e-08
+    9.224983429257445e-08
+    4.065638212233825e-07
+    2.461750480957951e-08
+    4.523998619743759e-08
+    1.494292359076047e-07
+    4.098863329909699e-07
+ 2.2e+09     
+    4.094298664416369e-07
+    1.493748881587196e-07
+    4.065560121111569e-07
+    4.523745435972639e-08
+    9.224228022392194e-08
+    4.064882742697863e-07
+    2.461722827330788e-08
+    4.523935918368662e-08
+    1.494217474540465e-07
+    4.098146420352995e-07
+ 2.3e+09     
+    4.093595239833183e-07
+    1.493675292252325e-07
+    4.064845794812584e-07
+    4.523818669136903e-08
+    9.223572273792599e-08
+    4.064171666066133e-07
+    2.461790994809888e-08
+    4.523995643717883e-08
+     1.49414462594482e-07
+    4.097468767800577e-07
+ 2.4e+09     
+    4.092933458013594e-07
+    1.493606370454434e-07
+    4.064175974018921e-07
+    4.524010615597025e-08
+    9.223020994405208e-08
+    4.063504677927401e-07
+     2.46195644676736e-08
+    4.524174364227123e-08
+    1.494076235203583e-07
+    4.096830540317826e-07
+ 2.5e+09     
+    4.092312900023529e-07
+    1.493544031765728e-07
+    4.063549915346874e-07
+    4.524317876088124e-08
+    9.222577362951162e-08
+    4.062881072488879e-07
+    2.462220032775121e-08
+    4.524468711332486e-08
+    1.494014228468374e-07
+    4.096231504808623e-07
+ 2.6e+09     
+    4.091732843531386e-07
+    1.493489786364307e-07
+    4.062966582201646e-07
+    4.524737178030726e-08
+    9.222243333326686e-08
+    4.062299850164576e-07
+    2.462582093337697e-08
+    4.524875427123748e-08
+    1.493960128306666e-07
+    4.095671121207048e-07
+ 2.7e+09     
+    4.091192344097723e-07
+    1.493444815994441e-07
+    4.062424732614232e-07
+    4.525265401994389e-08
+    9.222019954465399e-08
+    4.061759804652776e-07
+    2.463042551483398e-08
+     4.52539139619256e-08
+    1.493915129965701e-07
+    4.095148620343854e-07
+ 2.8e+09     
+      4.0906903010528e-07
+    1.493410037198305e-07
+    4.061922989263223e-07
+    4.525899598200881e-08
+    9.221907621081529e-08
+    4.061259592441941e-07
+    2.463600992169181e-08
+    4.526013665890548e-08
+    1.493880164062954e-07
+    4.094663067510442e-07
+ 2.9e+09     
+    4.090225510205294e-07
+    1.493386152994094e-07
+    4.061459894510836e-07
+    4.526636995651833e-08
+    9.221906269712533e-08
+    4.060797787523517e-07
+     2.46425673056276e-08
+    4.526739458060899e-08
+    1.493855947855661e-07
+    4.094213413728973e-07
+ 3e+09       
+    4.089796705472651e-07
+    1.493373694930812e-07
+     4.06103395301828e-07
+    4.527475005801593e-08
+      9.2220155314337e-08
+    4.060372923832822e-07
+    2.465008870308562e-08
+    4.527566174505443e-08
+    1.493843026996699e-07
+    4.093798536618128e-07
+ 3.1e+09     
+    4.089402591313958e-07
+    1.493373057190685e-07
+    4.060643664198978e-07
+    4.528411222224441e-08
+    9.222234850255064e-08
+    4.059983527639739e-07
+    2.465856352878247e-08
+    4.528491397878002e-08
+    1.493841809426332e-07
+    4.093417272567898e-07
+ 3.2e+09     
+    4.089041867614537e-07
+    1.493384524160676e-07
+    4.060287546453749e-07
+    4.529443417379594e-08
+    9.222563574351245e-08
+    4.059628141803072e-07
+    2.466797999065842e-08
+    4.529512889278028e-08
+    1.493852592802277e-07
+    4.093068441736196e-07
+ 3.3e+09     
+    4.088713248440005e-07
+    1.493408292666858e-07
+    4.059964154831658e-07
+    4.530569537317489e-08
+    9.223001025795967e-08
+    4.059305343508222e-07
+    2.467832543623307e-08
+    4.530628583507808e-08
+    1.493875586645733e-07
+    4.092750867176215e-07
+ 3.4e+09     
+    4.088415475859615e-07
+    1.493444489864686e-07
+    4.059672093486232e-07
+    4.531787694970617e-08
+    9.223546553287671e-08
+    4.059013756838879e-07
+    2.468958663953842e-08
+    4.531836582720742e-08
+    1.493910930183107e-07
+    4.092463389209088e-07
+ 3.5e+09     
+     4.08814732984097e-07
+    1.493493187604916e-07
+    4.059410024053749e-07
+    4.533096162515272e-08
+    9.224199571395571e-08
+    4.058752061294919e-07
+      2.4701750036943e-08
+    4.533135149005863e-08
+    1.493958706692399e-07
+    4.092204875978277e-07
+ 3.6e+09     
+    4.087907635044283e-07
+     1.49355441394795e-07
+     4.05917667087087e-07
+    4.534493363166005e-08
+     9.22495958908008e-08
+    4.058518997162644e-07
+    2.471480191930069e-08
+    4.534522696311692e-08
+     1.49401895501852e-07
+    4.091974230964375e-07
+ 3.7e+09     
+    4.087695265193804e-07
+    1.493628162376011e-07
+    4.058970823770488e-07
+     4.53597786266452e-08
+    9.225826229608253e-08
+    4.058313368468175e-07
+    2.472872858699275e-08
+    4.535997781999908e-08
+    1.494091678800329e-07
+    4.091770398101203e-07
+ 3.8e+09     
+    4.087509145576472e-07
+    1.493714399149974e-07
+    4.058791339045584e-07
+    4.537548360643753e-08
+    9.226799243465396e-08
+    4.058134044097934e-07
+    2.474351647360775e-08
+    4.537559098229628e-08
+    1.494176853851136e-07
+    4.091592365016814e-07
+ 3.9e+09     
+    4.087348254110721e-07
+    1.493813069173055e-07
+    4.058637139047522e-07
+    4.539203681981971e-08
+    9.227878515434993e-08
+    4.057979957548497e-07
+    2.475915224323742e-08
+    4.539205463301175e-08
+    1.494274434051084e-07
+    4.091439164823729e-07
+ 4e+09       
+    4.087211621339423e-07
+     1.49392410065391e-07
+    4.058507210783854e-07
+    4.540942768207498e-08
+    9.229064066661864e-08
+     4.05785010566824e-07
+    2.477562286566318e-08
+    4.540935813029554e-08
+    1.494384356041157e-07
+    4.091309876799879e-07
+ 4.1e+09     
+    4.087098329627925e-07
+    1.494047408804887e-07
+    4.058400603798532e-07
+    4.542764668970406e-08
+    9.230356052215821e-08
+    4.057743546671986e-07
+    2.479291567307586e-08
+    4.542749192170782e-08
+     1.49450654295255e-07
+    4.091203626233454e-07
+ 4.2e+09     
+    4.087007511788457e-07
+    1.494182898764783e-07
+    4.058316427551019e-07
+    4.544668533561009e-08
+    9.231754754423921e-08
+    4.057659397644145e-07
+     2.48110184014063e-08
+    4.544644745885507e-08
+    1.494640907359334e-07
+    4.091119583648378e-07
+ 4.3e+09     
+    4.086938349303913e-07
+    1.494330467897795e-07
+    4.058253848457408e-07
+    4.546653602425919e-08
+    9.233260572034684e-08
+    4.057596831693298e-07
+    2.482991921884824e-08
+    4.546621711193827e-08
+    1.494787353605221e-07
+    4.091056963581579e-07
+ 4.4e+09     
+    4.086890070284965e-07
+    1.494490007589947e-07
+    4.058212086714781e-07
+    4.548719198609819e-08
+    9.234874005114241e-08
+     4.05755507487924e-07
+    2.484960674372229e-08
+    4.548679408351688e-08
+    1.494945779625051e-07
+    4.091015023045944e-07
+ 4.5e+09     
+    4.086861947263421e-07
+    1.494661404639604e-07
+     4.05819041299644e-07
+    4.550864719035836e-08
+    9.236595635454792e-08
+    4.057533403000695e-07
+    2.487007005345912e-08
+     4.55081723206311e-08
+    1.495116078357358e-07
+    4.090993059783002e-07
+ 4.6e+09     
+    4.086853294899889e-07
+    1.494844542319057e-07
+    4.058188145080369e-07
+     4.55308962552967e-08
+    9.238426102205835e-08
+     4.05753113830647e-07
+    2.489129868616767e-08
+     4.55303464243447e-08
+    1.495298138824844e-07
+     4.09099041038543e-07
+ 4.7e+09     
+    4.086863467664257e-07
+    1.495039301168474e-07
+    4.058204644454064e-07
+    4.555393435494522e-08
+    9.240366072426511e-08
+    4.057547646173701e-07
+    2.491328263599811e-08
+    4.555331155578428e-08
+    1.495491846944044e-07
+    4.091006448350487e-07
+ 4.8e+09     
+    4.086891857532065e-07
+     1.49524555957117e-07
+    4.058239312925019e-07
+    4.557775712156647e-08
+    9.242416206316626e-08
+    4.057582331783373e-07
+    2.493601234330824e-08
+    4.557706333787823e-08
+    1.495697086113278e-07
+    4.091040582110345e-07
+ 4.9e+09     
+    4.086937891728094e-07
+    1.495463194149778e-07
+    4.058291589257685e-07
+    4.560236054327728e-08
+     9.24457711702715e-08
+    4.057634636814472e-07
+    2.495947868049514e-08
+    4.560159775225983e-08
+    1.495913737618602e-07
+    4.091092253073547e-07
+ 5e+09       
+    4.087001030539148e-07
+    1.495692080015831e-07
+    4.058360945853136e-07
+    4.562774085672047e-08
+    9.246849325192686e-08
+    4.057704036173788e-07
+    2.498367293425998e-08
+     4.56269110312166e-08
+    1.496141680890499e-07
+    4.091160933702753e-07
+ 5.1e+09     
+    4.087080765211242e-07
+    1.495932090900352e-07
+    4.058446885487346e-07
+    4.565389443525468e-08
+     9.24923320867915e-08
+    4.057790034777925e-07
+    2.500858678503305e-08
+    4.565299954515777e-08
+    1.496380793639137e-07
+    4.091246125646829e-07
+ 5.2e+09     
+    4.087176615941278e-07
+    1.496183099189963e-07
+    4.058548938127371e-07
+    4.568081767390155e-08
+    9.251728948503657e-08
+    4.057892164407469e-07
+    2.503421228429499e-08
+    4.567985968684198e-08
+    1.496630951892949e-07
+    4.091347357940314e-07
+ 5.3e+09     
+    4.087288129969606e-07
+    1.496444975891359e-07
+     4.05866665785082e-07
+    4.570850687322205e-08
+    9.254336472451398e-08
+    4.058009980659339e-07
+    2.506054183058369e-08
+    4.570748775453862e-08
+    1.496892029963643e-07
+    4.091464185279262e-07
+ 5.4e+09     
+    4.087414879777481e-07
+    1.496717590546601e-07
+    4.058799619902874e-07
+    4.573695812534938e-08
+    9.257055398560428e-08
+    4.058143060032072e-07
+    2.508756814506561e-08
+    4.573587983735425e-08
+    1.497163900360328e-07
+     4.09159618638007e-07
+ 5.5e+09     
+    4.087556461391599e-07
+    1.497000811122043e-07
+    4.058947417934993e-07
+    4.576616720650743e-08
+    9.259884981321986e-08
+    4.058290997188821e-07
+    2.511528424765979e-08
+    4.576503170705702e-08
+    1.497446433675838e-07
+    4.091742962425735e-07
+ 5.6e+09     
+    4.087712492796959e-07
+    1.497294503894423e-07
+    4.059109661479214e-07
+    4.579612948137131e-08
+    9.262824064075847e-08
+    4.058453402452312e-07
+     2.51436834348116e-08
+    4.579493872176047e-08
+    1.497739498469026e-07
+    4.091904135602996e-07
+ 5.7e+09     
+    4.087882612458661e-07
+    1.497598533358198e-07
+    4.059285973719765e-07
+    4.582683982542724e-08
+    9.265871041571115e-08
+    4.058629899593995e-07
+    2.517275926009542e-08
+    4.582559574763003e-08
+    1.498042961167303e-07
+    4.092079347732815e-07
+ 5.8e+09     
+    4.088066477952431e-07
+    1.497912762177886e-07
+    4.059475989627292e-07
+    4.585829257187629e-08
+    9.269023836897096e-08
+    4.058820123983109e-07
+    2.520250551884756e-08
+    4.585699710516303e-08
+    1.498356686013462e-07
+    4.092268258995951e-07
+ 5.9e+09     
+    4.088263764703481e-07
+    1.498237051207579e-07
+    4.059679354518679e-07
+    4.589048148941809e-08
+    9.272279896849879e-08
+    4.059023721158875e-07
+    2.523291623796485e-08
+    4.588913654638515e-08
+    1.498680535079129e-07
+    4.092470546754612e-07
+ 6e+09       
+    4.088474164831929e-07
+    1.498571259596207e-07
+    4.059895723094691e-07
+    4.592339979628763e-08
+    9.275636209190682e-08
+     4.05924034587852e-07
+    2.526398567182075e-08
+    4.592200726834258e-08
+    1.499014368363656e-07
+    4.092685904470076e-07
+ 6.1e+09     
+    4.088697386102286e-07
+     1.49891524499151e-07
+    4.060124758988596e-07
+    4.595704021412447e-08
+    9.279089344121714e-08
+    4.059469661674466e-07
+    2.529570830493868e-08
+    4.595560196647562e-08
+    1.499358043991594e-07
+    4.092914040714927e-07
+ 6.2e+09     
+    4.088933150972559e-07
+    1.499268863847879e-07
+    4.060366134830974e-07
+    4.599139506266215e-08
+    9.282635520675233e-08
+    4.059711340926153e-07
+    2.532807886162541e-08
+    4.598991292886582e-08
+    1.499711418514123e-07
+    4.093154678276763e-07
+ 6.3e+09     
+    4.089181195736908e-07
+    1.499631971833861e-07
+    4.060619532801327e-07
+     4.60264563930148e-08
+    9.286270696693983e-08
+    4.059965065417498e-07
+    2.536109232223321e-08
+    4.602493216913672e-08
+    1.500074347310431e-07
+    4.093407553348235e-07
+ 6.4e+09     
+     4.08944126975368e-07
+    1.500004424325026e-07
+    4.060884645599764e-07
+    4.606221615383864e-08
+    9.289990678880976e-08
+    4.060230527313307e-07
+     2.53947439451425e-08
+    4.606065159228734e-08
+    1.500446685074925e-07
+    4.093672414796303e-07
+ 6.5e+09     
+    4.089713134748844e-07
+    1.500386076958248e-07
+    4.061161177735898e-07
+    4.609866638129299e-08
+     9.29379124728876e-08
+    4.060507430452065e-07
+    2.542902929300582e-08
+    4.609706318438331e-08
+    1.500828286366504e-07
+    4.093949023501468e-07
+ 6.6e+09     
+    4.089996564183379e-07
+    1.500776786215622e-07
+    4.061448847002984e-07
+    4.613579940101421e-08
+    9.297668286910494e-08
+    4.060795491823401e-07
+    2.546394426134825e-08
+     4.61341592143167e-08
+    1.501219006188341e-07
+    4.094237151756371e-07
+ 6.7e+09     
+    4.090291342672457e-07
+    1.501176410001547e-07
+    4.061747385988234e-07
+    4.617360802868612e-08
+    9.301617918005863e-08
+    4.061094443081157e-07
+    2.549948510735133e-08
+    4.617193243421753e-08
+    1.501618700561846e-07
+    4.094536582712179e-07
+ 6.8e+09     
+    4.090597265444253e-07
+    1.501584808175565e-07
+    4.062056543467554e-07
+    4.621208575554942e-08
+     9.30563661663469e-08
+      4.0614040319407e-07
+    2.553564847660353e-08
+    4.621037626485716e-08
+    1.502027227057642e-07
+    4.094847109861263e-07
+ 6.9e+09     
+    4.090914137827329e-07
+    1.502001843006944e-07
+    4.062376085546886e-07
+    4.625122690643162e-08
+    9.309721317639995e-08
+    4.061724023322617e-07
+    2.557243142579845e-08
+    4.624948495362591e-08
+    1.502444445249669e-07
+    4.095168536545624e-07
+ 7e+09       
+    4.091241774757241e-07
+    1.502427379523943e-07
+    4.062705796440134e-07
+    4.629102676044681e-08
+    9.313869493924671e-08
+    4.062054200133021e-07
+    2.560983143977325e-08
+    4.628925369523709e-08
+    1.502870217065618e-07
+    4.095500675482188e-07
+ 7.1e+09     
+     4.09158000029542e-07
+    1.502861285740522e-07
+    4.063045478812187e-07
+    4.633148162804779e-08
+    9.318079208075042e-08
+    4.062394363609079e-07
+    2.564784644184897e-08
+    4.632967870884547e-08
+    1.503304407016603e-07
+    4.095843348298478e-07
+ 7.2e+09     
+    4.091928647156146e-07
+    1.503303432754276e-07
+    4.063394953658844e-07
+    4.637258888210278e-08
+    9.322349134881954e-08
+    4.062744333201719e-07
+    2.568647479707667e-08
+    4.637075726926206e-08
+    1.503746882300076e-07
+      4.0961963850748e-07
+ 7.3e+09     
+    4.092287556239809e-07
+    1.503753694720244e-07
+    4.063754059738074e-07
+    4.641434694457227e-08
+    9.326678555755506e-08
+    4.063103946009922e-07
+    2.572571530862236e-08
+    4.641248769385387e-08
+    1.504197512780835e-07
+    4.096559623891668e-07
+ 7.4e+09     
+    4.092656576173142e-07
+    1.504211948714511e-07
+    4.064122652603054e-07
+    4.645675523369895e-08
+    9.331067328121739e-08
+    4.063473055817362e-07
+    2.576556720806007e-08
+    4.645486929005751e-08
+    1.504656170864266e-07
+    4.096932910383204e-07
+ 7.5e+09     
+    4.093035562858608e-07
+    1.504678074508332e-07
+    4.064500603314332e-07
+    4.649981407905858e-08
+    9.335515834418185e-08
+     4.06385153180862e-07
+    2.580603014073476e-08
+    4.649790227087338e-08
+    1.505122731282745e-07
+    4.097316097299255e-07
+ 7.6e+09     
+    4.093424379036222e-07
+    1.505151954277323e-07
+    4.064887796923387e-07
+    4.654352461319751e-08
+    9.340024916172276e-08
+    4.064239257057408e-07
+    2.584710414757672e-08
+    4.654158764708753e-08
+    1.505597070819987e-07
+    4.097709044079605e-07
+ 7.7e+09     
+    4.093822893861435e-07
+    1.505633472271289e-07
+    4.065284130823865e-07
+    4.658788864892469e-08
+    9.344595798864494e-08
+    4.064636126883193e-07
+    2.588878964480273e-08
+    4.658592710531006e-08
+     1.50607906799913e-07
+    4.098111616444247e-07
+ 7.8e+09     
+      4.0942309825026e-07
+    1.506122514468702e-07
+    4.065689513061149e-07
+    4.663290855078723e-08
+    9.349230012945879e-08
+    4.065042047166916e-07
+    2.593108740285069e-08
+    4.663092288038301e-08
+    1.506568602758794e-07
+    4.098523686003373e-07
+ 7.9e+09     
+    4.094648525760839e-07
+    1.506618968236682e-07
+    4.066103860678542e-07
+    4.667858710808546e-08
+    9.353929315647189e-08
+    4.065456932704162e-07
+      2.5973998525703e-08
+    4.667657762953628e-08
+      1.5070655561382e-07
+    4.098945129890204e-07
+ 8e+09       
+     4.09507540971441e-07
+    1.507122722012888e-07
+     4.06652709816165e-07
+    4.672492741523335e-08
+    9.358695617250918e-08
+    4.065880705657425e-07
+    2.601752443150194e-08
+    4.672289431412051e-08
+    1.507569809988008e-07
+    4.099375830418906e-07
+ 8.1e+09     
+    4.095511525388789e-07
+    1.507633665021233e-07
+    4.066959156024772e-07
+    4.677193276359658e-08
+    9.363530914451711e-08
+    4.066313294151376e-07
+    2.606166683508899e-08
+    4.676987609307241e-08
+    1.508081246718998e-07
+    4.099815674768974e-07
+ 8.2e+09     
+    4.095956768452657e-07
+    1.508151687028703e-07
+    4.067399969565853e-07
+    4.681960654733223e-08
+    9.368437232427126e-08
+    4.066754631037784e-07
+    2.610642773283784e-08
+     4.68175262306583e-08
+    1.508599749096131e-07
+     4.10026455469646e-07
+ 8.3e+09     
+    4.096411038939411e-07
+    1.508676678146731e-07
+    4.067849477801544e-07
+    4.686795218434622e-08
+    9.373416576362626e-08
+    4.067204652841617e-07
+    2.615180938992273e-08
+    4.686584801963548e-08
+    1.509125200081684e-07
+     4.10072236627184e-07
+ 8.4e+09     
+     4.09687424099303e-07
+    1.509208528677399e-07
+    4.068307622581827e-07
+    4.691697305234978e-08
+    9.378470892467842e-08
+     4.06766329888794e-07
+    2.619781432997801e-08
+    4.691484471983358e-08
+    1.509657482727924e-07
+    4.101189009643458e-07
+ 8.5e+09     
+    4.097346282636889e-07
+    1.509747129002346e-07
+    4.068774347874695e-07
+    4.696667243915325e-08
+    9.383602037997868e-08
+    4.068130510600121e-07
+    2.624444532696726e-08
+    4.696451951131679e-08
+    1.510196480117475e-07
+    4.101664388825261e-07
+ 8.6e+09     
+    4.097827075563597e-07
+    1.510292369510738e-07
+     4.06924959920552e-07
+    4.701705350576906e-08
+     9.38881175944458e-08
+    4.068606230954044e-07
+    2.629170539898632e-08
+    4.701487546072037e-08
+     1.51074207534795e-07
+    4.102148411507124e-07
+ 8.7e+09     
+    4.098316534944032e-07
+    1.510844140561733e-07
+    4.069733323232308e-07
+    4.706811926056931e-08
+    9.394101677864521e-08
+    4.069090404069636e-07
+    2.633959780366949e-08
+    4.706591549902743e-08
+    1.511294151556453e-07
+     4.10264098888594e-07
+ 8.8e+09     
+    4.098814579253608e-07
+    1.511402332476461e-07
+    4.070225467436885e-07
+    4.711987254260525e-08
+    9.399473280231437e-08
+    4.069582974919705e-07
+    2.638812603484327e-08
+     4.71176424089148e-08
+    1.511852591979252e-07
+    4.103142035515659e-07
+ 8.9e+09     
+    4.099321130113789e-07
+    1.511966835554628e-07
+    4.070725979912127e-07
+    4.717231601219859e-08
+    9.404927915711642e-08
+    4.070083889136387e-07
+    2.643729382006884e-08
+    4.717005881979667e-08
+    1.512417280041854e-07
+    4.103651469174477e-07
+ 9e+09       
+     4.09983611214722e-07
+    1.512537540111057e-07
+    4.071234809226784e-07
+    4.722545214701104e-08
+    9.410466795830811e-08
+     4.07059309289675e-07
+    2.648710511872723e-08
+    4.722316720879156e-08
+    1.512988099475043e-07
+    4.104169210747473e-07
+ 9.1e+09     
+    4.100359452844671e-07
+       1.513114336528e-07
+    4.071751904351263e-07
+    4.727928324195023e-08
+    9.416090997607085e-08
+    4.071110532870864e-07
+    2.653756412032067e-08
+    4.727696990598729e-08
+    1.513564934452811e-07
+     4.10469518412313e-07
+ 9.2e+09     
+    4.100891082442404e-07
+    1.513697115319492e-07
+     4.07227721462982e-07
+     4.73338114114488e-08
+    9.421801468849313e-08
+    4.071636156218046e-07
+    2.658867524268917e-08
+     4.73314691025551e-08
+    1.514147669748672e-07
+     4.10522931610233e-07
+ 9.3e+09     
+    4.101430933808543e-07
+    1.514285767204626e-07
+    4.072810689787121e-07
+    4.738903859283559e-08
+    9.427599034947253e-08
+     4.07216991061907e-07
+    2.664044312986479e-08
+    4.738666686044352e-08
+    1.514736190907311e-07
+    4.105771536318505e-07
+ 9.4e+09     
+    4.101978942337303e-07
+    1.514880183187103e-07
+    4.073352279958921e-07
+    4.744496654968938e-08
+    9.433484406602834e-08
+    4.072711744334215e-07
+    2.669287264930924e-08
+    4.744256512255053e-08
+    1.515330384429035e-07
+    4.106321777167819e-07
+ 9.5e+09     
+    4.102535045849873e-07
+    1.515480254638849e-07
+    4.073901935738925e-07
+    4.750159687421887e-08
+    9.439458188063533e-08
+     4.07326160627923e-07
+    2.674596888829862e-08
+    4.749916572242081e-08
+     1.51593013796491e-07
+     4.10687997374834e-07
+ 9.6e+09     
+    4.103099184501171e-07
+    1.516085873385941e-07
+    4.074459608235262e-07
+    4.755893098784073e-08
+    9.445520885516762e-08
+    4.073819446112703e-07
+    2.679973714923369e-08
+    4.755647039263771e-08
+     1.51653534052083e-07
+    4.107446063807157e-07
+ 9.7e+09     
+    4.103671300691307e-07
+    1.516696931795363e-07
+    4.075025249131852e-07
+    4.761697013923001e-08
+    9.451672915387491e-08
+    4.074385214329989e-07
+    2.685418294366326e-08
+    4.761448077117688e-08
+    1.517145882669084e-07
+    4.108019987694732e-07
+ 9.8e+09     
+    4.104251338981197e-07
+    1.517313322861386e-07
+    4.075598810750708e-07
+    4.767571539919664e-08
+     9.45791461235002e-08
+    4.074958862359905e-07
+    2.690931198481371e-08
+    4.767319840505739e-08
+    1.517761656766153e-07
+    4.108601688325455e-07
+ 9.9e+09     
+     4.10483924601133e-07
+    1.517934940290589e-07
+    4.076180246112553e-07
+    4.773516765179519e-08
+    9.464246236920626e-08
+    4.075540342661486e-07
+    2.696513017841787e-08
+    4.773262475067459e-08
+    1.518382557175707e-07
+    4.109191111143805e-07
+ 1e+10       
+    4.105434970423134e-07
+    1.518561678584655e-07
+     4.07676950899373e-07
+    4.779532758111034e-08
+    9.470667982541157e-08
+    4.076129608818726e-07
+    2.702164361163332e-08
+    4.779276117022086e-08
+    1.519008480495785e-07
+     4.10978820409516e-07
+ 1.01e+10    
+    4.106110951656923e-07
+    1.519273025342471e-07
+    4.077549430048369e-07
+    4.785504308961082e-08
+    9.478647380220445e-08
+    4.076894347023091e-07
+    2.707573417174863e-08
+    4.785252242357304e-08
+        1.51971843142e-07
+    4.110465546055068e-07
+ 1.02e+10    
+    4.106787611991297e-07
+     1.51998319024758e-07
+    4.078322145698181e-07
+    4.791475399024049e-08
+    9.486546491378036e-08
+    4.077652949660089e-07
+     2.71298770855387e-08
+    4.791227568855205e-08
+    1.520427311604616e-07
+    4.111143566890004e-07
+ 1.03e+10    
+    4.107464926548918e-07
+    1.520692181781614e-07
+    4.079087915544738e-07
+    4.797445785520439e-08
+    9.494367977721384e-08
+    4.078405619198404e-07
+    2.718406592895193e-08
+    4.797201871873149e-08
+    1.521135123511141e-07
+    4.111822241444833e-07
+ 1.04e+10    
+    4.108142872161003e-07
+      1.5214000090289e-07
+    4.079846990766903e-07
+     4.80341522382307e-08
+    9.502114407999798e-08
+     4.07915255258691e-07
+    2.723829438747056e-08
+    4.803174924042631e-08
+    1.521841870516791e-07
+    4.112501546274875e-07
+ 1.05e+10    
+    4.108821427304378e-07
+    1.522106681646535e-07
+    4.080599614399694e-07
+    4.809383467817815e-08
+    9.509788261342445e-08
+    4.079893941384538e-07
+    2.729255625513876e-08
+    4.809146495674674e-08
+    1.522547556868204e-07
+    4.113181459583081e-07
+ 1.06e+10    
+    4.109500572040014e-07
+    1.522812209835173e-07
+    4.081346021604056e-07
+    4.815350270247947e-08
+    9.517391930485482e-08
+    4.080629971888928e-07
+    2.734684543356304e-08
+    4.815116355146551e-08
+    1.523252187636778e-07
+    4.113861961158774e-07
+ 1.07e+10    
+    4.110180287953074e-07
+    1.523516604310547e-07
+    4.082086439927822e-07
+    4.821315383042827e-08
+    9.524927724890638e-08
+    4.081360825263801e-07
+    2.740115593088803e-08
+    4.821084269270493e-08
+    1.523955768675544e-07
+    4.114543032317781e-07
+ 1.08e+10    
+    4.110860558094445e-07
+    1.524219876275756e-07
+     4.08282108955817e-07
+    4.827278557631001e-08
+    9.532397873757535e-08
+    4.082086677664845e-07
+    2.745548186074946e-08
+    4.827050003644675e-08
+    1.524658306577602e-07
+    4.115224655844161e-07
+ 1.09e+10    
+    4.111541366923815e-07
+    1.524922037394308e-07
+    4.083550183565772e-07
+    4.833239545238253e-08
+    9.539804528932146e-08
+    4.082807700364006e-07
+    2.750981744120685e-08
+    4.833013322987105e-08
+     1.52535980863606e-07
+    4.115906815933387e-07
+ 1.1e+10     
+    4.112222700254254e-07
+    1.525623099763978e-07
+    4.084273928141012e-07
+    4.839198097170756e-08
+     9.54714976771398e-08
+    4.083524059872037e-07
+    2.756415699365812e-08
+    4.838973991452914e-08
+    1.526060282805455e-07
+    4.116589498137091e-07
+ 1.11e+10    
+    4.112904545198304e-07
+     1.52632307589143e-07
+    4.084992522822392e-07
+    4.845153965084109e-08
+    9.554435595564644e-08
+    4.084235918059295e-07
+    2.761849494173803e-08
+    4.844931772935498e-08
+    1.526759737664626e-07
+    4.117272689309259e-07
+ 1.12e+10    
+    4.113586890115613e-07
+    1.527021978667647e-07
+    4.085706160717444e-07
+    4.851106901238323e-08
+    9.561663948720381e-08
+    4.084943432274587e-07
+    2.767282581020242e-08
+    4.850886431352023e-08
+    1.527458182381003e-07
+    4.117956377554021e-07
+ 1.13e+10    
+    4.114269724562029e-07
+    1.527719821344158e-07
+    4.086415028716358e-07
+    4.857056658739233e-08
+    9.568836696711341e-08
+     4.08564675546208e-07
+    2.772714422380007e-08
+    4.856837730913872e-08
+    1.528155626676286e-07
+    4.118640552174843e-07
+ 1.14e+10    
+    4.114953039240238e-07
+    1.528416617510058e-07
+    4.087119307698566e-07
+    4.863002991766933e-08
+    9.575955644790272e-08
+    4.086346036276199e-07
+    2.778144490613395e-08
+    4.862785436382382e-08
+    1.528852080793468e-07
+    4.119325203625282e-07
+ 1.15e+10    
+    4.115636825951822e-07
+    1.529112381069819e-07
+    4.087819172732503e-07
+     4.86894565579144e-08
+    9.583022536273372e-08
+    4.087041419194396e-07
+    2.783572267851358e-08
+    4.868729313310568e-08
+    1.529547555465174e-07
+    4.120010323461175e-07
+ 1.16e+10    
+    4.116321077550824e-07
+    1.529807126221874e-07
+    4.088514793268706e-07
+    4.874884407776012e-08
+    9.590039054795953e-08
+    4.087733044627861e-07
+    2.788997245879962e-08
+    4.874669128271093e-08
+    1.530242061883288e-07
+    4.120695904294292e-07
+ 1.17e+10    
+    4.117005787898727e-07
+    1.530500867437993e-07
+    4.089206333326555e-07
+    4.880819006368688e-08
+    9.597006826485728e-08
+    4.088421049030043e-07
+     2.79441892602428e-08
+    4.880604649071155e-08
+    1.530935611669814e-07
+    4.121381939747439e-07
+ 1.18e+10    
+      4.1176909518209e-07
+    1.531193619443411e-07
+    4.089893951674812e-07
+    4.886749212082298e-08
+    9.603927422056228e-08
+    4.089105565003015e-07
+    2.799836819031801e-08
+    4.886535644954684e-08
+    1.531628216848955e-07
+    4.122068424410949e-07
+ 1.19e+10    
+    4.118376565064383e-07
+    1.531885397197711e-07
+     4.09057780200609e-07
+    4.892674787463412e-08
+    9.610802358823098e-08
+     4.08978672140163e-07
+    2.805250444955519e-08
+    4.892461886792318e-08
+     1.53231988982036e-07
+    4.122755353800619e-07
+ 1.2e+10     
+    4.119062624257091e-07
+    1.532576215876447e-07
+    4.091258033105585e-07
+    4.898595497250548e-08
+    9.617633102645769e-08
+    4.090464643435501e-07
+     2.81065933303677e-08
+     4.89838314725953e-08
+    1.533010643333514e-07
+    4.123442724316948e-07
+ 1.21e+10    
+    4.119749126868364e-07
+     1.53326609085349e-07
+    4.091934789014098e-07
+    4.904511108522101e-08
+    9.624421069797039e-08
+    4.091139452768735e-07
+    2.816063021588009e-08
+    4.904299201003595e-08
+    1.533700490463225e-07
+    4.124130533205819e-07
+ 1.22e+10    
+    4.120436071170844e-07
+    1.533955037684086e-07
+    4.092608209185686e-07
+    4.910421390834488e-08
+    9.631167628763162e-08
+    4.091811267617487e-07
+    2.821461057875569e-08
+    4.910209824799546e-08
+    1.534389444586176e-07
+    4.124818778520379e-07
+ 1.23e+10    
+    4.121123456203644e-07
+    1.534643072088606e-07
+    4.093278428639982e-07
+    4.916326116350451e-08
+    9.637874101976683e-08
+    4.092480202845309e-07
+    2.826852998002492e-08
+    4.916114797695653e-08
+    1.535077519358525e-07
+     4.12550745908435e-07
+ 1.24e+10    
+    4.121811281736798e-07
+    1.535330209936973e-07
+    4.093945578109426e-07
+    4.922225059958522e-08
+    9.644541767484521e-08
+    4.093146370056269e-07
+    2.832238406791593e-08
+    4.922013901148938e-08
+    1.535764728694467e-07
+    4.126196574456463e-07
+ 1.25e+10    
+    4.122499548236938e-07
+    1.536016467233747e-07
+    4.094609784181564e-07
+    4.928117999383324e-08
+    9.651171860553548e-08
+    4.093809877685945e-07
+     2.83761685766877e-08
+     4.92790691915102e-08
+    1.536451086745804e-07
+     4.12688612489628e-07
+ 1.26e+10    
+    4.123188256834226e-07
+    1.536701860103857e-07
+    4.095271169436572e-07
+    4.934004715287758e-08
+    9.657765575215976e-08
+    4.094470831090203e-07
+    2.842987932546677e-08
+    4.933793638344646e-08
+    1.537136607882406e-07
+    4.127576111331096e-07
+ 1.27e+10    
+     4.12387740929041e-07
+    1.537386404778948e-07
+    4.095929852580155e-07
+    4.939884991366676e-08
+    9.664324065756586e-08
+    4.095129332631846e-07
+    2.848351221708814e-08
+     4.93967384813141e-08
+    1.537821306673585e-07
+    4.128266535324099e-07
+ 1.28e+10    
+    4.124567007968108e-07
+    1.538070117584344e-07
+    4.096585948571951e-07
+    4.945758614433036e-08
+    9.670848448144121e-08
+    4.095785481765157e-07
+    2.853706323694113e-08
+    4.945547340770957e-08
+    1.538505197870334e-07
+    4.128957399043655e-07
+ 1.29e+10    
+    4.125257055801161e-07
+    1.538753014926592e-07
+    4.097239568749673e-07
+    4.951625374496443e-08
+    9.677339801408703e-08
+    4.096439375118301e-07
+    2.859052845182084e-08
+    4.951413911471972e-08
+     1.53918829638839e-07
+    4.129648705233728e-07
+ 1.3e+10     
+    4.125947556266106e-07
+    1.539435113281575e-07
+    4.097890820949004e-07
+    4.957485064834492e-08
+    9.683799168967424e-08
+    4.097091106573712e-07
+    2.864390400878551e-08
+    4.957273358475467e-08
+      1.5398706172921e-07
+    4.130340457185366e-07
+ 1.31e+10    
+    4.126638513354727e-07
+    1.540116429183181e-07
+    4.098539809619487e-07
+    4.963337482057365e-08
+    9.690227559899935e-08
+    4.097740767346374e-07
+    2.869718613402086e-08
+    4.963125483130555e-08
+    1.540552175779054e-07
+    4.131032658709279e-07
+ 1.32e+10    
+    4.127329931547609e-07
+    1.540796979212493e-07
+    4.099186635936508e-07
+    4.969182426165731e-08
+    9.696625950175915e-08
+     4.09838844606014e-07
+    2.875037113171112e-08
+     4.96897008996307e-08
+    1.541232987165465e-07
+    4.131725314109414e-07
+ 1.33e+10    
+    4.128021815788749e-07
+    1.541476779987512e-07
+    4.099831397909484e-07
+    4.975019700602414e-08
+    9.702995283836349e-08
+    4.099034228822034e-07
+    2.880345538291806e-08
+    4.974806986737462e-08
+    1.541913066872252e-07
+    4.132418428157597e-07
+ 1.34e+10    
+    4.128714171461087e-07
+    1.542155848153354e-07
+    4.100474190486395e-07
+     4.98084911229808e-08
+    9.709336474130095e-08
+    4.099678199294632e-07
+    2.885643534446751e-08
+    4.980635984511996e-08
+    1.542592430411809e-07
+    4.133112006069064e-07
+ 1.35e+10    
+    4.129407004363057e-07
+    1.542834200372947e-07
+    4.101115105654819e-07
+    4.986670471711166e-08
+    9.715650404607773e-08
+    4.100320438766505e-07
+    2.890930754784463e-08
+    4.986456897687947e-08
+    1.543271093375429e-07
+    4.133806053479002e-07
+ 1.36e+10    
+    4.130100320685974e-07
+    1.543511853318175e-07
+    4.101754232539531e-07
+    4.992483592862266e-08
+    9.721937930174271e-08
+    4.100961026220791e-07
+    2.896206859809745e-08
+    4.992269544052705e-08
+    1.543949071421354e-07
+    4.134500576419976e-07
+ 1.37e+10    
+    4.130794126992398e-07
+    1.544188823661466e-07
+    4.102391657496784e-07
+    4.998288293363436e-08
+    9.728199878101682e-08
+    4.101600038401947e-07
+    2.901471517274954e-08
+    4.998073744817323e-08
+    1.544626380263431e-07
+    4.135195581300273e-07
+ 1.38e+10    
+    4.131488430195282e-07
+    1.544865128067818e-07
+    4.103027464205456e-07
+    5.004084394442387e-08
+    9.734437049004026e-08
+    4.102237549880639e-07
+    2.906724402072179e-08
+     5.00386932464856e-08
+     1.54530303566034e-07
+    4.135891074883043e-07
+ 1.39e+10    
+    4.132183237538037e-07
+    1.545540783187226e-07
+    4.103661733755058e-07
+     5.00987172096201e-08
+    9.740650217775349e-08
+    4.102873633116912e-07
+    2.911965196126379e-08
+     5.00965611169597e-08
+    1.545979053405382e-07
+    4.136587064266343e-07
+ 1.4e+10     
+    4.132878556575329e-07
+    1.546215805647505e-07
+    4.104294544730818e-07
+    5.015650101435373e-08
+    9.746840134492482e-08
+    4.103508358521598e-07
+    2.917193588289457e-08
+    5.015433937613928e-08
+    1.546654449316788e-07
+    4.137283556863962e-07
+ 1.41e+10    
+    4.133574395154705e-07
+    1.546890212047495e-07
+    4.104925973295854e-07
+    5.021419368036398e-08
+    9.753007525283892e-08
+    4.104141794516043e-07
+     2.92240927423533e-08
+    5.021202637579106e-08
+    1.547329239228544e-07
+     4.13798056038699e-07
+ 1.42e+10    
+    4.134270761398974e-07
+    1.547564018950632e-07
+    4.105556093270604e-07
+    5.027179356606507e-08
+    9.759153093165967e-08
+    4.104774007590154e-07
+    2.927611956356011e-08
+    5.026962050303557e-08
+     1.54800343898169e-07
+    4.138678082826209e-07
+ 1.43e+10    
+    4.134967663689298e-07
+    1.548237242878852e-07
+    4.106184976209505e-07
+     5.03292990665735e-08
+    9.765277518847804e-08
+    4.105405062358841e-07
+    2.932801343658675e-08
+    5.032712018043507e-08
+    1.548677064416092e-07
+    4.139376132435123e-07
+ 1.44e+10    
+    4.135665110648993e-07
+    1.548909900306854e-07
+    4.106812691475186e-07
+    5.038670861369879e-08
+    9.771381461506017e-08
+    4.106035021616852e-07
+    2.937977151663773e-08
+     5.03845238660432e-08
+    1.549350131362651e-07
+     4.14007471771379e-07
+ 1.45e+10    
+    4.136363111128021e-07
+    1.549582007656655e-07
+    4.107439306310038e-07
+    5.044402067589966e-08
+    9.777465559530416e-08
+    4.106663946392082e-07
+    2.943139102304166e-08
+    5.044183005341569e-08
+    1.550022655635937e-07
+    4.140773847393234e-07
+ 1.46e+10    
+    4.137061674188149e-07
+     1.55025358129248e-07
+    4.108064885905456e-07
+    5.050123375820654e-08
+    9.783530431241866e-08
+    4.107291895997357e-07
+    2.948286923825311e-08
+    5.049903727158555e-08
+    1.550694653027228e-07
+    4.141473530420598e-07
+ 1.47e+10    
+    4.137760809088698e-07
+     1.55092463751592e-07
+    4.108689493468706e-07
+    5.055834640211324e-08
+    9.789576675583413e-08
+    4.107918928080737e-07
+    2.953420350686476e-08
+    5.055614408500585e-08
+     1.55136613929793e-07
+    4.142173775944844e-07
+ 1.48e+10    
+    4.138460525272946e-07
+    1.551595192561382e-07
+    4.109313190287527e-07
+    5.061535718543997e-08
+    9.795604872785545e-08
+    4.108545098674377e-07
+    2.958539123463043e-08
+    5.061314909345833e-08
+    1.552037130173375e-07
+    4.142874593303145e-07
+ 1.49e+10    
+     4.13916083235511e-07
+    1.552265262591812e-07
+    4.109936035792572e-07
+    5.067226472216627e-08
+    9.801615585006787e-08
+    4.109170462242011e-07
+    2.963642988749828e-08
+    5.067005093193381e-08
+    1.552707641336962e-07
+    4.143575992007797e-07
+ 1.5e+10     
+    4.139861740107873e-07
+     1.55293486369466e-07
+    4.110558087617729e-07
+    5.072906766224067e-08
+    9.807609356950466e-08
+    4.109795071725012e-07
+    2.968731699065496e-08
+    5.072684827048309e-08
+    1.553377688424632e-07
+    4.144277981733728e-07
+ 1.51e+10    
+    4.140563258450495e-07
+    1.553604011878101e-07
+    4.111179401658407e-07
+    5.078576469136312e-08
+    9.813586716458587e-08
+     4.11041897858717e-07
+    2.973805012758015e-08
+     5.07835398140415e-08
+     1.55404728701967e-07
+    4.144980572306546e-07
+ 1.52e+10    
+    4.141265397437405e-07
+    1.554272723067483e-07
+    4.111800032127886e-07
+    5.084235453074532e-08
+    9.819548175083749e-08
+    4.111042232858148e-07
+    2.978862693911184e-08
+    5.084012430222802e-08
+    1.554716452647807e-07
+    4.145683773691112e-07
+ 1.53e+10    
+    4.141968167247345e-07
+    1.554941013102001e-07
+    4.112420031611715e-07
+    5.089883593684948e-08
+    9.825494228639893e-08
+     4.11166488317566e-07
+    2.983904512252221e-08
+    5.089660050912103e-08
+    1.555385200772609e-07
+    4.146387595980596e-07
+ 1.54e+10    
+    4.142671578172954e-07
+    1.555608897731583e-07
+    4.113039451120333e-07
+    5.095520770110553e-08
+    9.831425357732749e-08
+     4.11228697682643e-07
+     2.98893024306039e-08
+    5.095296724301072e-08
+    1.556053546791151e-07
+    4.147092049386058e-07
+ 1.55e+10    
+    4.143375640610857e-07
+     1.55627639261397e-07
+    4.113658340139874e-07
+    5.101146864961034e-08
+    9.837342028270739e-08
+    4.112908559785955e-07
+    2.993939667076725e-08
+    5.100922334613257e-08
+    1.556721506029944e-07
+    4.147797144226453e-07
+ 1.56e+10    
+    4.144080365052198e-07
+    1.556943513312007e-07
+    4.114276746681306e-07
+    5.106761764280799e-08
+    9.843244691957094e-08
+    4.113529676757058e-07
+    2.998932570414765e-08
+    5.106536769437944e-08
+    1.557389093741117e-07
+    4.148502890919118e-07
+ 1.57e+10    
+    4.144785762073579e-07
+    1.557610275291095e-07
+     4.11489471732788e-07
+     5.11236535751544e-08
+    9.849133786763919e-08
+    4.114150371207367e-07
+     3.00390874447237e-08
+    5.112139919699603e-08
+    1.558056325098845e-07
+    4.149209299970677e-07
+ 1.58e+10    
+    4.145491842328449e-07
+     1.55827669391684e-07
+    4.115512297281003e-07
+    5.117957537476545e-08
+    9.855009737388955e-08
+    4.114770685405652e-07
+    3.008867985844575e-08
+     5.11773167962573e-08
+    1.558723215195986e-07
+    4.149916381968341e-07
+ 1.59e+10    
+    4.146198616538863e-07
+    1.558942784452847e-07
+    4.116129530404573e-07
+    5.123538200305096e-08
+    9.860872955695551e-08
+    4.115390660457073e-07
+     3.01381009623746e-08
+    5.123311946712928e-08
+    1.559389779040951e-07
+     4.15062414757165e-07
+ 1.6e+10     
+    4.146906095487654e-07
+    1.559608562058688e-07
+    4.116746459267817e-07
+    5.129107245433582e-08
+    9.866723841136655e-08
+     4.11601033633738e-07
+    3.018734882383103e-08
+    5.128880621691675e-08
+     1.56005603155477e-07
+    4.151332607504545e-07
+ 1.61e+10    
+    4.147614290010948e-07
+    1.560274041788018e-07
+    4.117363125186704e-07
+    5.134664575546793e-08
+    9.872562781163431e-08
+    4.116629751926164e-07
+    3.023642155955511e-08
+    5.134437608489648e-08
+    1.560721987568353e-07
+    4.152041772547855e-07
+ 1.62e+10    
+    4.148323210991033e-07
+    1.560939238586826e-07
+    4.117979568263967e-07
+    5.140210096541518e-08
+    9.878390151618935e-08
+    4.117248945039013e-07
+    3.028531733487614e-08
+    5.139982814193815e-08
+    1.561387661819945e-07
+     4.15275165353211e-07
+ 1.63e+10    
+    4.149032869349586e-07
+    1.561604167291828e-07
+    4.118595827427758e-07
+    5.145743717485189e-08
+    9.884206317117592e-08
+    4.117867952458785e-07
+    3.033403436289246e-08
+    5.145516149011374e-08
+     1.56205306895274e-07
+     4.15346226133069e-07
+ 1.64e+10    
+    4.149743276041218e-07
+    1.562268842628994e-07
+    4.119211940469083e-07
+    5.151265350573619e-08
+    9.890011631410994e-08
+    4.118486809965915e-07
+    3.038257090366162e-08
+    5.151037526229605e-08
+     1.56271822351268e-07
+    4.154173606853306e-07
+ 1.65e+10    
+    4.150454442047321e-07
+    1.562933279212185e-07
+    4.119827944077882e-07
+    5.156774911087768e-08
+    9.895806437740425e-08
+    4.119105552367819e-07
+    3.043092526340029e-08
+     5.15654686217478e-08
+    1.563383139946403e-07
+    4.154885701039807e-07
+ 1.66e+10    
+    4.151166378370214e-07
+    1.563597491541918e-07
+    4.120443873878005e-07
+    5.162272317349801e-08
+    9.901591069176787e-08
+    4.119724213527426e-07
+    3.047909579369426e-08
+    5.162044076170166e-08
+    1.564047832599346e-07
+    4.155598554854246e-07
+ 1.67e+10    
+    4.151879096027588e-07
+    1.564261494004233e-07
+    4.121059764460945e-07
+    5.167757490678421e-08
+    9.907365848948276e-08
+    4.120342826390814e-07
+    3.052708089071835e-08
+    5.167529090493263e-08
+    1.564712315713985e-07
+    4.156312179279277e-07
+ 1.68e+10    
+    4.152592606047222e-07
+    1.564925300869681e-07
+    4.121675649418508e-07
+    5.173230355343565e-08
+     9.91313109075639e-08
+    4.120961423014085e-07
+    3.057487899446607e-08
+    5.173001830332263e-08
+    1.565376603428219e-07
+    4.157026585310803e-07
+ 1.69e+10    
+    4.153306919461958e-07
+    1.565588926292378e-07
+    4.122291561374322e-07
+     5.17869083852052e-08
+     9.91888709908056e-08
+    4.121580034589367e-07
+    3.062248858798887e-08
+    5.178462223741907e-08
+    1.566040709773877e-07
+    4.157741783952879e-07
+ 1.7e+10     
+    4.154022047304921e-07
+    1.566252384309199e-07
+    4.122907532014381e-07
+    5.184138870243532e-08
+    9.924634169472028e-08
+    4.122198691470047e-07
+    3.066990819664508e-08
+    5.183910201598739e-08
+    1.566704648675343e-07
+    4.158457786212881e-07
+ 1.71e+10    
+    4.154738000605006e-07
+    1.566915688839017e-07
+    4.123523592116505e-07
+    5.189574383359066e-08
+    9.930372588837261e-08
+    4.122817423195285e-07
+    3.071713638735858e-08
+    5.189345697555895e-08
+    1.567368433948321e-07
+    4.159174603096933e-07
+ 1.72e+10    
+    4.155454790382563e-07
+    1.567578853682061e-07
+    4.124139771578861e-07
+    5.194997313478616e-08
+    9.936102635711266e-08
+    4.123436258513714e-07
+    3.076417176788656e-08
+    5.194768647997399e-08
+    1.568032079298668e-07
+    4.159892245605509e-07
+ 1.73e+10    
+    4.156172427645337e-07
+    1.568241892519333e-07
+    4.124756099447521e-07
+    5.200407598931192e-08
+    9.941824580521347e-08
+    4.124055225406503e-07
+    3.081101298609704e-08
+    5.200178991992152e-08
+    1.568695598321372e-07
+    4.160610724729335e-07
+ 1.74e+10    
+     4.15689092338459e-07
+    1.568904818912111e-07
+    4.125372603943106e-07
+    5.205805180715669e-08
+    9.947538685841485e-08
+    4.124674351109658e-07
+    3.085765872925536e-08
+    5.205576671247504e-08
+    1.569359004499603e-07
+     4.16133005144542e-07
+ 1.75e+10    
+    4.157610288571432e-07
+    1.569567646301517e-07
+    4.125989312486569e-07
+    5.211190002452813e-08
+    9.953245206637811e-08
+    4.125293662135679e-07
+    3.090410772332001e-08
+    5.210961630062669e-08
+    1.570022311203872e-07
+    4.162050236713368e-07
+ 1.76e+10    
+    4.158330534153378e-07
+    1.570230388008162e-07
+    4.126606251724079e-07
+    5.216562010337198e-08
+    9.958944390505479e-08
+    4.125913184294559e-07
+    3.095035873224768e-08
+    5.216333815281877e-08
+    1.570685531691265e-07
+    4.162771291471821e-07
+ 1.77e+10    
+    4.159051671051037e-07
+    1.570893057231846e-07
+    4.127223447551137e-07
+    5.221921153089089e-08
+    9.964636477897271e-08
+    4.126532942714153e-07
+    3.099641055730705e-08
+    5.221693176247368e-08
+    1.571348679104776e-07
+    4.163493226635125e-07
+ 1.78e+10    
+    4.159773710155039e-07
+    1.571555667051325e-07
+    4.127840925135855e-07
+    5.227267381906158e-08
+     9.97032170234421e-08
+    4.127152961859909e-07
+    3.104226203640189e-08
+    5.227039664752308e-08
+    1.572011766472708e-07
+    4.164216053090162e-07
+ 1.79e+10    
+     4.16049666232306e-07
+    1.572218230424137e-07
+    4.128458708941493e-07
+    5.232600650415284e-08
+      9.9760002906685e-08
+    4.127773265554015e-07
+    3.108791204340269e-08
+    5.232373234993618e-08
+    1.572674806708151e-07
+    4.164939781693344e-07
+ 1.8e+10     
+     4.16122053837709e-07
+    1.572880760186475e-07
+    4.129076822748242e-07
+    5.237920914624333e-08
+    9.981672463189152e-08
+    4.128393876993967e-07
+    3.113335948748736e-08
+    5.237693843524825e-08
+    1.573337812608539e-07
+    4.165664423267807e-07
+ 1.81e+10    
+    4.161945349100777e-07
+    1.573543269053112e-07
+    4.129695289674274e-07
+     5.24322813287405e-08
+    9.987338433920424e-08
+    4.129014818770572e-07
+     3.11786033124903e-08
+    5.243001449208862e-08
+    1.574000796855261e-07
+    4.166389988600685e-07
+ 1.82e+10    
+    4.162671105236994e-07
+    1.574205769617387e-07
+    4.130314132196147e-07
+    5.248522265789981e-08
+    9.992998410763486e-08
+    4.129636112885389e-07
+    3.122364249626034e-08
+    5.248296013171022e-08
+     1.57466377201335e-07
+     4.16711648844063e-07
+ 1.83e+10    
+    4.163397817485478e-07
+    1.574868274351221e-07
+     4.13093337216847e-07
+    5.253803276234651e-08
+    9.998652595691467e-08
+    4.130257780767686e-07
+    3.126847605002714e-08
+    5.253577498751956e-08
+    1.575326750531221e-07
+    4.167843933495383e-07
+ 1.84e+10    
+    4.164125496500659e-07
+    1.575530795605183e-07
+    4.131553030843017e-07
+    5.259071129259795e-08
+    1.000430118492821e-07
+    4.130879843290806e-07
+    3.131310301777587e-08
+    5.258845871460813e-08
+     1.57598974474047e-07
+    4.168572334429549e-07
+ 1.85e+10    
+    4.164854152889584e-07
+    1.576193345608601e-07
+    4.132173128887092e-07
+    5.264325792058921e-08
+    1.000994436912087e-07
+    4.131502320788127e-07
+    3.135752247563057e-08
+    5.264101098928603e-08
+    1.576652766855731e-07
+    4.169301701862464e-07
+ 1.86e+10    
+    4.165583797210001e-07
+    1.576855936469704e-07
+    4.132793686401442e-07
+    5.269567233920024e-08
+    1.001558233350669e-07
+    4.132125233068459e-07
+    3.140173353124542e-08
+    5.269343150861649e-08
+    1.577315828974573e-07
+    4.170032046366189e-07
+ 1.87e+10    
+    4.166314439968489e-07
+    1.577518580175802e-07
+    4.133414722937424e-07
+    5.274795426178541e-08
+     1.00212152580741e-07
+     4.13274859943103e-07
+    3.144573532320439e-08
+    5.274571998995389e-08
+    1.577978943077461e-07
+    4.170763378463652e-07
+ 1.88e+10    
+    4.167046091618797e-07
+    1.578181288593502e-07
+    4.134036257513759e-07
+      5.2800103421707e-08
+    1.002684331771836e-07
+     4.13337243867997e-07
+    3.148952702042899e-08
+    5.279787617048369e-08
+     1.57864212102774e-07
+    4.171495708626853e-07
+ 1.89e+10    
+    4.167778762560224e-07
+    1.578844073468959e-07
+     4.13465830863262e-07
+    5.285211957187119e-08
+    1.003246668239197e-07
+    4.133996769138414e-07
+    3.153310782159417e-08
+    5.284989980676536e-08
+     1.57930537457169e-07
+    4.172229047275229e-07
+ 1.9e+10     
+    4.168512463136104e-07
+    1.579506946428152e-07
+      4.1352808942953e-07
+    5.290400248426711e-08
+    1.003808551725008e-07
+    4.134621608662108e-07
+    3.157647695455176e-08
+    5.290179067427834e-08
+    1.579968715338595e-07
+    4.172963404774081e-07
+ 1.91e+10    
+    4.169247203632423e-07
+    1.580169918977184e-07
+    4.135904032017264e-07
+    5.295575194951035e-08
+     1.00436999827909e-07
+    4.135246974652666e-07
+    3.161963367576228e-08
+    5.295354856697134e-08
+    1.580632154840865e-07
+    4.173698791433134e-07
+ 1.92e+10    
+    4.169982994276507e-07
+    1.580833002502625e-07
+    4.136527738842816e-07
+    5.300736777638937e-08
+    1.004931023499156e-07
+    4.135872884070378e-07
+    3.166257726973425e-08
+    5.300517329681532e-08
+    1.581295704474191e-07
+    4.174435217505148e-07
+ 1.93e+10    
+    4.170719845235793e-07
+    1.581496208271866e-07
+    4.137152031359211e-07
+    5.305884979141677e-08
+    1.005491642543942e-07
+    4.136499353446667e-07
+    3.170530704847124e-08
+    5.305666469335993e-08
+    1.581959375517734e-07
+    4.175172693184675e-07
+ 1.94e+10    
+      4.1714577666167e-07
+    1.582159547433493e-07
+    4.137776925710344e-07
+    5.311019783838371e-08
+    1.006051870145894e-07
+    4.137126398896137e-07
+    3.174782235092661e-08
+    5.310802260329391e-08
+    1.582623179134343e-07
+    4.175911228606846e-07
+ 1.95e+10    
+    4.172196768463577e-07
+    1.582823031017706e-07
+    4.138402437610019e-07
+    5.316141177791958e-08
+     1.00661172062345e-07
+     4.13775403612828e-07
+    3.179012254246591e-08
+    5.315924689000993e-08
+    1.583287126370808e-07
+    4.176650833846279e-07
+ 1.96e+10    
+    4.172936860757706e-07
+    1.583486669936731e-07
+     4.13902858235472e-07
+    5.321249148705561e-08
+    1.007171207892909e-07
+    4.138382280458811e-07
+     3.18322070143364e-08
+    5.321033743317303e-08
+    1.583951228158134e-07
+    4.177391518916034e-07
+ 1.97e+10    
+    4.173678053416442e-07
+    1.584150474985271e-07
+    4.139655374836047e-07
+     5.32634368587934e-08
+    1.007730345479911e-07
+    4.139011146820679e-07
+    3.187407518314452e-08
+    5.326129412829422e-08
+    1.584615495311852e-07
+    4.178133293766674e-07
+ 1.98e+10    
+    4.174420356292325e-07
+    1.584814456840968e-07
+    4.140282829552703e-07
+    5.331424780167748e-08
+    1.008289146530545e-07
+    4.139640649774738e-07
+    3.191572649034019e-08
+    5.331211688630788e-08
+     1.58527993853235e-07
+    4.178876168285385e-07
+ 1.99e+10    
+     4.17516377917234e-07
+    1.585478626064875e-07
+    4.140910960622099e-07
+    5.336492423937398e-08
+    1.008847623822094e-07
+     4.14027080352007e-07
+    3.195716040170866e-08
+    5.336280563315417e-08
+    1.585944568405216e-07
+    4.179620152295124e-07
+ 2e+10       
+    4.175908331777218e-07
+    1.586142993101965e-07
+    4.141539781791618e-07
+    5.341546611025287e-08
+    1.009405789773435e-07
+    4.140901621904053e-07
+     3.19983764068695e-08
+    5.341336030936657e-08
+    1.586609395401631e-07
+    4.180365255553917e-07
+ 2.01e+10    
+    4.176654023760778e-07
+    1.586807568281629e-07
+    4.142169306449481e-07
+    5.346587336697636e-08
+    1.009963656455095e-07
+     4.14153311843207e-07
+    3.203937401878259e-08
+    5.346378086966345e-08
+    1.587274429878754e-07
+    4.181111487754123e-07
+ 2.02e+10    
+    4.177400864709345e-07
+    1.587472361818211e-07
+    4.142799547635274e-07
+    5.351614597609179e-08
+    1.010521235598987e-07
+    4.142165306276953e-07
+    3.208015277326139e-08
+    5.351406728254537e-08
+    1.587939682080146e-07
+    4.181858858521836e-07
+ 2.03e+10    
+    4.178148864141229e-07
+    1.588137383811537e-07
+    4.143430518050161e-07
+     5.35662839176299e-08
+     1.01107853860784e-07
+    4.142798198288142e-07
+    3.212071222849287e-08
+      5.3564219529897e-08
+    1.588605162136198e-07
+    4.182607377416276e-07
+ 2.04e+10    
+    4.178898031506219e-07
+     1.58880264424747e-07
+    4.144062230066736e-07
+    5.361628718470859e-08
+    1.011635576564321e-07
+    4.143431807000563e-07
+    3.216105196456458e-08
+    5.361423760659464e-08
+    1.589270880064592e-07
+    4.183357053929283e-07
+ 2.05e+10    
+     4.17964837618518e-07
+    1.589468152998471e-07
+    4.144694695738582e-07
+    5.366615578314179e-08
+    1.012192360239859e-07
+    4.144066144643229e-07
+    3.220117158299853e-08
+    5.366412152011826e-08
+    1.589936845770763e-07
+    4.184107897484847e-07
+ 2.06e+10    
+    4.180399907489652e-07
+    1.590133919824169e-07
+     4.14532792680952e-07
+    5.371588973105386e-08
+    1.012748900103213e-07
+    4.144701223147623e-07
+    3.224107070629166e-08
+     5.37138712901695e-08
+     1.59060306904839e-07
+    4.184859917438663e-07
+ 2.07e+10    
+    4.181152634661532e-07
+    1.590799954371943e-07
+    4.145961934722572e-07
+    5.376548905849945e-08
+    1.013305206328745e-07
+    4.145337054155771e-07
+    3.228074897746321e-08
+    5.376348694829468e-08
+    1.591269559579886e-07
+    4.185613123077759e-07
+ 2.08e+10    
+    4.181906566872743e-07
+    1.591466266177511e-07
+    4.146596730628627e-07
+    5.381495380708885e-08
+    1.013861288804441e-07
+    4.145973649028119e-07
+    3.232020605960865e-08
+    5.381296853751314e-08
+    1.591936326936917e-07
+    4.186367523620175e-07
+ 2.09e+10    
+    4.182661713225018e-07
+    1.592132864665539e-07
+    4.147232325394836e-07
+    5.386428402961878e-08
+    1.014417157139687e-07
+    4.146611018851161e-07
+    3.235944163546002e-08
+     5.38623161119511e-08
+    1.592603380580918e-07
+    4.187123128214632e-07
+ 2.1e+10     
+    4.183418082749658e-07
+    1.592799759150229e-07
+    4.147868729612724e-07
+    5.391347978970916e-08
+    1.014972820672793e-07
+    4.147249174444817e-07
+    3.239845540695308e-08
+    5.391152973648108e-08
+    1.593270729863637e-07
+      4.1878799459403e-07
+ 2.11e+10    
+    4.184175684407356e-07
+    1.593466958835951e-07
+    4.148505953606105e-07
+    5.396254116144469e-08
+    1.015528288478292e-07
+    4.147888126369643e-07
+    3.243724709480047e-08
+    5.396060948636649e-08
+    1.593938384027675e-07
+    4.188637985806579e-07
+ 2.12e+10    
+    4.184934527088057e-07
+    1.594134472817852e-07
+    4.149144007438666e-07
+    5.401146822902286e-08
+    1.016083569374002e-07
+    4.148527884933759e-07
+    3.247581643807166e-08
+    5.400955544691212e-08
+    1.594606352207045e-07
+    4.189397256752901e-07
+ 2.13e+10    
+    4.185694619610843e-07
+    1.594802310082494e-07
+    4.149782900921374e-07
+    5.406026108640742e-08
+    1.016638671927883e-07
+    4.149168460199637e-07
+    3.251416319377889e-08
+    5.405836771311979e-08
+    1.595274643427738e-07
+    4.190157767648583e-07
+ 2.14e+10    
+    4.186455970723847e-07
+    1.595470479508469e-07
+    4.150422643619611e-07
+    5.410891983698647e-08
+    1.017193604464669e-07
+    4.149809861990626e-07
+    3.255228713646934e-08
+    5.410704638934976e-08
+    1.595943266608295e-07
+    4.190919527292714e-07
+ 2.15e+10    
+    4.187218589104205e-07
+    1.596138989867055e-07
+    4.151063244860115e-07
+    5.415744459323796e-08
+    1.017748375072314e-07
+    4.150452099897337e-07
+    3.259018805782378e-08
+    5.415559158898753e-08
+    1.596612230560392e-07
+    4.191682544414072e-07
+ 2.16e+10    
+    4.187982483358026e-07
+    1.596807849822845e-07
+    4.151704713737688e-07
+    5.420583547639934e-08
+    1.018302991608228e-07
+    4.151095183283792e-07
+    3.262786576626089e-08
+    5.420400343411645e-08
+    1.597281543989426e-07
+    4.192446827671041e-07
+ 2.17e+10    
+    4.188747662020405e-07
+    1.597477067934399e-07
+    4.152347059121686e-07
+    5.425409261614339e-08
+    1.018857461705327e-07
+    4.151739121293431e-07
+     3.26653200865479e-08
+    5.425228205519541e-08
+    1.597951215495119e-07
+    4.193212385651605e-07
+ 2.18e+10    
+    4.189514133555438e-07
+    1.598146652654889e-07
+    4.152990289662314e-07
+    5.430221615025982e-08
+    1.019411792777907e-07
+    4.152383922854923e-07
+    3.270255085941718e-08
+    5.430042759074259e-08
+    1.598621253572115e-07
+    4.193979226873327e-07
+ 2.19e+10    
+    4.190281906356292e-07
+    1.598816612332757e-07
+    4.153634413796742e-07
+      5.4350206224342e-08
+    1.019965992027332e-07
+    4.153029596687778e-07
+    3.273955794118856e-08
+    5.434844018702423e-08
+    1.599291666610586e-07
+     4.19474735978337e-07
+ 2.2e+10     
+    4.191050988745256e-07
+    1.599486955212369e-07
+       4.154279439755e-07
+    5.439806299147981e-08
+    1.020520066447561e-07
+    4.153676151307865e-07
+    3.277634120339774e-08
+    5.439631999774925e-08
+    1.599962462896857e-07
+    4.195516792758543e-07
+ 2.21e+10    
+    4.191821388973855e-07
+    1.600157689434677e-07
+    4.154925375565719e-07
+     5.44457866119576e-08
+    1.021074022830502e-07
+    4.154323595032682e-07
+    3.281290053243036e-08
+     5.44440671837694e-08
+    1.600633650614017e-07
+     4.19628753410537e-07
+ 2.22e+10    
+    4.192593115222952e-07
+    1.600828823037871e-07
+    4.155572229061647e-07
+    5.449337725295783e-08
+     1.02162786777121e-07
+    4.154971935986541e-07
+     3.28492358291616e-08
+    5.449168191278429e-08
+    1.601305237842541e-07
+     4.19705959206015e-07
+ 2.23e+10    
+    4.193366175602896e-07
+    1.601500363958053e-07
+    4.156220007885065e-07
+    5.454083508827038e-08
+    1.022181607672935e-07
+    4.155621182105548e-07
+    3.288534700860201e-08
+    5.453916435905282e-08
+    1.601977232560927e-07
+    4.197832974789092e-07
+ 2.24e+10    
+    4.194140578153682e-07
+    1.602172320029896e-07
+    4.156868719492971e-07
+    5.458816029800715e-08
+    1.022735248752019e-07
+    4.156271341142484e-07
+     3.29212339995483e-08
+    5.458651470310906e-08
+    1.602649642646318e-07
+    4.198607690388427e-07
+ 2.25e+10    
+    4.194916330845079e-07
+    1.602844698987308e-07
+    4.157518371162137e-07
+    5.463535306832192e-08
+    1.023288797042646e-07
+     4.15692242067151e-07
+    3.295689674423996e-08
+    5.463373313148405e-08
+    1.603322475875141e-07
+    4.199383746884544e-07
+ 2.26e+10    
+    4.195693441576865e-07
+    1.603517508464109e-07
+    4.158168969994008e-07
+    5.468241359113632e-08
+    1.023842258401462e-07
+    4.157574428092745e-07
+    3.299233519802159e-08
+    5.468081983643302e-08
+    1.603995739923746e-07
+    4.200161152234153e-07
+ 2.27e+10    
+    4.196471918179022e-07
+    1.604190755994691e-07
+    4.158820522919429e-07
+    5.472934206387002e-08
+     1.02439563851205e-07
+    4.158227370636701e-07
+    3.302754932901014e-08
+    5.472777501566751e-08
+    1.604669442369041e-07
+    4.200939914324464e-07
+ 2.28e+10    
+    4.197251768411909e-07
+    1.604864449014687e-07
+     4.15947303670326e-07
+    5.477613868917752e-08
+    1.024948942889286e-07
+    4.158881255368616e-07
+    3.306253911776796e-08
+      5.4774598872093e-08
+    1.605343590689141e-07
+    4.201720040973369e-07
+ 2.29e+10    
+    4.198032999966558e-07
+    1.605538594861647e-07
+    4.160126517948819e-07
+    5.482280367468912e-08
+    1.025502176883564e-07
+    4.159536089192639e-07
+    3.309730455698098e-08
+    5.482129161355185e-08
+    1.606018192264007e-07
+    4.202501539929652e-07
+ 2.3e+10     
+     4.19881562046485e-07
+    1.606213200775698e-07
+    4.160780973102203e-07
+    5.486933723275792e-08
+    1.026055345684902e-07
+    4.160191878855881e-07
+    3.313184565114211e-08
+    5.486785345257125e-08
+    1.606693254376097e-07
+    4.203284418873202e-07
+ 2.31e+10    
+    4.199599637459816e-07
+    1.606888273900229e-07
+    4.161436408456498e-07
+    5.491573958021147e-08
+     1.02660845432693e-07
+    4.160848630952378e-07
+    3.316616241623985e-08
+    5.491428460611646e-08
+    1.607368784211008e-07
+    4.204068685415237e-07
+ 2.32e+10    
+    4.200385058435891e-07
+    1.607563821282547e-07
+    4.162092830155812e-07
+    5.496201093810899e-08
+    1.027161507690768e-07
+    4.161506351926945e-07
+    3.320025487945214e-08
+    5.496058529534894e-08
+    1.608044788858133e-07
+    4.204854347098568e-07
+ 2.33e+10    
+    4.201171890809179e-07
+    1.608239849874549e-07
+    4.162750244199215e-07
+    5.500815153150322e-08
+    1.027714510508788e-07
+     4.16216504807886e-07
+    3.323412307884511e-08
+     5.50067557453898e-08
+    1.608721275311302e-07
+    4.205641411397816e-07
+ 2.34e+10    
+    4.201960141927759e-07
+      1.6089163665334e-07
+    4.163408656444578e-07
+    5.505416158920781e-08
+    1.028267467368278e-07
+    4.162824725565518e-07
+    3.326776706307702e-08
+    5.505279618508806e-08
+     1.60939825046944e-07
+    4.206429885719717e-07
+ 2.35e+10    
+    4.202749819071943e-07
+    1.609593378022186e-07
+    4.164068072612251e-07
+    5.510004134356934e-08
+       1.028820382715e-07
+    4.163485390405934e-07
+    3.330118689110697e-08
+    5.509870684679393e-08
+     1.61007572113721e-07
+    4.207219777403355e-07
+ 2.36e+10    
+    4.203540929454631e-07
+    1.610270891010597e-07
+     4.16472849828867e-07
+     5.51457910302443e-08
+    1.029373260856647e-07
+    4.164147048484149e-07
+    3.333438263190875e-08
+    5.514448796613684e-08
+    1.610753694025675e-07
+    4.208011093720481e-07
+ 2.37e+10    
+    4.204333480221599e-07
+    1.610948912075589e-07
+    4.165389938929836e-07
+    5.519141088798117e-08
+    1.029926105966209e-07
+    4.164809705552546e-07
+    3.336735436418934e-08
+    5.519013978180879e-08
+     1.61143217575294e-07
+    4.208803841875774e-07
+ 2.38e+10    
+    4.205127478451802e-07
+     1.61162744770204e-07
+    4.166052399864689e-07
+    5.523690115840716e-08
+    1.030478922085243e-07
+    4.165473367235091e-07
+    3.340010217611232e-08
+    5.523566253535163e-08
+    1.612111172844809e-07
+    4.209598029007168e-07
+ 2.39e+10    
+    4.205922931157729e-07
+    1.612306504283428e-07
+    4.166715886298375e-07
+    5.528226208581976e-08
+    1.031031713127054e-07
+    4.166138039030447e-07
+    3.343262616502594e-08
+    5.528105647095016e-08
+    1.612790691735433e-07
+    4.210393662186136e-07
+ 2.4e+10     
+    4.206719845285737e-07
+    1.612986088122487e-07
+    4.167380403315446e-07
+    5.532749391698281e-08
+    1.031584482879785e-07
+    4.166803726314997e-07
+    3.346492643719595e-08
+    5.532632183522873e-08
+    1.613470738767961e-07
+    4.211190748418022e-07
+ 2.41e+10    
+    4.207518227716356e-07
+    1.613666205431872e-07
+    4.168045955882935e-07
+    5.537259690092773e-08
+    1.032137235009442e-07
+    4.167470434345843e-07
+    3.349700310754304e-08
+    5.537145887705369e-08
+    1.614151320195195e-07
+    4.211989294642352e-07
+ 2.42e+10    
+    4.208318085264685e-07
+    1.614346862334811e-07
+    4.168712548853328e-07
+    5.541757128875871e-08
+    1.032689973062804e-07
+    4.168138168263637e-07
+    3.352885629938479e-08
+    5.541646784733923e-08
+    1.614832442180231e-07
+    4.212789307733168e-07
+ 2.43e+10    
+    4.209119424680712e-07
+    1.615028064865777e-07
+    4.169380186967493e-07
+    5.546241733346288e-08
+    1.033242700470285e-07
+     4.16880693309539e-07
+    3.356048614418229e-08
+    5.546134899885869e-08
+    1.615514110797115e-07
+    4.213590794499359e-07
+ 2.44e+10    
+     4.20992225264967e-07
+    1.615709818971131e-07
+    4.170048874857485e-07
+    5.550713528972485e-08
+    1.033795420548708e-07
+    4.169476733757177e-07
+    3.359189278129101e-08
+    5.550610258605962e-08
+    1.616196332031483e-07
+    4.214393761685001e-07
+ 2.45e+10    
+    4.210726575792413e-07
+    1.616392130509787e-07
+     4.17071861704928e-07
+     5.55517254137456e-08
+    1.034348136503998e-07
+    4.170147575056774e-07
+    3.362307635771641e-08
+    5.555072886488386e-08
+    1.616879111781221e-07
+    4.215198215969714e-07
+ 2.46e+10    
+    4.211532400665775e-07
+    1.617075005253859e-07
+    4.171389417965419e-07
+    5.559618796306567e-08
+    1.034900851433819e-07
+    4.170819461696213e-07
+    3.365403702787347e-08
+    5.559522809259111e-08
+     1.61756245585709e-07
+    4.216004163968973e-07
+ 2.47e+10    
+    4.212339733762937e-07
+    1.617758448889317e-07
+    4.172061281927602e-07
+    5.564052319639294e-08
+    1.035453568330131e-07
+    4.171492398274295e-07
+    3.368477495335103e-08
+    5.563960052758778e-08
+    1.618246369983388e-07
+    4.216811612234513e-07
+ 2.48e+10    
+    4.213148581513801e-07
+    1.618442467016627e-07
+    4.172734213159164e-07
+    5.568473137343427e-08
+    1.036006290081677e-07
+    4.172166389288974e-07
+    3.371529030268001e-08
+    5.568384642925928e-08
+     1.61893085979858e-07
+    4.217620567254647e-07
+ 2.49e+10    
+    4.213958950285363e-07
+    1.619127065151409e-07
+    4.173408215787517e-07
+    5.572881275473145e-08
+     1.03655901947642e-07
+     4.17284143913974e-07
+    3.374558325110592e-08
+    5.572796605780676e-08
+    1.619615930855947e-07
+    4.218431035454648e-07
+ 2.5e+10     
+    4.214770846382108e-07
+    1.619812248725072e-07
+    4.174083293846499e-07
+    5.577276760150158e-08
+    1.037111759203897e-07
+    4.173517552129902e-07
+    3.377565398036577e-08
+    5.577195967408793e-08
+    1.620301588624219e-07
+    4.219243023197111e-07
+ 2.51e+10    
+    4.215584276046363e-07
+    1.620498023085461e-07
+    4.174759451278656e-07
+    5.581659617548085e-08
+    1.037664511857531e-07
+    4.174194732468791e-07
+    3.380550267846874e-08
+    5.581582753946193e-08
+    1.620987838488214e-07
+     4.22005653678231e-07
+ 2.52e+10    
+    4.216399245458717e-07
+    1.621184393497495e-07
+    4.175436691937464e-07
+     5.58602987387732e-08
+    1.038217279936871e-07
+    4.174872984273962e-07
+    3.383512953948112e-08
+    5.585956991563805e-08
+    1.621674685749474e-07
+    4.220871582448575e-07
+ 2.53e+10    
+    4.217215760738366e-07
+    1.621871365143806e-07
+    4.176115019589494e-07
+    5.590387555370171e-08
+    1.038770065849777e-07
+    4.175552311573253e-07
+    3.386453476331518e-08
+    5.590318706452856e-08
+    1.622362135626898e-07
+    4.221688166372683e-07
+ 2.54e+10    
+    4.218033827943547e-07
+    1.622558943125372e-07
+    4.176794437916492e-07
+    5.594732688266511e-08
+    1.039322871914555e-07
+    4.176232718306873e-07
+    3.389371855552207e-08
+    5.594667924810515e-08
+    1.623050193257372e-07
+    4.222506294670199e-07
+ 2.55e+10    
+    4.218853453071887e-07
+    1.623247132462146e-07
+    4.177474950517408e-07
+    5.599065298799736e-08
+    1.039875700362032e-07
+    4.176914208329358e-07
+    3.392268112708848e-08
+     5.59900467282593e-08
+    1.623738863696397e-07
+    4.223325973395882e-07
+ 2.56e+10    
+    4.219674642060822e-07
+    1.623935938093694e-07
+    4.178156560910388e-07
+    5.603385413183127e-08
+    1.040428553337581e-07
+    4.177596785411546e-07
+    3.395142269423739e-08
+    5.603328976666661e-08
+    1.624428151918722e-07
+    4.224147208544059e-07
+ 2.57e+10    
+    4.220497400787974e-07
+    1.624625364879813e-07
+    4.178839272534683e-07
+    5.607693057596539e-08
+    1.040981432903095e-07
+    4.178280453242409e-07
+    3.397994347823237e-08
+    5.607640862465427e-08
+    1.625118062818959e-07
+       4.224970006049e-07
+ 2.58e+10    
+    4.221321735071562e-07
+    1.625315417601163e-07
+     4.17952308875251e-07
+    5.611988258173531e-08
+    1.041534341038913e-07
+    4.178965215430937e-07
+    3.400824370518584e-08
+    5.611940356307262e-08
+    1.625808601212214e-07
+    4.225794371785307e-07
+ 2.59e+10    
+    4.222147650670776e-07
+    1.626006100959881e-07
+    4.180208012850856e-07
+    5.616271040988762e-08
+    1.042087279645693e-07
+    4.179651075507885e-07
+    3.403632360587088e-08
+    5.616227484216999e-08
+    1.626499771834702e-07
+    4.226620311568289e-07
+ 2.6e+10     
+    4.222975153286188e-07
+    1.626697419580205e-07
+    4.180894048043248e-07
+     5.62054143204581e-08
+    1.042640250546249e-07
+    4.180338036927534e-07
+    3.406418341553695e-08
+     5.62050227214713e-08
+    1.627191579344363e-07
+    4.227447831154372e-07
+ 2.61e+10    
+    4.223804248560146e-07
+    1.627389378009089e-07
+    4.181581197471465e-07
+    5.624799457265313e-08
+    1.043193255487334e-07
+    4.181026103069355e-07
+     3.40918233737289e-08
+    5.624764745965964e-08
+    1.627884028321482e-07
+    4.228276936241452e-07
+ 2.62e+10    
+    4.224634942077168e-07
+    1.628081980716813e-07
+    4.182269464207177e-07
+    5.629045142473431e-08
+     1.04374629614138e-07
+    4.181715277239671e-07
+    3.411924372410984e-08
+    5.629014931446184e-08
+    1.628577123269297e-07
+    4.229107632469306e-07
+ 2.63e+10    
+    4.225467239364333e-07
+    1.628775232097596e-07
+    4.182958851253581e-07
+    5.633278513390657e-08
+    1.044299374108198e-07
+    4.182405562673247e-07
+    3.414644471428738e-08
+    5.633252854253704e-08
+     1.62927086861461e-07
+    4.229939925419974e-07
+ 2.64e+10    
+    4.226301145891692e-07
+    1.629469136470205e-07
+    4.183649361546956e-07
+    5.637499595620977e-08
+    1.044852490916644e-07
+    4.183096962534857e-07
+    3.417342659564336e-08
+    5.637478539936813e-08
+    1.629965268708396e-07
+    4.230773820618144e-07
+ 2.65e+10    
+    4.227136667072661e-07
+    1.630163698078553e-07
+    4.184340997958201e-07
+    5.641708414641302e-08
+    1.045405648026226e-07
+    4.183789479920788e-07
+    3.420018962316711e-08
+    5.641692013915746e-08
+      1.6306603278264e-07
+    4.231609323531543e-07
+ 2.66e+10    
+      4.2279738082644e-07
+    1.630858921092304e-07
+    4.185033763294303e-07
+    5.645904995791273e-08
+    1.045958846828695e-07
+    4.184483117860326e-07
+    3.422673405529198e-08
+    5.645893301472444e-08
+    1.631356050169751e-07
+     4.23244643957133e-07
+ 2.67e+10    
+    4.228812574768245e-07
+    1.631554809607474e-07
+    4.185727660299787e-07
+    5.650089364263327e-08
+    1.046512088649581e-07
+    4.185177879317176e-07
+    3.425306015373528e-08
+    5.650082427740722e-08
+    1.632052439865545e-07
+    4.233285174092478e-07
+ 2.68e+10    
+    4.229652971830072e-07
+    1.632251367647021e-07
+    4.186422691658112e-07
+    5.654261545093122e-08
+      1.0470653747497e-07
+    4.185873767190904e-07
+    3.427916818334149e-08
+      5.6542594176967e-08
+    1.632749500967457e-07
+     4.23412553239417e-07
+ 2.69e+10    
+    4.230495004640712e-07
+     1.63294859916144e-07
+    4.187118859993041e-07
+    5.658421563150197e-08
+    1.047618706326628e-07
+     4.18657078431824e-07
+    3.430505841192877e-08
+    5.658424296149528e-08
+    1.633447237456321e-07
+    4.234967519720189e-07
+ 2.7e+10     
+    4.231338678336336e-07
+     1.63364650802935e-07
+    4.187816167869954e-07
+    5.662569443128986e-08
+    1.048172084516128e-07
+    4.187268933474453e-07
+     3.43307311101386e-08
+    5.662577087732416e-08
+    1.634145653240726e-07
+    4.235811141259281e-07
+ 2.71e+10    
+    4.232183997998859e-07
+     1.63434509805808e-07
+    4.188514617797153e-07
+    5.666705209540083e-08
+    1.048725510393564e-07
+    4.187968217374619e-07
+    3.435618655128869e-08
+    5.666717816893959e-08
+    1.634844752157603e-07
+    4.236656402145601e-07
+ 2.72e+10    
+    4.233030968656331e-07
+    1.635044372984258e-07
+    4.189214212227109e-07
+    5.670828886701827e-08
+    1.049278984975262e-07
+    4.188668638674901e-07
+    3.438142501122894e-08
+    5.670846507889732e-08
+    1.635544537972811e-07
+    4.237503307459035e-07
+ 2.73e+10    
+    4.233879595283324e-07
+    1.635744336474381e-07
+    4.189914953557671e-07
+    5.674940498732112e-08
+    1.049832509219853e-07
+    4.189370199973755e-07
+    3.440644676820044e-08
+     5.67496318477416e-08
+     1.63624501438171e-07
+    4.238351862225624e-07
+ 2.74e+10    
+    4.234729882801331e-07
+    1.636444992125396e-07
+    4.190616844133271e-07
+    5.679040069540528e-08
+    1.050386084029577e-07
+    4.190072903813139e-07
+     3.44312521026977e-08
+    5.679067871392686e-08
+    1.636946185009751e-07
+    4.239202071417955e-07
+ 2.75e+10    
+    4.235581836079156e-07
+    1.637146343465273e-07
+    4.191319886246057e-07
+    5.683127622820728e-08
+    1.050939710251561e-07
+    4.190776752679686e-07
+    3.445584129733358e-08
+    5.683160591374154e-08
+    1.637648053413038e-07
+    4.240053939955527e-07
+ 2.76e+10    
+    4.236435459933312e-07
+    1.637848393953577e-07
+    4.192024082137053e-07
+    5.687203182043089e-08
+    1.051493388679071e-07
+    4.191481749005813e-07
+    3.448021463670756e-08
+    5.687241368123531e-08
+    1.638350623078913e-07
+    4.240907472705143e-07
+ 2.77e+10    
+    4.237290759128399e-07
+    1.638551146982034e-07
+    4.192729433997215e-07
+    5.691266770447598e-08
+    1.052047120052728e-07
+    4.192187895170865e-07
+    3.450437240727648e-08
+     5.69131022481481e-08
+    1.639053897426517e-07
+    4.241762674481304e-07
+ 2.78e+10    
+    4.238147738377493e-07
+    1.639254605875089e-07
+    4.193435943968508e-07
+    5.695318411037034e-08
+    1.052600905061701e-07
+    4.192895193502152e-07
+    3.452831489722857e-08
+    5.695367184384209e-08
+    1.639757879807357e-07
+    4.242619550046583e-07
+ 2.79e+10    
+    4.239006402342541e-07
+    1.639958773890475e-07
+    4.194143614144957e-07
+    5.699358126570349e-08
+    1.053154744344876e-07
+    4.193603646276052e-07
+    3.455204239636006e-08
+    5.699412269523623e-08
+    1.640462573505869e-07
+    4.243478104112012e-07
+ 2.8e+10     
+     4.23986675563474e-07
+    1.640663654219762e-07
+    4.194852446573631e-07
+     5.70338593955634e-08
+    1.053708638491991e-07
+    4.194313255718985e-07
+    3.457555519595456e-08
+    5.703445502674267e-08
+    1.641167981739978e-07
+    4.244338341337452e-07
+ 2.81e+10    
+    4.240728802814926e-07
+    1.641369249988919e-07
+    4.195562443255649e-07
+    5.707401872247516e-08
+    1.054262588044754e-07
+    4.195024024008453e-07
+    3.459885358866547e-08
+    5.707466906020633e-08
+    1.641874107661656e-07
+    4.245200266332001e-07
+ 2.82e+10    
+    4.241592548393951e-07
+    1.642075564258859e-07
+    4.196273606147126e-07
+    5.711405946634238e-08
+    1.054816593497933e-07
+    4.195735953273997e-07
+    3.462193786840075e-08
+    5.711476501484611e-08
+    1.642580954357473e-07
+    4.246063883654331e-07
+ 2.83e+10    
+    4.242457996833084e-07
+    1.642782600025988e-07
+    4.196985937160097e-07
+    5.715398184439072e-08
+    1.055370655300417e-07
+    4.196449045598151e-07
+    3.464480833021072e-08
+    5.715474310719873e-08
+    1.643288524849145e-07
+    4.246929197813112e-07
+ 2.84e+10    
+    4.243325152544347e-07
+    1.643490360222747e-07
+    4.197699438163449e-07
+    5.719378607111349e-08
+    1.055924773856267e-07
+    4.197163303017381e-07
+    3.466746527017815e-08
+    5.719460355106496e-08
+    1.643996822094088e-07
+    4.247796213267352e-07
+ 2.85e+10    
+    4.244194019890951e-07
+    1.644198847718156e-07
+     4.19841411098377e-07
+    5.723347235821968e-08
+     1.05647894952573e-07
+    4.197878727522975e-07
+    3.468990898531119e-08
+    5.723434655745758e-08
+    1.644705848985952e-07
+      4.2486649344268e-07
+ 2.86e+10    
+     4.24506460318762e-07
+    1.644908065318354e-07
+    4.199129957406254e-07
+    5.727304091458422e-08
+    1.057033182626234e-07
+    4.198595321061931e-07
+    3.471213977343884e-08
+    5.727397233455187e-08
+    1.645415608355172e-07
+    4.249535365652295e-07
+ 2.87e+10    
+    4.245936906701009e-07
+     1.64561801576712e-07
+    4.199846979175495e-07
+    5.731249194620008e-08
+     1.05758747343337e-07
+    4.199313085537828e-07
+     3.47341579331088e-08
+    5.731348108763807e-08
+    1.646126102969493e-07
+    4.250407511256157e-07
+ 2.88e+10    
+    4.246810934650059e-07
+    1.646328701746423e-07
+     4.20056517799634e-07
+    5.735182565613271e-08
+    1.058141822181849e-07
+    4.200032022811671e-07
+    3.475596376348804e-08
+    5.735287301907598e-08
+    1.646837335534514e-07
+    4.251281375502547e-07
+ 2.89e+10    
+    4.247686691206352e-07
+    1.647040125876934e-07
+    4.201284555534668e-07
+     5.73910422444761e-08
+    1.058696229066427e-07
+    4.200752134702687e-07
+    3.477755756426555e-08
+    5.739214832825142e-08
+    1.647549308694218e-07
+    4.252156962607857e-07
+ 2.9e+10     
+    4.248564180494519e-07
+    1.647752290718557e-07
+    4.202005113418179e-07
+     5.74301419083115e-08
+    1.059250694242828e-07
+    4.201473422989155e-07
+    3.479893963555771e-08
+    5.743130721153487e-08
+     1.64826202503149e-07
+    4.253034276741039e-07
+ 2.91e+10    
+    4.249443406592578e-07
+    1.648465198770951e-07
+    4.202726853237142e-07
+    5.746912484166739e-08
+     1.05980521782864e-07
+    4.202195889409176e-07
+    3.482011027781609e-08
+    5.747034986224197e-08
+    1.648975487068652e-07
+    4.253913322024018e-07
+ 2.92e+10    
+     4.25032437353232e-07
+    1.649178852474043e-07
+    4.203449776545133e-07
+     5.75079912354819e-08
+    1.060359799904183e-07
+     4.20291953566144e-07
+    3.484106979173727e-08
+    5.750927647059571e-08
+    1.649689697267977e-07
+    4.254794102532017e-07
+ 2.93e+10    
+    4.251207085299661e-07
+    1.649893254208547e-07
+    4.204173884859769e-07
+    5.754674127756659e-08
+     1.06091444051338e-07
+    4.203644363405967e-07
+    3.486181847817536e-08
+    5.754808722369103e-08
+    1.650404658032212e-07
+    4.255676622293958e-07
+ 2.94e+10    
+    4.252091545835008e-07
+     1.65060840629647e-07
+    4.204899179663392e-07
+    5.758537515257248e-08
+    1.061469139664585e-07
+    4.204370374264844e-07
+    3.488235663805656e-08
+    5.758678230546047e-08
+    1.651120371705085e-07
+    4.256560885292783e-07
+ 2.95e+10    
+    4.252977759033634e-07
+    1.651324311001629e-07
+    4.205625662403781e-07
+    5.762389304195786e-08
+    1.062023897331417e-07
+    4.205097569822948e-07
+    3.490268457229606e-08
+     5.76253618966424e-08
+    1.651836840571824e-07
+    4.257446895465853e-07
+ 2.96e+10    
+     4.25386572874602e-07
+    1.652040970530144e-07
+    4.206353334494782e-07
+    5.766229512395719e-08
+    1.062578713453554e-07
+    4.205825951628596e-07
+    3.492280258171706e-08
+    5.766382617475035e-08
+    1.652554066859659e-07
+    4.258334656705278e-07
+ 2.97e+10    
+    4.254755458778226e-07
+    1.652758387030945e-07
+    4.207082197316998e-07
+    5.770058157355291e-08
+    1.063133587937533e-07
+    4.206555521194289e-07
+    3.494271096697212e-08
+    5.770217531404437e-08
+     1.65327205273833e-07
+    4.259224172858299e-07
+ 2.98e+10    
+    4.255646952892233e-07
+     1.65347656259627e-07
+    4.207812252218405e-07
+    5.773875256244762e-08
+    1.063688520657519e-07
+    4.207286279997327e-07
+    3.496241002846649e-08
+    5.774040948550408e-08
+    1.653990800320584e-07
+    4.260115447727613e-07
+ 2.99e+10    
+    4.256540214806321e-07
+     1.65419549926216e-07
+    4.208543500514981e-07
+     5.77768082590388e-08
+     1.06424351145606e-07
+    4.208018229480481e-07
+    3.498190006628359e-08
+    5.777852885680313e-08
+    1.654710311662679e-07
+    4.261008485071754e-07
+ 3e+10       
+    4.257435248195398e-07
+    1.654915199008949e-07
+    4.209275943491312e-07
+     5.78147488283949e-08
+    1.064798560144831e-07
+     4.20875137105262e-07
+    3.500118138011272e-08
+    5.781653359228551e-08
+    1.655430588764872e-07
+    4.261903288605434e-07
+ 3.01e+10    
+    4.258332056691353e-07
+    1.655635663761747e-07
+    4.210009582401166e-07
+    5.785257443223268e-08
+     1.06535366650536e-07
+    4.209485706089326e-07
+    3.502025426917855e-08
+    5.785442385294326e-08
+    1.656151633571916e-07
+    4.262799861999891e-07
+ 3.02e+10    
+    4.259230643883433e-07
+    1.656356895390939e-07
+    4.210744418468115e-07
+    5.789028522889668e-08
+    1.065908830289745e-07
+    4.210221235933519e-07
+    3.503911903217294e-08
+    5.789219979639571e-08
+    1.656873447973545e-07
+    4.263698208883238e-07
+ 3.03e+10    
+    4.260131013318549e-07
+    1.657078895712648e-07
+    4.211480452886048e-07
+     5.79278813733396e-08
+    1.066464051221344e-07
+     4.21095796189603e-07
+    3.505777596718841e-08
+    5.792986157687039e-08
+    1.657596033804958e-07
+    4.264598332840812e-07
+ 3.04e+10    
+    4.261033168501655e-07
+    1.657801666489231e-07
+    4.212217686819758e-07
+    5.796536301710438e-08
+    1.067019328995465e-07
+    4.211695885256191e-07
+    3.507622537165384e-08
+    5.796740934518508e-08
+    1.658319392847303e-07
+    4.265500237415522e-07
+ 3.05e+10    
+    4.261937112896057e-07
+    1.658525209429735e-07
+    4.212956121405462e-07
+    5.800273030830792e-08
+    1.067574663280034e-07
+    4.212435007262397e-07
+    3.509446754227191e-08
+    5.800484324873174e-08
+    1.659043526828154e-07
+    4.266403926108182e-07
+ 3.06e+10    
+    4.262842849923796e-07
+    1.659249526190387e-07
+    4.213695757751345e-07
+    5.803998339162589e-08
+    1.068130053716253e-07
+    4.213175329132669e-07
+     3.51125027749586e-08
+    5.804216343146124e-08
+    1.659768437421988e-07
+    4.267309402377868e-07
+ 3.07e+10    
+    4.263750382965952e-07
+    1.659974618375053e-07
+    4.214436596938049e-07
+    5.807712240827908e-08
+    1.068685499919243e-07
+    4.213916852055184e-07
+    3.513033136478445e-08
+    5.807937003387011e-08
+    1.660494126250651e-07
+    4.268216669642231e-07
+ 3.08e+10    
+    4.264659715363003e-07
+    1.660700487535701e-07
+    4.215178640019198e-07
+    5.811414749602098e-08
+    1.069241001478678e-07
+    4.214659577188811e-07
+    3.514795360591761e-08
+    5.811646319298821e-08
+    1.661220594883832e-07
+     4.26912573127787e-07
+ 3.09e+10    
+    4.265570850415143e-07
+    1.661427135172868e-07
+    4.215921888021873e-07
+     5.81510587891268e-08
+    1.069796557959403e-07
+    4.215403505663643e-07
+     3.51653697915688e-08
+    5.815344304236759e-08
+    1.661947844839531e-07
+    4.270036590620635e-07
+ 3.1e+10     
+    4.266483791382627e-07
+    1.662154562736117e-07
+    4.216666341947112e-07
+    5.818785641838363e-08
+    1.070352168902039e-07
+    4.216148638581489e-07
+    3.518258021393799e-08
+    5.819030971207317e-08
+    1.662675877584509e-07
+    4.270949250965983e-07
+ 3.11e+10    
+    4.267398541486109e-07
+    1.662882771624494e-07
+    4.217412002770352e-07
+    5.822454051108202e-08
+    1.070907833823583e-07
+    4.216894977016371e-07
+    3.519958516416291e-08
+    5.822706332867423e-08
+    1.663404694534761e-07
+    4.271863715569294e-07
+ 3.12e+10    
+    4.268315103906949e-07
+    1.663611763186975e-07
+     4.21815887144191e-07
+    5.826111119100852e-08
+    1.071463552217987e-07
+    4.217642522015025e-07
+    3.521638493226916e-08
+    5.826370401523695e-08
+    1.664134297055961e-07
+    4.272779987646218e-07
+ 3.13e+10    
+    4.269233481787565e-07
+    1.664341538722919e-07
+    4.218906948887423e-07
+    5.829756857843969e-08
+    1.072019323556736e-07
+    4.218391274597368e-07
+    3.523297980712205e-08
+    5.830023189131882e-08
+    1.664864686463919e-07
+    4.273698070372988e-07
+ 3.14e+10    
+    4.270153678231739e-07
+    1.665072099482516e-07
+    4.219656236008283e-07
+    5.833391279013716e-08
+    1.072575147289404e-07
+    4.219141235756968e-07
+     3.52493700763803e-08
+    5.833664707296356e-08
+    1.665595864025032e-07
+    4.274617966886754e-07
+ 3.15e+10    
+    4.271075696304958e-07
+    1.665803446667226e-07
+    4.220406733682079e-07
+     5.83701439393438e-08
+    1.073131022844211e-07
+    4.219892406461509e-07
+    3.526555602645102e-08
+    5.837294967269733e-08
+    1.666327830956726e-07
+    4.275539680285915e-07
+ 3.16e+10    
+    4.271999539034721e-07
+    1.666535581430217e-07
+    4.221158442763003e-07
+    5.840626213578089e-08
+    1.073686949628559e-07
+    4.220644787653209e-07
+    3.528153794244661e-08
+    5.840913979952646e-08
+    1.667060588427899e-07
+    4.276463213630422e-07
+ 3.17e+10    
+    4.272925209410876e-07
+    1.667268504876808e-07
+    4.221911364082271e-07
+    5.844226748564681e-08
+    1.074242927029563e-07
+    4.221398380249311e-07
+    3.529731610814315e-08
+    5.844521755893551e-08
+    1.667794137559361e-07
+     4.27738856994211e-07
+ 3.18e+10    
+    4.273852710385909e-07
+    1.668002218064892e-07
+    4.222665498448514e-07
+    5.847816009161611e-08
+    1.074798954414575e-07
+    4.222153185142454e-07
+    3.531289080594039e-08
+    5.848118305288723e-08
+    1.668528479424275e-07
+    4.278315752205035e-07
+ 3.19e+10    
+    4.274782044875295e-07
+    1.668736722005381e-07
+    4.223420846648195e-07
+    5.851394005284035e-08
+    1.075355031131691e-07
+    4.222909203201149e-07
+    3.532826231682308e-08
+    5.851703637982274e-08
+    1.669263615048584e-07
+    4.279244763365756e-07
+ 3.2e+10     
+    4.275713215757794e-07
+    1.669472017662612e-07
+     4.22417740944596e-07
+    5.854960746494928e-08
+    1.075911156510253e-07
+    4.223666435270152e-07
+    3.534343092032418e-08
+    5.855277763466334e-08
+    1.669999545411442e-07
+    4.280175606333676e-07
+ 3.21e+10    
+    4.276646225875759e-07
+    1.670208105954794e-07
+    4.224935187585048e-07
+    5.858516242005355e-08
+    1.076467329861341e-07
+    4.224424882170881e-07
+    3.535839689448926e-08
+    5.858840690881306e-08
+    1.670736271445645e-07
+    4.281108283981352e-07
+ 3.22e+10    
+    4.277581078035451e-07
+    1.670944987754406e-07
+    4.225694181787633e-07
+      5.8620605006748e-08
+    1.077023550478258e-07
+    4.225184544701838e-07
+     3.53731605158424e-08
+    5.862392429016195e-08
+     1.67147379403805e-07
+    4.282042799144797e-07
+ 3.23e+10    
+    4.278517775007359e-07
+    1.671682663888637e-07
+     4.22645439275522e-07
+     5.86559353101161e-08
+    1.077579817636997e-07
+    4.225945423638952e-07
+    3.538772205935377e-08
+    5.865932986309089e-08
+    1.672212114030001e-07
+    4.282979154623793e-07
+ 3.24e+10    
+    4.279456319526494e-07
+    1.672421135139782e-07
+    4.227215821168966e-07
+    5.869115341173518e-08
+    1.078136130596716e-07
+    4.226707519735987e-07
+    3.540208179840828e-08
+    5.869462370847656e-08
+     1.67295123221774e-07
+    4.283917353182216e-07
+ 3.25e+10    
+    4.280396714292689e-07
+    1.673160402245661e-07
+     4.22797846769004e-07
+    5.872625938968268e-08
+    1.078692488600185e-07
+    4.227470833724929e-07
+    3.541624000477592e-08
+    5.872980590369799e-08
+    1.673691149352826e-07
+    4.284857397548314e-07
+ 3.26e+10    
+    4.281338961970909e-07
+     1.67390046590003e-07
+    4.228742332959976e-07
+    5.876125331854316e-08
+    1.079248890874242e-07
+    4.228235366316325e-07
+    3.543019694858324e-08
+    5.876487652264345e-08
+    1.674431866142547e-07
+    4.285799290415034e-07
+ 3.27e+10    
+    4.282283065191557e-07
+     1.67464132675298e-07
+    4.229507417600986e-07
+    5.879613526941609e-08
+    1.079805336630225e-07
+     4.22900111819966e-07
+    3.544395289828644e-08
+     5.87998356357186e-08
+    1.675173383250326e-07
+    4.286743034440315e-07
+ 3.28e+10    
+    4.283229026550773e-07
+    1.675382985411345e-07
+    4.230273722216302e-07
+    5.883090530992485e-08
+    1.080361825064413e-07
+    4.229768090043703e-07
+    3.545750812064552e-08
+     5.88346833098551e-08
+    1.675915701296124e-07
+    4.287688632247391e-07
+ 3.29e+10    
+    4.284176848610709e-07
+    1.676125442439096e-07
+    4.231041247390494e-07
+    5.886556350422599e-08
+    1.080918355358445e-07
+    4.230536282496867e-07
+    3.547086288069992e-08
+    5.886941960852038e-08
+     1.67665882085685e-07
+    4.288636086425082e-07
+ 3.3e+10     
+    4.285126533899858e-07
+    1.676868698357742e-07
+     4.23180999368977e-07
+    5.890010991301968e-08
+    1.081474926679735e-07
+    4.231305696187528e-07
+    3.548401744174533e-08
+    5.890404459172781e-08
+    1.677402742466753e-07
+    4.289585399528118e-07
+ 3.31e+10    
+    4.286078084913317e-07
+    1.677612753646721e-07
+    4.232579961662318e-07
+    5.893454459356069e-08
+    1.082031538181888e-07
+    4.232076331724376e-07
+    3.549697206531186e-08
+      5.8938558316048e-08
+    1.678147466617818e-07
+    4.290536574077392e-07
+ 3.32e+10    
+    4.287031504113107e-07
+     1.67835760874379e-07
+    4.233351151838575e-07
+    5.896886759967048e-08
+    1.082588189005095e-07
+    4.232848189696735e-07
+    3.550972701114341e-08
+    5.897296083462062e-08
+    1.678892993760166e-07
+    4.291489612560288e-07
+ 3.33e+10    
+    4.287986793928424e-07
+     1.67910326404541e-07
+    4.234123564731538e-07
+    5.900307898174928e-08
+     1.08314487827653e-07
+    4.233621270674884e-07
+    3.552228253717816e-08
+    5.900725219716698e-08
+    1.679639324302438e-07
+    4.292444517430958e-07
+ 3.34e+10    
+    4.288943956755977e-07
+    1.679849719907136e-07
+     4.23489720083705e-07
+    5.903717878678999e-08
+    1.083701605110741e-07
+    4.234395575210386e-07
+    3.553463889953051e-08
+     5.90414324500033e-08
+    1.680386458612183e-07
+    4.293401291110616e-07
+ 3.35e+10    
+    4.289902994960233e-07
+    1.680596976643998e-07
+    4.235672060634105e-07
+    5.907116705839167e-08
+    1.084258368610029e-07
+    4.235171103836385e-07
+    3.554679635247402e-08
+    5.907550163605509e-08
+     1.68113439701625e-07
+    4.294359935987838e-07
+ 3.36e+10    
+    4.290863910873714e-07
+    1.681345034530869e-07
+    4.236448144585094e-07
+    5.910504383677421e-08
+    1.084815167864819e-07
+    4.235947857067913e-07
+     3.55587551484253e-08
+    5.910945979487109e-08
+    1.681883139801151e-07
+    4.295320454418814e-07
+ 3.37e+10    
+    4.291826706797278e-07
+    1.682093893802852e-07
+    4.237225453136119e-07
+    5.913880915879382e-08
+    1.085372001954032e-07
+    4.236725835402185e-07
+    3.557051553792963e-08
+    5.914330696263934e-08
+    1.682632687213457e-07
+    4.296282848727663e-07
+ 3.38e+10    
+    4.292791385000421e-07
+    1.682843554655655e-07
+    4.238003986717237e-07
+    5.917246305795885e-08
+    1.085928869945444e-07
+    4.237505039318911e-07
+    3.558207776964713e-08
+    5.917704317220272e-08
+    1.683383039460173e-07
+    4.297247121206716e-07
+ 3.39e+10    
+    4.293757947721516e-07
+    1.683594017245944e-07
+    4.238783745742723e-07
+    5.920600556444641e-08
+    1.086485770896043e-07
+    4.238285469280568e-07
+    3.559344209034033e-08
+     5.92106684530756e-08
+    1.684134196709094e-07
+    4.298213274116778e-07
+ 3.4e+10     
+    4.294726397168119e-07
+    1.684345281691728e-07
+    4.239564730611364e-07
+    5.923943670511935e-08
+    1.087042703852377e-07
+    4.239067125732691e-07
+    3.560460874486266e-08
+    5.924418283146112e-08
+    1.684886159089192e-07
+    4.299181309687415e-07
+ 3.41e+10    
+     4.29569673551724e-07
+    1.685097348072712e-07
+    4.240346941706669e-07
+    5.927275650354423e-08
+    1.087599667850895e-07
+    4.239850009104152e-07
+    3.561557797614823e-08
+    5.927758633026886e-08
+    1.685638926690976e-07
+    4.300151230117247e-07
+ 3.42e+10    
+    4.296668964915605e-07
+    1.685850216430665e-07
+    4.241130379397161e-07
+    5.930596498000942e-08
+    1.088156661918287e-07
+    4.240634119807431e-07
+     3.56263500252024e-08
+    5.931087896913328e-08
+    1.686392499566853e-07
+    4.301123037574197e-07
+ 3.43e+10    
+    4.297643087479935e-07
+    1.686603886769773e-07
+    4.241915044036599e-07
+    5.933906215154408e-08
+    1.088713685071812e-07
+    4.241419458238896e-07
+    3.563692513109357e-08
+    5.934406076443254e-08
+    1.687146877731495e-07
+    4.302096734195794e-07
+ 3.44e+10    
+    4.298619105297225e-07
+    1.687358359056997e-07
+    4.242700935964237e-07
+    5.937204803193773e-08
+    1.089270736319629e-07
+    4.242206024779056e-07
+    3.564730353094587e-08
+    5.937713172930795e-08
+    1.687902061162191e-07
+    4.303072322089418e-07
+ 3.45e+10    
+    4.299597020424995e-07
+    1.688113633222426e-07
+    4.243488055505044e-07
+    5.940492263175985e-08
+     1.08982781466111e-07
+    4.242993819792828e-07
+    3.565748545993289e-08
+    5.941009187368392e-08
+    1.688658049799209e-07
+    4.304049803332586e-07
+ 3.46e+10    
+    4.300576834891571e-07
+    1.688869709159628e-07
+    4.244276402969962e-07
+    5.943768595838062e-08
+    1.090384919087159e-07
+    4.243782843629798e-07
+    3.566747115127239e-08
+    5.944294120428855e-08
+    1.689414843546144e-07
+    4.305029179973221e-07
+ 3.47e+10    
+     4.30155855069633e-07
+    1.689626586725991e-07
+    4.245065978656124e-07
+    5.947033801599173e-08
+     1.09094204858052e-07
+    4.244573096624463e-07
+    3.567726083622194e-08
+    5.947567972467441e-08
+    1.690172442270266e-07
+    4.306010454029913e-07
+ 3.48e+10    
+    4.302542169809982e-07
+    1.690384265743079e-07
+    4.245856782847081e-07
+     5.95028788056279e-08
+    1.091499202116082e-07
+    4.245364579096485e-07
+    3.568685474407554e-08
+    5.950830743524013e-08
+    1.690930845802874e-07
+    4.306993627492193e-07
+ 3.49e+10    
+    4.303527694174839e-07
+    1.691142745996963e-07
+    4.246648815813019e-07
+    5.953530832518873e-08
+    1.092056378661177e-07
+     4.24615729135095e-07
+    3.569625310216115e-08
+    5.954082433325225e-08
+    1.691690053939633e-07
+    4.307978702320786e-07
+ 3.5e+10     
+    4.304515125705032e-07
+    1.691902027238563e-07
+    4.247442077811002e-07
+    5.956762656946109e-08
+    1.092613577175873e-07
+    4.246951233678581e-07
+    3.570545613583908e-08
+    5.957323041286764e-08
+    1.692450066440919e-07
+    4.308965680447878e-07
+ 3.51e+10    
+    4.305504466286822e-07
+    1.692662109183988e-07
+     4.24823656908516e-07
+    5.959983353014186e-08
+    1.093170796613266e-07
+    4.247746406355987e-07
+    3.571446406850145e-08
+    5.960552566515632e-08
+    1.693210883032158e-07
+    4.309954563777383e-07
+ 3.52e+10    
+    4.306495717778819e-07
+    1.693422991514869e-07
+    4.249032289866925e-07
+    5.963192919586147e-08
+    1.093728035919764e-07
+     4.24854280964591e-07
+    3.572327712157225e-08
+    5.963771007812471e-08
+    1.693972503404161e-07
+     4.31094535418519e-07
+ 3.53e+10    
+     4.30748888201225e-07
+    1.694184673878682e-07
+    4.249829240375229e-07
+    5.966391355220701e-08
+     1.09428529403536e-07
+    4.249340443797431e-07
+    3.573189551450848e-08
+    5.966978363673923e-08
+    1.694734927213457e-07
+    4.311938053519427e-07
+ 3.54e+10    
+     4.30848396079121e-07
+     1.69494715588909e-07
+    4.250627420816698e-07
+    5.969578658174687e-08
+    1.094842569893916e-07
+    4.250139309046217e-07
+    3.574031946480214e-08
+    5.970174632295043e-08
+    1.695498154082625e-07
+    4.312932663600727e-07
+ 3.55e+10    
+    4.309480955892915e-07
+    1.695710437126253e-07
+    4.251426831385876e-07
+    5.972754826405484e-08
+    1.095399862423431e-07
+    4.250939405614726e-07
+    3.574854918798281e-08
+    5.973359811571741e-08
+     1.69626218360062e-07
+    4.313929186222446e-07
+ 3.56e+10    
+    4.310479869067949e-07
+    1.696474517137167e-07
+    4.252227472265429e-07
+    5.975919857573507e-08
+    1.095957170546301e-07
+    4.251740733712443e-07
+    3.575658489762147e-08
+    5.976533899103277e-08
+      1.6970270153231e-07
+    4.314927623150968e-07
+ 3.57e+10    
+    4.311480702040503e-07
+    1.697239395435971e-07
+    4.253029343626314e-07
+    5.979073749044724e-08
+    1.096514493179589e-07
+    4.252543293536068e-07
+    3.576442680533463e-08
+    5.979696892194772e-08
+     1.69779264877275e-07
+    4.315927976125906e-07
+ 3.58e+10    
+    4.312483456508653e-07
+    1.698005071504273e-07
+    4.253832445627983e-07
+    5.982216497893233e-08
+    1.097071829235276e-07
+    4.253347085269772e-07
+    3.577207512078968e-08
+    5.982848787859759e-08
+    1.698559083439598e-07
+    4.316930246860376e-07
+ 3.59e+10    
+    4.313488134144552e-07
+    1.698771544791464e-07
+    4.254636778418596e-07
+    5.985348100903814e-08
+    1.097629177620519e-07
+    4.254152109085363e-07
+    3.577953005171068e-08
+    5.985989582822793e-08
+    1.699326318781334e-07
+    4.317934437041246e-07
+ 3.6e+10     
+    4.314494736594725e-07
+    1.699538814715028e-07
+    4.255442342135185e-07
+    5.988468554574599e-08
+    1.098186537237898e-07
+     4.25495836514252e-07
+    3.578679180388527e-08
+    5.989119273522067e-08
+    1.700094354223629e-07
+    4.318940548329376e-07
+ 3.61e+10    
+    4.315503265480279e-07
+    1.700306880660854e-07
+    4.256249136903832e-07
+    5.991577855119704e-08
+     1.09874390698566e-07
+    4.255765853588982e-07
+    3.579386058117187e-08
+    5.992237856112057e-08
+    1.700863189160439e-07
+    4.319948582359855e-07
+ 3.62e+10    
+    4.316513722397152e-07
+    1.701075741983543e-07
+    4.257057162839883e-07
+    5.994675998471928e-08
+    1.099301285757961e-07
+    4.256574574560763e-07
+    3.580073658550804e-08
+    5.995345326466243e-08
+    1.701632822954327e-07
+     4.32095854074226e-07
+ 3.63e+10    
+    4.317526108916344e-07
+    1.701845398006712e-07
+    4.257866420048099e-07
+    5.997762980285465e-08
+    1.099858672445107e-07
+    4.257384528182326e-07
+     3.58074200169193e-08
+    5.998441680179798e-08
+    1.702403254936757e-07
+    4.321970425060883e-07
+ 3.64e+10    
+    4.318540426584178e-07
+    1.702615848023308e-07
+    4.258676908622851e-07
+    6.000838795938678e-08
+    1.100416065933781e-07
+    4.258195714566803e-07
+    3.581391107352879e-08
+    6.001526912572351e-08
+    1.703174484408405e-07
+    4.322984236874973e-07
+ 3.65e+10    
+     4.31955667692249e-07
+    1.703387091295883e-07
+     4.25948862864827e-07
+    6.003903440536847e-08
+    1.100973465107277e-07
+    4.259008133816175e-07
+    3.582020995156748e-08
+     6.00460101869076e-08
+    1.703946510639466e-07
+    4.323999977718977e-07
+ 3.66e+10    
+    4.320574861428912e-07
+    1.704159127056921e-07
+    4.260301580198465e-07
+    6.006956908915001e-08
+    1.101530868845727e-07
+    4.259821786021453e-07
+    3.582631684538532e-08
+    6.007663993311933e-08
+    1.704719332869941e-07
+    4.325017649102772e-07
+ 3.67e+10    
+    4.321594981577071e-07
+    1.704931954509111e-07
+    4.261115763337633e-07
+    6.009999195640744e-08
+    1.102088276026322e-07
+    4.260636671262889e-07
+    3.583223194746272e-08
+    6.010715830945639e-08
+    1.705492950309948e-07
+    4.326037252511917e-07
+ 3.68e+10    
+    4.322617038816828e-07
+    1.705705572825653e-07
+    4.261931178120283e-07
+    6.013030295017106e-08
+     1.10264568552353e-07
+    4.261452789610126e-07
+     3.58379554484229e-08
+    6.013756525837376e-08
+    1.706267362140007e-07
+    4.327058789407849e-07
+ 3.69e+10    
+    4.323641034574509e-07
+    1.706479981150541e-07
+     4.26274782459136e-07
+    6.016050201085446e-08
+    1.103203096209313e-07
+    4.262270141122414e-07
+    3.584348753704497e-08
+    6.016786071971251e-08
+    1.707042567511339e-07
+    4.328082261228159e-07
+ 3.7e+10     
+    4.324666970253127e-07
+    1.707255178598856e-07
+    4.263565702786424e-07
+    6.019058907628345e-08
+    1.103760506953341e-07
+    4.263088725848762e-07
+    3.584882840027732e-08
+      6.0198044630729e-08
+    1.707818565546148e-07
+    4.329107669386783e-07
+ 3.71e+10    
+    4.325694847232612e-07
+    1.708031164257048e-07
+    4.264384812731817e-07
+    6.022056408172537e-08
+    1.104317916623199e-07
+    4.263908543828129e-07
+    3.585397822325198e-08
+    6.022811692612397e-08
+    1.708595355337919e-07
+    4.330135015274265e-07
+ 3.72e+10    
+    4.326724666870044e-07
+    1.708807937183221e-07
+     4.26520515444481e-07
+    6.025042695991889e-08
+    1.104875324084593e-07
+    4.264729595089605e-07
+    3.585893718929932e-08
+    6.025807753807222e-08
+    1.709372935951695e-07
+    4.331164300257957e-07
+ 3.73e+10    
+    4.327756430499847e-07
+    1.709585496407413e-07
+    4.266026727933759e-07
+    6.028017764110336e-08
+    1.105432728201554e-07
+    4.265551879652549e-07
+    3.586370547996351e-08
+    6.028792639625227e-08
+    1.710151306424361e-07
+    4.332195525682253e-07
+ 3.74e+10    
+    4.328790139434045e-07
+    1.710363840931877e-07
+     4.26684953319828e-07
+    6.030981605304923e-08
+    1.105990127836635e-07
+    4.266375397526806e-07
+    3.586828327501853e-08
+     6.03176634278763e-08
+    1.710930465764926e-07
+    4.333228692868816e-07
+ 3.75e+10    
+    4.329825794962459e-07
+    1.711142969731353e-07
+    4.267673570229361e-07
+    6.033934212108788e-08
+     1.10654752185111e-07
+    4.267200148712841e-07
+    3.587267075248472e-08
+    6.034728855772038e-08
+    1.711710412954801e-07
+    4.334263803116811e-07
+ 3.76e+10    
+    4.330863398352931e-07
+    1.711922881753349e-07
+    4.268498839009557e-07
+    6.036875576814206e-08
+    1.107104909105167e-07
+    4.268026133201908e-07
+    3.587686808864586e-08
+    6.037680170815473e-08
+    1.712491146948076e-07
+    4.335300857703098e-07
+ 3.77e+10    
+    4.331902950851539e-07
+    1.712703575918403e-07
+    4.269325339513117e-07
+    6.039805691475665e-08
+    1.107662288458098e-07
+    4.268853350976226e-07
+    3.588087545806691e-08
+    6.040620279917423e-08
+    1.713272666671787e-07
+    4.336339857882477e-07
+ 3.78e+10    
+    4.332944453682814e-07
+    1.713485051120358e-07
+     4.27015307170611e-07
+    6.042724547912896e-08
+    1.108219658768485e-07
+    4.269681802009134e-07
+     3.58846930336122e-08
+    6.043549174842915e-08
+    1.714054971026196e-07
+    4.337380804887897e-07
+ 3.79e+10    
+    4.333987908049962e-07
+    1.714267306226633e-07
+    4.270982035546615e-07
+    6.045632137714016e-08
+    1.108777018894389e-07
+    4.270511486265244e-07
+    3.588832098646426e-08
+    6.046466847125602e-08
+    1.714838058885054e-07
+    4.338423699930672e-07
+ 3.8e+10     
+    4.335033315135059e-07
+    1.715050340078476e-07
+    4.271812230984821e-07
+     6.04852845223859e-08
+    1.109334367693527e-07
+    4.271342403700601e-07
+     3.58917594861429e-08
+    6.049373288070855e-08
+    1.715621929095867e-07
+    4.339468544200694e-07
+ 3.81e+10    
+    4.336080676099266e-07
+    1.715834151491242e-07
+    4.272643657963209e-07
+    6.051413482620768e-08
+    1.109891704023456e-07
+    4.272174554262846e-07
+    3.589500870052525e-08
+    6.052268488758909e-08
+    1.716406580480165e-07
+    4.340515338866658e-07
+ 3.82e+10    
+    4.337129992083059e-07
+    1.716618739254643e-07
+    4.273476316416653e-07
+    6.054287219772422e-08
+    1.110449026741744e-07
+    4.273007937891355e-07
+    3.589806879586577e-08
+    6.055152440047954e-08
+     1.71719201183376e-07
+     4.34156408507626e-07
+ 3.83e+10    
+    4.338181264206411e-07
+    1.717404102133003e-07
+    4.274310206272569e-07
+    6.057149654386305e-08
+    1.111006334706152e-07
+      4.2738425545174e-07
+    3.590093993681724e-08
+    6.058025132577313e-08
+    1.717978221927005e-07
+     4.34261478395641e-07
+ 3.84e+10    
+    4.339234493569009e-07
+     1.71819023886553e-07
+    4.275145327451075e-07
+    6.060000776939204e-08
+    1.111563626774798e-07
+      4.2746784040643e-07
+    3.590362228645198e-08
+    6.060886556770607e-08
+    1.718765209505058e-07
+    4.343667436613464e-07
+ 3.85e+10    
+    4.340289681250454e-07
+    1.718977148166548e-07
+    4.275981679865093e-07
+    6.062840577695111e-08
+    1.112120901806327e-07
+    4.275515486447565e-07
+    3.590611600628335e-08
+    6.063736702838902e-08
+    1.719552973288131e-07
+    4.344722044133395e-07
+ 3.86e+10    
+     4.34134682831048e-07
+    1.719764828725772e-07
+    4.276819263420486e-07
+    6.065669046708427e-08
+    1.112678158660081e-07
+    4.276353801575023e-07
+    3.590842125628822e-08
+    6.066575560783903e-08
+    1.720341511971742e-07
+    4.345778607582031e-07
+ 3.87e+10    
+    4.342405935789142e-07
+    1.720553279208539e-07
+    4.277658078016224e-07
+    6.068486173827167e-08
+    1.113235396196262e-07
+    4.277193349347006e-07
+    3.591053819492941e-08
+    6.069403120401176e-08
+    1.721130824226974e-07
+    4.346837128005235e-07
+ 3.88e+10    
+    4.343467004707015e-07
+    1.721342498256063e-07
+    4.278498123544466e-07
+    6.071291948696146e-08
+    1.113792613276087e-07
+    4.278034129656444e-07
+    3.591246697917884e-08
+    6.072219371283317e-08
+    1.721920908700716e-07
+    4.347897606429141e-07
+ 3.89e+10    
+    4.344530036065405e-07
+    1.722132484485682e-07
+    4.279339399890717e-07
+     6.07408636076024e-08
+    1.114349808761957e-07
+    4.278876142389054e-07
+      3.5914207764541e-08
+    6.075024302823209e-08
+    1.722711764015915e-07
+    4.348960043860321e-07
+ 3.9e+10     
+    4.345595030846539e-07
+    1.722923236491096e-07
+    4.280181906933945e-07
+    6.076869399267577e-08
+    1.114906981517607e-07
+    4.279719387423431e-07
+    3.591576070507685e-08
+    6.077817904217217e-08
+    1.723503388771818e-07
+    4.350024441286017e-07
+ 3.91e+10    
+    4.346661990013761e-07
+    1.723714752842614e-07
+    4.281025644546713e-07
+    6.079641053272818e-08
+    1.115464130408264e-07
+    4.280563864631214e-07
+    3.591712595342824e-08
+    6.080600164468457e-08
+    1.724295781544214e-07
+    4.351090799674312e-07
+ 3.92e+10    
+    4.347730914511742e-07
+     1.72450703208739e-07
+    4.281870612595294e-07
+    6.082401311640387e-08
+    1.116021254300797e-07
+    4.281409573877223e-07
+    3.591830366084258e-08
+    6.083371072390012e-08
+    1.725088940885677e-07
+    4.352159119974357e-07
+ 3.93e+10    
+    4.348801805266652e-07
+    1.725300072749662e-07
+    4.282716810939801e-07
+     6.08515016304774e-08
+    1.116578352063867e-07
+    4.282256515019581e-07
+    3.591929397719803e-08
+    6.086130616608219e-08
+    1.725882865325803e-07
+    4.353229403116544e-07
+ 3.94e+10    
+    4.349874663186368e-07
+    1.726093873330979e-07
+    4.283564239434298e-07
+    6.087887595988611e-08
+    1.117135422568076e-07
+    4.283104687909841e-07
+    3.592009705102891e-08
+    6.088878785565903e-08
+    1.726677553371447e-07
+     4.35430165001272e-07
+ 3.95e+10    
+    4.350949489160661e-07
+    1.726888432310448e-07
+    4.284412897926941e-07
+    6.090613598776324e-08
+    1.117692464686115e-07
+    4.283954092393143e-07
+    3.592071302955175e-08
+     6.09161556752567e-08
+    1.727473003506955e-07
+    4.355375861556368e-07
+ 3.96e+10    
+    4.352026284061382e-07
+    1.727683748144955e-07
+     4.28526278626006e-07
+     6.09332815954705e-08
+    1.118249477292905e-07
+    4.284804728308316e-07
+    3.592114205869152e-08
+    6.094340950573166e-08
+    1.728269214194401e-07
+    4.356452038622816e-07
+ 3.97e+10    
+    4.353105048742663e-07
+    1.728479819269392e-07
+    4.286113904270316e-07
+    6.096031266263088e-08
+    1.118806459265735e-07
+    4.285656595488011e-07
+    3.592138428310817e-08
+    6.097054922620374e-08
+    1.729066183873811e-07
+    4.357530182069403e-07
+ 3.98e+10    
+    4.354185784041085e-07
+    1.729276644096895e-07
+    4.286966251788788e-07
+    6.098722906716176e-08
+    1.119363409484411e-07
+    4.286509693758841e-07
+    3.592143984622373e-08
+    6.099757471408887e-08
+    1.729863910963397e-07
+      4.3586102927357e-07
+ 3.99e+10    
+    4.355268490775891e-07
+    1.730074221019061e-07
+    4.287819828641107e-07
+    6.101403068530792e-08
+    1.119920326831386e-07
+    4.287364022941502e-07
+    3.592130889024964e-08
+    6.102448584513221e-08
+    1.730662393859781e-07
+    4.359692371443673e-07
+ 4e+10       
+    4.356353169749146e-07
+     1.73087254840617e-07
+    4.288674634647542e-07
+    6.104071739167439e-08
+    1.120477210191898e-07
+    4.288219582850884e-07
+    3.592099155621433e-08
+    6.105128249344097e-08
+    1.731461630938217e-07
+    4.360776418997881e-07
+ 4.01e+10    
+    4.357439821745933e-07
+     1.73167162460741e-07
+     4.28953066962315e-07
+     6.10672890592597e-08
+    1.121034058454106e-07
+    4.289076373296205e-07
+    3.592048798399133e-08
+     6.10779645315176e-08
+     1.73226162055282e-07
+    4.361862436185685e-07
+ 4.02e+10    
+    4.358528447534529e-07
+    1.732471447951098e-07
+    4.290387933377859e-07
+    6.109374555948887e-08
+    1.121590870509218e-07
+    4.289934394081126e-07
+    3.591979831232747e-08
+    6.110453183029263e-08
+    1.733062361036776e-07
+    4.362950423777387e-07
+ 4.03e+10    
+    4.359619047866602e-07
+    1.733272016744893e-07
+    4.291246425716585e-07
+    6.112008676224676e-08
+    1.122147645251625e-07
+    4.290793645003875e-07
+    3.591892267887169e-08
+    6.113098425915804e-08
+    1.733863850702574e-07
+    4.364040382526449e-07
+ 4.04e+10    
+    4.360711623477359e-07
+    1.734073329276011e-07
+    4.292106146439339e-07
+    6.114631253591099e-08
+    1.122704381579028e-07
+    4.291654125857366e-07
+    3.591786122020377e-08
+    6.115732168600015e-08
+     1.73466608784221e-07
+    4.365132313169672e-07
+ 4.05e+10    
+    4.361806175085762e-07
+    1.734875383811443e-07
+     4.29296709534134e-07
+    6.117242274738539e-08
+    1.123261078392562e-07
+    4.292515836429303e-07
+    3.591661407186372e-08
+    6.118354397723295e-08
+    1.735469070727406e-07
+    4.366226216427359e-07
+ 4.06e+10    
+    4.362902703394683e-07
+    1.735678178598162e-07
+    4.293829272213112e-07
+    6.119841726213312e-08
+    1.123817734596926e-07
+    4.293378776502323e-07
+    3.591518136838128e-08
+    6.120965099783117e-08
+    1.736272797609831e-07
+    4.367322093003517e-07
+ 4.07e+10    
+     4.36400120909108e-07
+    1.736481711863341e-07
+    4.294692676840602e-07
+    6.122429594420992e-08
+    1.124374349100501e-07
+    4.294242945854077e-07
+     3.59135632433057e-08
+    6.123564261136361e-08
+    1.737077266721297e-07
+    4.368419943586023e-07
+ 4.08e+10    
+    4.365101692846178e-07
+    1.737285981814545e-07
+    4.295557309005267e-07
+    6.125005865629731e-08
+    1.124930920815473e-07
+     4.29510834425736e-07
+     3.59117598292358e-08
+    6.126151868002609e-08
+    1.737882476273977e-07
+    4.369519768846799e-07
+ 4.09e+10    
+    4.366204155315641e-07
+    1.738090986639958e-07
+    4.296423168484202e-07
+    6.127570525973614e-08
+    1.125487448657959e-07
+    4.295974971480238e-07
+    3.590977125785048e-08
+    6.128727906467503e-08
+    1.738688424460618e-07
+    4.370621569442009e-07
+ 4.1e+10     
+    4.367308597139756e-07
+    1.738896724508573e-07
+    4.297290255050215e-07
+    6.130123561455964e-08
+    1.126043931548113e-07
+    4.296842827286133e-07
+    3.590759765993918e-08
+    6.131292362486041e-08
+    1.739495109454732e-07
+    4.371725346012217e-07
+ 4.11e+10    
+    4.368415018943575e-07
+    1.739703193570394e-07
+     4.29815856847193e-07
+    6.132664957952659e-08
+    1.126600368410251e-07
+    4.297711911433932e-07
+    3.590523916543275e-08
+    6.133845221885894e-08
+    1.740302529410809e-07
+    4.372831099182543e-07
+ 4.12e+10    
+    4.369523421337113e-07
+    1.740510391956649e-07
+    4.299028108513922e-07
+    6.135194701215491e-08
+    1.127156758172967e-07
+    4.298582223678126e-07
+    3.590269590343472e-08
+    6.136386470370758e-08
+    1.741110682464518e-07
+    4.373938829562886e-07
+ 4.13e+10    
+    4.370633804915497e-07
+    1.741318317779977e-07
+    4.299898874936777e-07
+    6.137712776875476e-08
+    1.127713099769241e-07
+     4.29945376376888e-07
+    3.589996800225252e-08
+    6.138916093523651e-08
+    1.741919566732905e-07
+    4.375048537748038e-07
+ 4.14e+10    
+    4.371746170259163e-07
+    1.742126969134631e-07
+    4.300770867497195e-07
+    6.140219170446184e-08
+    1.128269392136555e-07
+     4.30032653145217e-07
+    3.589705558942915e-08
+    6.141434076810243e-08
+    1.742729180314595e-07
+    4.376160224317908e-07
+ 4.15e+10    
+    4.372860517933976e-07
+    1.742936344096667e-07
+    4.301644085948099e-07
+    6.142713867327062e-08
+    1.128825634216999e-07
+     4.30120052646987e-07
+    3.589395879177496e-08
+    6.143940405582172e-08
+    1.743539521289983e-07
+    4.377273889837652e-07
+ 4.16e+10    
+    4.373976848491445e-07
+    1.743746440724153e-07
+    4.302518530038744e-07
+    6.145196852806763e-08
+    1.129381824957387e-07
+    4.302075748559854e-07
+    3.589067773539974e-08
+    6.146435065080368e-08
+     1.74435058772143e-07
+    4.378389534857859e-07
+ 4.17e+10    
+    4.375095162468843e-07
+    1.744557257057343e-07
+    4.303394199514772e-07
+    6.147668112066464e-08
+    1.129937963309358e-07
+    4.302952197456117e-07
+    3.588721254574487e-08
+    6.148918040438358e-08
+    1.745162377653461e-07
+    4.379507159914702e-07
+ 4.18e+10    
+    4.376215460389412e-07
+    1.745368791118879e-07
+    4.304271094118345e-07
+    6.150127630183198e-08
+    1.130494048229485e-07
+    4.303829872888856e-07
+    3.588356334761594e-08
+    6.151389316685593e-08
+     1.74597488911295e-07
+    4.380626765530131e-07
+ 4.19e+10    
+    4.377337742762477e-07
+    1.746181040913974e-07
+     4.30514921358821e-07
+    6.152575392133142e-08
+    1.131050078679379e-07
+     4.30470877458458e-07
+    3.587973026521525e-08
+    6.153848878750748e-08
+    1.746788120109315e-07
+    4.381748352212017e-07
+ 4.2e+10     
+    4.378462010083655e-07
+    1.746994004430603e-07
+    4.306028557659817e-07
+    6.155011382794962e-08
+    1.131606053625792e-07
+    4.305588902266219e-07
+    3.587571342217482e-08
+    6.156296711465042e-08
+    1.747602068634699e-07
+    4.382871920454307e-07
+ 4.21e+10    
+    4.379588262834983e-07
+    1.747807679639685e-07
+    4.306909126065385e-07
+    6.157435586953117e-08
+    1.132161972040721e-07
+    4.306470255653206e-07
+    3.587151294158926e-08
+    6.158732799565516e-08
+    1.748416732664165e-07
+    4.383997470737214e-07
+ 4.22e+10    
+    4.380716501485085e-07
+    1.748622064495272e-07
+    4.307790918534013e-07
+    6.159847989301159e-08
+    1.132717832901505e-07
+    4.307352834461579e-07
+    3.586712894604915e-08
+    6.161157127698379e-08
+    1.749232110155872e-07
+    4.385125003527351e-07
+ 4.23e+10    
+    4.381846726489315e-07
+    1.749437156934719e-07
+    4.308673934791752e-07
+    6.162248574445032e-08
+    1.133273635190929e-07
+    4.308236638404089e-07
+    3.586256155767431e-08
+    6.163569680422261e-08
+    1.750048199051264e-07
+    4.386254519277909e-07
+ 4.24e+10    
+     4.38297893828995e-07
+    1.750252954878879e-07
+    4.309558174561712e-07
+    6.164637326906387e-08
+    1.133829377897316e-07
+     4.30912166719028e-07
+    3.585781089814746e-08
+     6.16597044221153e-08
+    1.750864997275246e-07
+    4.387386018428802e-07
+ 4.25e+10    
+    4.384113137316314e-07
+    1.751069456232277e-07
+    4.310443637564133e-07
+    6.167014231125878e-08
+     1.13438506001463e-07
+    4.310007920526598e-07
+     3.58528770887479e-08
+    6.168359397459578e-08
+    1.751682502736371e-07
+     4.38851950140684e-07
+ 4.26e+10    
+    4.385249323984924e-07
+    1.751886658883279e-07
+    4.311330323516487e-07
+    6.169379271466431e-08
+    1.134940680542567e-07
+    4.310895398116476e-07
+    3.584776025038538e-08
+    6.170736530482094e-08
+    1.752500713327008e-07
+    4.389654968625864e-07
+ 4.27e+10    
+    4.386387498699675e-07
+    1.752704560704275e-07
+    4.312218232133544e-07
+    6.171732432216545e-08
+    1.135496238486652e-07
+    4.311784099660423e-07
+    3.584246050363414e-08
+     6.17310182552036e-08
+    1.753319626923527e-07
+    4.390792420486924e-07
+ 4.28e+10    
+    4.387527661851968e-07
+    1.753523159551861e-07
+    4.313107363127493e-07
+    6.174073697593588e-08
+    1.136051732858332e-07
+    4.312674024856131e-07
+    3.583697796876717e-08
+    6.175455266744516e-08
+     1.75413924138647e-07
+    4.391931857378409e-07
+ 4.29e+10    
+    4.388669813820867e-07
+    1.754342453266988e-07
+    4.313997716207973e-07
+    6.176403051747028e-08
+    1.136607162675063e-07
+    4.313565173398547e-07
+     3.58313127657903e-08
+     6.17779683825681e-08
+    1.754959554560723e-07
+     4.39307327967623e-07
+ 4.3e+10     
+    4.389813954973243e-07
+     1.75516243967516e-07
+    4.314889291082212e-07
+    6.178720478761745e-08
+    1.137162526960407e-07
+    4.314457544979979e-07
+    3.582546501447689e-08
+    6.180126524094896e-08
+    1.755780564275689e-07
+    4.394216687743935e-07
+ 4.31e+10    
+    4.390960085663926e-07
+    1.755983116586583e-07
+    4.315782087455078e-07
+    6.181025962661268e-08
+    1.137717824744121e-07
+    4.315351139290174e-07
+    3.581943483440223e-08
+    6.182444308235056e-08
+    1.756602268345457e-07
+    4.395362081932891e-07
+ 4.32e+10    
+    4.392108206235857e-07
+     1.75680448179634e-07
+    4.316676105029167e-07
+    6.183319487411048e-08
+    1.138273055062241e-07
+    4.316245956016423e-07
+    3.581322234497836e-08
+    6.184750174595484e-08
+     1.75742466456898e-07
+    4.396509462582429e-07
+ 4.33e+10    
+    4.393258317020223e-07
+    1.757626533084565e-07
+     4.31757134350488e-07
+     6.18560103692169e-08
+    1.138828216957173e-07
+    4.317141994843618e-07
+    3.580682766548868e-08
+    6.187044107039479e-08
+    1.758247750730218e-07
+    4.397658830019964e-07
+ 4.34e+10    
+    4.394410418336612e-07
+    1.758449268216589e-07
+    4.318467802580523e-07
+    6.187870595052205e-08
+    1.139383309477777e-07
+    4.318039255454376e-07
+    3.580025091512304e-08
+    6.189326089378727e-08
+     1.75907152459833e-07
+    4.398810184561173e-07
+ 4.35e+10    
+    4.395564510493149e-07
+    1.759272684943124e-07
+    4.319365481952363e-07
+    6.190128145613252e-08
+    1.139938331679455e-07
+     4.31893773752909e-07
+    3.579349221301275e-08
+    6.191596105376515e-08
+    1.759895983927824e-07
+    4.399963526510139e-07
+ 4.36e+10    
+    4.396720593786644e-07
+     1.76009678100041e-07
+    4.320264381314724e-07
+    6.192373672370354e-08
+    1.140493282624233e-07
+    4.319837440746039e-07
+    3.578655167826549e-08
+    6.193854138750942e-08
+     1.76072112645872e-07
+    4.401118856159479e-07
+ 4.37e+10    
+    4.397878668502735e-07
+     1.76092155411038e-07
+    4.321164500360051e-07
+     6.19460715904712e-08
+    1.141048161380843e-07
+    4.320738364781463e-07
+    3.577942943000068e-08
+    6.196100173178135e-08
+    1.761546949916714e-07
+    4.402276173790493e-07
+ 4.38e+10    
+     4.39903873491601e-07
+    1.761747001980822e-07
+    4.322065838779007e-07
+    6.196828589328467e-08
+    1.141602967024806e-07
+    4.321640509309631e-07
+    3.577212558738475e-08
+    6.198334192295471e-08
+    1.762373452013335e-07
+    4.403435479673322e-07
+ 4.39e+10    
+    4.400200793290173e-07
+    1.762573122305527e-07
+    4.322968396260524e-07
+    6.199037946863806e-08
+    1.142157698638515e-07
+    4.322543874002954e-07
+    3.576464026966641e-08
+    6.200556179704746e-08
+    1.763200630446103e-07
+    4.404596774067073e-07
+ 4.4e+10     
+    4.401364843878177e-07
+    1.763399912764459e-07
+    4.323872172491909e-07
+    6.201235215270277e-08
+    1.142712355311315e-07
+    4.323448458532053e-07
+    3.575697359621223e-08
+    6.202766118975395e-08
+    1.764028482898689e-07
+    4.405760057219968e-07
+ 4.41e+10    
+    4.402530886922338e-07
+    1.764227371023897e-07
+    4.324777167158895e-07
+    6.203420378135869e-08
+    1.143266936139574e-07
+    4.324354262565817e-07
+    3.574912568654196e-08
+    6.204963993647643e-08
+    1.764857007041065e-07
+    4.406925329369479e-07
+ 4.42e+10    
+      4.4036989226545e-07
+    1.765055494736591e-07
+    4.325683379945724e-07
+    6.205593419022671e-08
+    1.143821440226774e-07
+    4.325261285771521e-07
+    3.574109666036419e-08
+    6.207149787235692e-08
+    1.765686200529658e-07
+    4.408092590742465e-07
+ 4.43e+10    
+    4.404868951296149e-07
+    1.765884281541915e-07
+    4.326590810535231e-07
+    6.207754321469987e-08
+    1.144375866683576e-07
+    4.326169527814876e-07
+    3.573288663761204e-08
+    6.209323483230886e-08
+    1.766516061007507e-07
+     4.40926184155532e-07
+ 4.44e+10    
+    4.406040973058567e-07
+    1.766713729066022e-07
+    4.327499458608895e-07
+    6.209903068997534e-08
+    1.144930214627905e-07
+    4.327078988360127e-07
+    3.572449573847873e-08
+    6.211485065104856e-08
+    1.767346586104409e-07
+    4.410433082014099e-07
+ 4.45e+10    
+    4.407214988142936e-07
+    1.767543834921982e-07
+    4.328409323846938e-07
+    6.212039645108561e-08
+     1.14548448318502e-07
+    4.327989667070117e-07
+    3.571592408345327e-08
+    6.213634516312658e-08
+    1.768177773437068e-07
+    4.411606312314661e-07
+ 4.46e+10    
+    4.408390996740508e-07
+    1.768374596709936e-07
+    4.329320405928376e-07
+    6.214164033293012e-08
+     1.14603867148759e-07
+     4.32890156360637e-07
+    3.570717179335638e-08
+    6.215771820295921e-08
+    1.769009620609246e-07
+    4.412781532642794e-07
+ 4.47e+10    
+    4.409568999032706e-07
+    1.769206012017241e-07
+    4.330232704531098e-07
+    6.216276217030648e-08
+    1.146592778675765e-07
+    4.329814677629154e-07
+     3.56982389893761e-08
+    6.217896960485953e-08
+    1.769842125211908e-07
+    4.413958743174351e-07
+ 4.48e+10    
+    4.410748995191272e-07
+    1.770038078418615e-07
+    4.331146219331951e-07
+    6.218376179794171e-08
+    1.147146803897255e-07
+    4.330729008797589e-07
+    3.568912579310379e-08
+    6.220009920306882e-08
+    1.770675284823365e-07
+    4.415137944075397e-07
+ 4.49e+10    
+    4.411930985378372e-07
+     1.77087079347628e-07
+    4.332060950006779e-07
+    6.220463905052323e-08
+    1.147700746307393e-07
+    4.331644556769686e-07
+    3.567983232656981e-08
+    6.222110683178723e-08
+     1.77150909700942e-07
+    4.416319135502318e-07
+ 4.5e+10     
+    4.413114969746762e-07
+    1.771704154740103e-07
+    4.332976896230515e-07
+    6.222539376273009e-08
+    1.148254605069211e-07
+    4.332561321202439e-07
+    3.567035871227955e-08
+    6.224199232520495e-08
+    1.772343559323512e-07
+     4.41750231760196e-07
+ 4.51e+10    
+    4.414300948439871e-07
+    1.772538159747736e-07
+    4.333894057677248e-07
+    6.224602576926357e-08
+     1.14880837935351e-07
+    4.333479301751889e-07
+    3.566070507324919e-08
+    6.226275551753294e-08
+    1.773178669306851e-07
+    4.418687490511774e-07
+ 4.52e+10    
+    4.415488921591964e-07
+    1.773372806024755e-07
+    4.334812434020283e-07
+    6.226653490487803e-08
+    1.149362068338924e-07
+    4.334398498073205e-07
+    3.565087153304165e-08
+    6.228339624303367e-08
+    1.774014424488565e-07
+     4.41987465435991e-07
+ 4.53e+10    
+    4.416678889328247e-07
+    1.774208091084802e-07
+    4.335732024932222e-07
+    6.228692100441195e-08
+    1.149915671211998e-07
+    4.335318909820762e-07
+    3.564085821580252e-08
+    6.230391433605169e-08
+    1.774850822385832e-07
+    4.421063809265378e-07
+ 4.54e+10    
+    4.417870851764989e-07
+    1.775044012429717e-07
+    4.336652830085006e-07
+    6.230718390281785e-08
+    1.150469187167243e-07
+     4.33624053664818e-07
+    3.563066524629585e-08
+      6.2324309631044e-08
+    1.775687860504021e-07
+    4.422254955338153e-07
+ 4.55e+10    
+    4.419064809009677e-07
+    1.775880567549674e-07
+    4.337574849150009e-07
+    6.232732343519327e-08
+     1.15102261540721e-07
+    4.337163378208434e-07
+    3.562029274994017e-08
+    6.234458196261071e-08
+    1.776525536336824e-07
+    4.423448092679306e-07
+ 4.56e+10    
+    4.420260761161075e-07
+    1.776717753923318e-07
+    4.338498081798093e-07
+    6.234733943681072e-08
+    1.151575955142556e-07
+    4.338087434153898e-07
+    3.560974085284426e-08
+     6.23647311655249e-08
+    1.777363847366396e-07
+    4.424643221381137e-07
+ 4.57e+10    
+    4.421458708309419e-07
+    1.777555569017892e-07
+    4.339422527699656e-07
+    6.236723174314812e-08
+    1.152129205592108e-07
+    4.339012704136423e-07
+     3.55990096818431e-08
+    6.238475707476305e-08
+    1.778202791063483e-07
+    4.425840341527285e-07
+ 4.58e+10    
+    4.422658650536478e-07
+    1.778394010289374e-07
+    4.340348186524728e-07
+    6.238700018991871e-08
+    1.152682365982923e-07
+    4.339939187807402e-07
+    3.558809936453365e-08
+    6.240465952553492e-08
+    1.779042364887557e-07
+    4.427039453192851e-07
+ 4.59e+10    
+    4.423860587915701e-07
+    1.779233075182603e-07
+    4.341275057943011e-07
+    6.240664461310119e-08
+    1.153235435550358e-07
+    4.340866884817842e-07
+    3.557701002931065e-08
+    6.242443835331335e-08
+    1.779882566286939e-07
+    4.428240556444528e-07
+ 4.6e+10     
+    4.425064520512328e-07
+    1.780072761131411e-07
+    4.342203141623953e-07
+    6.242616484896926e-08
+    1.153788413538128e-07
+    4.341795794818417e-07
+    3.556574180540245e-08
+    6.244409339386423e-08
+    1.780723392698942e-07
+    4.429443651340719e-07
+ 4.61e+10    
+    4.426270448383521e-07
+    1.780913065558751e-07
+    4.343132437236807e-07
+    6.244556073412168e-08
+    1.154341299198368e-07
+    4.342725917459558e-07
+    3.555429482290675e-08
+    6.246362448327594e-08
+    1.781564841549986e-07
+     4.43064873793165e-07
+ 4.62e+10    
+    4.427478371578454e-07
+    1.781753985876818e-07
+     4.34406294445068e-07
+    6.246483210551156e-08
+      1.1548940917917e-07
+    4.343657252391504e-07
+    3.554266921282627e-08
+    6.248303145798879e-08
+    1.782406910255733e-07
+    4.431855816259485e-07
+ 4.63e+10    
+    4.428688290138457e-07
+    1.782595519487178e-07
+    4.344994662934631e-07
+    6.248397880047592e-08
+    1.155446790587285e-07
+    4.344589799264358e-07
+    3.553086510710446e-08
+    6.250231415482473e-08
+    1.783249596221205e-07
+    4.433064886358467e-07
+ 4.64e+10    
+    4.429900204097089e-07
+    1.783437663780896e-07
+    4.345927592357682e-07
+    6.250300065676493e-08
+    1.155999394862886e-07
+     4.34552355772816e-07
+    3.551888263866096e-08
+    6.252147241101612e-08
+    1.784092896840916e-07
+    4.434275948254991e-07
+ 4.65e+10    
+    4.431114113480305e-07
+    1.784280416138649e-07
+    4.346861732388928e-07
+    6.252189751257121e-08
+    1.156551903904931e-07
+    4.346458527432967e-07
+    3.550672194142739e-08
+    6.254050606423526e-08
+    1.784936809498991e-07
+    4.435489001967776e-07
+ 4.66e+10    
+     4.43233001830653e-07
+    1.785123773930858e-07
+    4.347797082697559e-07
+     6.25406692065588e-08
+    1.157104317008566e-07
+    4.347394708028887e-07
+    3.549438315038257e-08
+    6.255941495262302e-08
+    1.785781331569287e-07
+     4.43670404750792e-07
+ 4.67e+10    
+     4.43354791858678e-07
+    1.785967734517798e-07
+    4.348733642952932e-07
+    6.255931557789191e-08
+    1.157656633477712e-07
+    4.348332099166157e-07
+    3.548186640158815e-08
+    6.257819891481791e-08
+    1.786626460415518e-07
+    4.437921084879064e-07
+ 4.68e+10    
+    4.434767814324779e-07
+    1.786812295249726e-07
+    4.349671412824638e-07
+    6.257783646626402e-08
+    1.158208852625129e-07
+      4.3492707004952e-07
+    3.546917183222385e-08
+    6.259685778998459e-08
+    1.787472193391368e-07
+    4.439140114077462e-07
+ 4.69e+10    
+    4.435989705517054e-07
+    1.787657453466995e-07
+    4.350610391982551e-07
+    6.259623171192617e-08
+    1.158760973772467e-07
+    4.350210511666692e-07
+     3.54562995806227e-08
+    6.261539141784258e-08
+    1.788318527840613e-07
+    4.440361135092125e-07
+ 4.7e+10     
+    4.437213592153058e-07
+    1.788503206500169e-07
+    4.351550580096876e-07
+    6.261450115571562e-08
+    1.159312996250315e-07
+    4.351151532331613e-07
+    3.544324978630635e-08
+    6.263379963869442e-08
+    1.789165461097238e-07
+    4.441584147904914e-07
+ 4.71e+10    
+    4.438439474215278e-07
+    1.789349551670143e-07
+    4.352491976838228e-07
+    6.263264463908413e-08
+    1.159864919398272e-07
+    4.352093762141315e-07
+    3.543002259002007e-08
+     6.26520822934543e-08
+    1.790012990485555e-07
+    4.442809152490654e-07
+ 4.72e+10    
+    4.439667351679324e-07
+    1.790196486288253e-07
+    4.353434581877675e-07
+     6.26506620041262e-08
+    1.160416742564988e-07
+    4.353037200747588e-07
+    3.541661813376776e-08
+    6.267023922367579e-08
+    1.790861113320312e-07
+    4.444036148817242e-07
+ 4.73e+10    
+    4.440897224514056e-07
+    1.791044007656393e-07
+    4.354378394886789e-07
+    6.266855309360706e-08
+    1.160968465108221e-07
+    4.353981847802688e-07
+    3.540303656084697e-08
+    6.268827027158004e-08
+     1.79170982690681e-07
+    4.445265136845756e-07
+ 4.74e+10    
+    4.442129092681673e-07
+    1.791892113067125e-07
+    4.355323415537707e-07
+    6.268631775099047e-08
+    1.161520086394891e-07
+    4.354927702959424e-07
+    3.538927801588362e-08
+     6.27061752800836e-08
+    1.792559128541019e-07
+    4.446496116530568e-07
+ 4.75e+10    
+    4.443362956137825e-07
+     1.79274079980379e-07
+    4.356269643503198e-07
+    6.270395582046667e-08
+    1.162071605801134e-07
+     4.35587476587121e-07
+    3.537534264486666e-08
+    6.272395409282588e-08
+    1.793409015509677e-07
+    4.447729087819411e-07
+ 4.76e+10    
+    4.444598814831725e-07
+     1.79359006514062e-07
+    4.357217078456694e-07
+    6.272146714697992e-08
+    1.162623022712349e-07
+    4.356823036192117e-07
+     3.53612305951829e-08
+      6.2741606554197e-08
+    1.794259485090418e-07
+    4.448964050653557e-07
+ 4.77e+10    
+    4.445836668706218e-07
+    1.794439906342843e-07
+    4.358165720072354e-07
+     6.27388515762557e-08
+    1.163174336523253e-07
+    4.357772513576924e-07
+     3.53469420156512e-08
+    6.275913250936481e-08
+    1.795110534551866e-07
+    4.450201004967854e-07
+ 4.78e+10    
+    4.447076517697919e-07
+    1.795290320666797e-07
+    4.359115568025127e-07
+     6.27561089548283e-08
+    1.163725546637929e-07
+    4.358723197681192e-07
+    3.533247705655703e-08
+    6.277653180430237e-08
+     1.79596216115375e-07
+    4.451439950690857e-07
+ 4.79e+10    
+      4.4483183617373e-07
+    1.796141305360027e-07
+    4.360066621990777e-07
+    6.277323913006775e-08
+    1.164276652469877e-07
+     4.35967508816129e-07
+    3.531783586968668e-08
+    6.279380428581479e-08
+    1.796814362147009e-07
+    4.452680887744922e-07
+ 4.8e+10     
+    4.449562200748785e-07
+      1.7969928576614e-07
+    4.361018881645975e-07
+    6.279024195020694e-08
+    1.164827653442065e-07
+    4.360628184674478e-07
+    3.530301860836132e-08
+    6.281094980156622e-08
+    1.797667134773897e-07
+     4.45392381604632e-07
+ 4.81e+10    
+    4.450808034650846e-07
+    1.797844974801207e-07
+    4.361972346668313e-07
+    6.280711726436829e-08
+    1.165378548986972e-07
+    4.361582486878944e-07
+    3.528802542747107e-08
+    6.282796820010673e-08
+     1.79852047626809e-07
+    4.455168735505321e-07
+ 4.82e+10    
+    4.452055863356111e-07
+     1.79869765400126e-07
+    4.362927016736368e-07
+    6.282386492259037e-08
+    1.165929338546642e-07
+    4.362537994433869e-07
+    3.527285648350872e-08
+    6.284485933089857e-08
+    1.799374383854788e-07
+    4.456415646026305e-07
+ 4.83e+10    
+     4.45330568677146e-07
+    1.799550892475002e-07
+    4.363882891529775e-07
+    6.284048477585453e-08
+    1.166480021572728e-07
+    4.363494706999457e-07
+    3.525751193460351e-08
+    6.286162304434279e-08
+    1.800228854750815e-07
+    4.457664547507855e-07
+ 4.84e+10    
+    4.454557504798102e-07
+    1.800404687427606e-07
+    4.364839970729227e-07
+    6.285697667611117e-08
+    1.167030597526543e-07
+    4.364452624237021e-07
+    3.524199194055472e-08
+    6.287825919180554e-08
+    1.801083886164728e-07
+    4.458915439842851e-07
+ 4.85e+10    
+    4.455811317331707e-07
+    1.801259036056072e-07
+    4.365798254016579e-07
+     6.28733404763058e-08
+    1.167581065879098e-07
+    4.365411745809003e-07
+    3.522629666286494e-08
+    6.289476762564386e-08
+    1.801939475296905e-07
+    4.460168322918569e-07
+ 4.86e+10    
+    4.457067124262448e-07
+    1.802113935549332e-07
+    4.366757741074857e-07
+    6.288957603040513e-08
+    1.168131426111157e-07
+    4.366372071379041e-07
+    3.521042626477346e-08
+    6.291114819923202e-08
+    1.802795619339657e-07
+    4.461423196616789e-07
+ 4.87e+10    
+     4.45832492547515e-07
+    1.802969383088342e-07
+     4.36771843158832e-07
+    6.290568319342287e-08
+    1.168681677713276e-07
+    4.367333600612026e-07
+    3.519438091128924e-08
+     6.29274007669869e-08
+    1.803652315477318e-07
+    4.462680060813868e-07
+ 4.88e+10    
+    4.459584720849341e-07
+    1.803825375846182e-07
+    4.368680325242525e-07
+    6.292166182144533e-08
+    1.169231820185851e-07
+    4.368296333174122e-07
+    3.517816076922388e-08
+    6.294352518439377e-08
+    1.804509560886347e-07
+    4.463938915380845e-07
+ 4.89e+10    
+    4.460846510259362e-07
+    1.804681910988152e-07
+    4.369643421724339e-07
+    6.293751177165691e-08
+    1.169781853039158e-07
+    4.369260268732855e-07
+    3.516176600722438e-08
+    6.295952130803155e-08
+    1.805367352735419e-07
+    4.465199760183535e-07
+ 4.9e+10     
+    4.462110293574451e-07
+    1.805538985671871e-07
+    4.370607720722015e-07
+    6.295323290236552e-08
+    1.170331775793403e-07
+    4.370225406957136e-07
+    3.514519679580566e-08
+    6.297538899559825e-08
+    1.806225688185525e-07
+    4.466462595082626e-07
+ 4.91e+10    
+    4.463376070658829e-07
+    1.806396597047357e-07
+    4.371573221925225e-07
+    6.296882507302747e-08
+    1.170881587978759e-07
+    4.371191747517313e-07
+    3.512845330738297e-08
+    6.299112810593586e-08
+    1.807084564390063e-07
+    4.467727419933744e-07
+ 4.92e+10    
+    4.464643841371817e-07
+     1.80725474225714e-07
+    4.372539925025113e-07
+    6.298428814427277e-08
+    1.171431289135409e-07
+     4.37215929008522e-07
+    3.511153571630416e-08
+    6.300673849905522e-08
+    1.807943978494932e-07
+    4.468994234587582e-07
+ 4.93e+10    
+    4.465913605567875e-07
+    1.808113418436336e-07
+    4.373507829714328e-07
+    6.299962197792955e-08
+    1.171980878813594e-07
+     4.37312803433424e-07
+    3.509444419888163e-08
+    6.302222003616097e-08
+    1.808803927638626e-07
+    4.470263038889959e-07
+ 4.94e+10    
+    4.467185363096733e-07
+    1.808972622712752e-07
+    4.374476935687085e-07
+    6.301482643704893e-08
+    1.172530356573643e-07
+    4.374097979939307e-07
+    3.507717893342415e-08
+    6.303757257967578e-08
+    1.809664408952322e-07
+    4.471533832681922e-07
+ 4.95e+10    
+    4.468459113803448e-07
+    1.809832352206964e-07
+    4.375447242639203e-07
+    6.302990138592929e-08
+    1.173079721986025e-07
+    4.375069126577026e-07
+    3.505974010026857e-08
+    6.305279599326494e-08
+    1.810525419559971e-07
+    4.472806615799827e-07
+ 4.96e+10    
+    4.469734857528519e-07
+    1.810692604032416e-07
+    4.376418750268143e-07
+    6.304484669014064e-08
+    1.173628974631386e-07
+    4.376041473925634e-07
+    3.504212788181119e-08
+    6.306789014186037e-08
+    1.811386956578388e-07
+    4.474081388075435e-07
+ 4.97e+10    
+    4.471012594107929e-07
+    1.811553375295501e-07
+    4.377391458273057e-07
+    6.305966221654853e-08
+    1.174178114100582e-07
+    4.377015021665106e-07
+    3.502434246253897e-08
+    6.308285489168475e-08
+     1.81224901711734e-07
+    4.475358149335984e-07
+ 4.98e+10    
+    4.472292323373276e-07
+    1.812414663095654e-07
+    4.378365366354835e-07
+    6.307434783333811e-08
+     1.17472713999473e-07
+     4.37798976947718e-07
+    3.500638402906063e-08
+    6.309769011027523e-08
+    1.813111598279632e-07
+    4.476636899404291e-07
+ 4.99e+10    
+    4.473574045151822e-07
+    1.813276464525432e-07
+    4.379340474216136e-07
+    6.308890341003766e-08
+    1.175276051925236e-07
+    4.378965717045393e-07
+    3.498825277013735e-08
+    6.311239566650715e-08
+    1.813974697161195e-07
+    4.477917638098821e-07
+ 5e+10       
+    4.474857759266584e-07
+    1.814138776670604e-07
+    4.380316781561442e-07
+    6.310332881754226e-08
+    1.175824849513841e-07
+    4.379942864055146e-07
+    3.496994887671342e-08
+    6.312697143061748e-08
+    1.814838310851171e-07
+    4.479200365233771e-07
+ 5.01e+10    
+     4.47614346553642e-07
+     1.81500159661023e-07
+    4.381294288097091e-07
+    6.311762392813693e-08
+    1.176373532392651e-07
+    4.380921210193717e-07
+    3.495147254194655e-08
+     6.31414172742279e-08
+    1.815702436431992e-07
+    4.480485080619174e-07
+ 5.02e+10    
+    4.477431163776115e-07
+    1.815864921416756e-07
+    4.382272993531327e-07
+    6.313178861551997e-08
+    1.176922100204184e-07
+    4.381900755150331e-07
+     3.49328239612381e-08
+    6.315573307036817e-08
+    1.816567070979475e-07
+    4.481771784060948e-07
+ 5.03e+10    
+    4.478720853796439e-07
+    1.816728748156081e-07
+    4.383252897574335e-07
+    6.314582275482583e-08
+      1.1774705526014e-07
+    4.382881498616192e-07
+    3.491400333226282e-08
+    6.316991869349881e-08
+    1.817432211562892e-07
+    4.483060475360998e-07
+ 5.04e+10    
+    4.480012535404239e-07
+    1.817593073887643e-07
+    4.384233999938273e-07
+    6.315972622264772e-08
+    1.178018889247735e-07
+    4.383863440284518e-07
+    3.489501085499862e-08
+    6.318397401953381e-08
+    1.818297855245057e-07
+    4.484351154317294e-07
+ 5.05e+10    
+     4.48130620840253e-07
+    1.818457895664513e-07
+    4.385216300337325e-07
+    6.317349889706049e-08
+    1.178567109817144e-07
+    4.384846579850588e-07
+    3.487584673175606e-08
+    6.319789892586325e-08
+     1.81916399908241e-07
+    4.485643820723938e-07
+ 5.06e+10    
+    4.482601872590556e-07
+    1.819323210533457e-07
+     4.38619979848774e-07
+    6.318714065764275e-08
+    1.179115213994132e-07
+    4.385830917011786e-07
+    3.485651116720739e-08
+     6.32116932913755e-08
+    1.820030640125089e-07
+    4.486938474371261e-07
+ 5.07e+10    
+    4.483899527763849e-07
+    1.820189015535021e-07
+    4.387184494107871e-07
+    6.320065138549915e-08
+    1.179663201473791e-07
+     4.38681645146764e-07
+     3.48370043684155e-08
+    6.322535699647937e-08
+    1.820897775417015e-07
+    4.488235115045883e-07
+ 5.08e+10    
+    4.485199173714345e-07
+     1.82105530770361e-07
+    4.388170386918193e-07
+    6.321403096328233e-08
+    1.180211071961829e-07
+    4.387803182919859e-07
+    3.481732654486274e-08
+    6.323888992312611e-08
+    1.821765401995968e-07
+    4.489533742530804e-07
+ 5.09e+10    
+     4.48650081023043e-07
+    1.821922084067567e-07
+    4.389157476641368e-07
+    6.322727927521486e-08
+     1.18075882517461e-07
+    4.388791111072361e-07
+    3.479747790847918e-08
+    6.325229195483101e-08
+    1.822633516893661e-07
+    4.490834356605456e-07
+ 5.1e+10     
+    4.487804437097021e-07
+    1.822789341649244e-07
+    4.390145763002274e-07
+     6.32403962071106e-08
+    1.181306460839185e-07
+    4.389780235631345e-07
+    3.477745867367087e-08
+    6.326556297669513e-08
+    1.823502117135822e-07
+    4.492136957045819e-07
+ 5.11e+10    
+    4.489110054095642e-07
+    1.823657077465079e-07
+    4.391135245728032e-07
+    6.325338164639634e-08
+    1.181853978693326e-07
+     4.39077055630529e-07
+    3.475726905734765e-08
+    6.327870287542635e-08
+    1.824371199742263e-07
+    4.493441543624441e-07
+ 5.12e+10    
+    4.490417661004502e-07
+    1.824525288525675e-07
+    4.392125924548057e-07
+    6.326623548213286e-08
+    1.182401378485554e-07
+    4.391762072805017e-07
+    3.473690927895097e-08
+    6.329171153936087e-08
+    1.825240761726956e-07
+    4.494748116110562e-07
+ 5.13e+10    
+    4.491727257598529e-07
+    1.825393971835866e-07
+     4.39311779919409e-07
+    6.327895760503595e-08
+    1.182948659975178e-07
+    4.392754784843719e-07
+    3.471637956048101e-08
+    6.330458885848394e-08
+    1.826110800098113e-07
+    4.496056674270164e-07
+ 5.14e+10    
+      4.4930388436495e-07
+    1.826263124394791e-07
+    4.394110869400217e-07
+    6.329154790749724e-08
+    1.183495822932319e-07
+    4.393748692137002e-07
+    3.469568012652384e-08
+    6.331733472445049e-08
+    1.826981311858246e-07
+    4.497367217866021e-07
+ 5.15e+10    
+     4.49435241892608e-07
+    1.827132743195975e-07
+    4.395105134902941e-07
+     6.33040062836049e-08
+    1.184042867137948e-07
+    4.394743794402915e-07
+    3.467481120427838e-08
+      6.3329949030606e-08
+    1.827852294004252e-07
+    4.498679746657821e-07
+ 5.16e+10    
+    4.495667983193859e-07
+    1.828002825227384e-07
+    4.396100595441172e-07
+    6.331633262916381e-08
+    1.184589792383911e-07
+    4.395740091361998e-07
+    3.465377302358266e-08
+    6.334243167200652e-08
+    1.828723743527472e-07
+    4.499994260402186e-07
+ 5.17e+10    
+    4.496985536215495e-07
+    1.828873367471508e-07
+    4.397097250756304e-07
+    6.332852684171588e-08
+    1.185136598472961e-07
+    4.396737582737283e-07
+    3.463256581694024e-08
+    6.335478254543913e-08
+     1.82959565741377e-07
+    4.501310758852774e-07
+ 5.18e+10    
+    4.498305077750703e-07
+    1.829744366905426e-07
+     4.39809510059222e-07
+    6.334058882056019e-08
+    1.185683285218791e-07
+    4.397736268254385e-07
+    3.461118981954603e-08
+    6.336700154944156e-08
+    1.830468032643598e-07
+     4.50262924176033e-07
+ 5.19e+10    
+    4.499626607556386e-07
+    1.830615820500874e-07
+    4.399094144695338e-07
+    6.335251846677254e-08
+    1.186229852446058e-07
+    4.398736147641494e-07
+    3.458964526931202e-08
+    6.337908858432207e-08
+    1.831340866192063e-07
+    4.503949708872763e-07
+ 5.2e+10     
+    4.500950125386655e-07
+    1.831487725224311e-07
+     4.40009438281464e-07
+     6.33643156832251e-08
+    1.186776299990414e-07
+    4.399737220629416e-07
+    3.456793240689251e-08
+    6.339104355217892e-08
+    1.832214155028999e-07
+    4.505272159935197e-07
+ 5.21e+10    
+    4.502275630992912e-07
+    1.832360078036989e-07
+    4.401095814701708e-07
+    6.337598037460588e-08
+    1.187322627698534e-07
+    4.400739486951622e-07
+    3.454605147570929e-08
+    6.340286635691993e-08
+    1.833087896119029e-07
+    4.506596594690068e-07
+ 5.22e+10    
+    4.503603124123927e-07
+    1.833232875895016e-07
+    4.402098440110755e-07
+    6.338751244743784e-08
+    1.187868835428146e-07
+     4.40174294634427e-07
+    3.452400272197621e-08
+    6.341455690428117e-08
+    1.833962086421636e-07
+    4.507923012877153e-07
+ 5.23e+10    
+    4.504932604525886e-07
+    1.834106115749425e-07
+    4.403102258798659e-07
+    6.339891181009778e-08
+    1.188414923048055e-07
+    4.402747598546234e-07
+    3.450178639472373e-08
+     6.34261151018462e-08
+    1.834836722891221e-07
+    4.509251414233658e-07
+ 5.24e+10    
+    4.506264071942438e-07
+    1.834979794546233e-07
+    4.404107270524992e-07
+    6.341017837283507e-08
+    1.188960890438172e-07
+    4.403753443299145e-07
+     3.44794027458229e-08
+    6.343754085906457e-08
+    1.835711802477172e-07
+    4.510581798494275e-07
+ 5.25e+10    
+    4.507597526114803e-07
+    1.835853909226508e-07
+    4.405113475052049e-07
+    6.342131204779045e-08
+    1.189506737489539e-07
+     4.40476048034742e-07
+    3.445685203000926e-08
+    6.344883408727045e-08
+     1.83658732212393e-07
+    4.511914165391251e-07
+ 5.26e+10    
+    4.508932966781787e-07
+    1.836728456726431e-07
+    4.406120872144888e-07
+    6.343231274901402e-08
+    1.190052464104357e-07
+    4.405768709438297e-07
+    3.443413450490623e-08
+    6.345999469970078e-08
+    1.837463278771043e-07
+    4.513248514654432e-07
+ 5.27e+10    
+    4.510270393679868e-07
+     1.83760343397736e-07
+    4.407129461571349e-07
+    6.344318039248354e-08
+    1.190598070196013e-07
+    4.406778130321859e-07
+    3.441125043104825e-08
+    6.347102261151342e-08
+    1.838339669353237e-07
+    4.514584846011345e-07
+ 5.28e+10    
+    4.511609806543252e-07
+    1.838478837905886e-07
+    4.408139243102087e-07
+    6.345391489612219e-08
+    1.191143555689097e-07
+    4.407788742751068e-07
+    3.438820007190361e-08
+    6.348191773980489e-08
+    1.839216490800473e-07
+    4.515923159187248e-07
+ 5.29e+10    
+    4.512951205103927e-07
+    1.839354665433898e-07
+    4.409150216510615e-07
+     6.34645161798165e-08
+     1.19168892051944e-07
+    4.408800546481794e-07
+    3.436498369389688e-08
+    6.349268000362812e-08
+    1.840093740038004e-07
+    4.517263453905192e-07
+ 5.3e+10     
+     4.51429458909173e-07
+    1.840230913478641e-07
+    4.410162381573324e-07
+    6.347498416543353e-08
+    1.192234164634126e-07
+    4.409813541272857e-07
+    3.434160156643111e-08
+    6.350330932400976e-08
+     1.84097141398644e-07
+    4.518605729886074e-07
+ 5.31e+10    
+     4.51563995823438e-07
+    1.841107578952772e-07
+    4.411175738069484e-07
+    6.348531877683829e-08
+    1.192779287991523e-07
+    4.410827726886028e-07
+    3.431805396190958e-08
+    6.351380562396754e-08
+    1.841849509561805e-07
+    4.519949986848713e-07
+ 5.32e+10    
+    4.516987312257584e-07
+     1.84198465876443e-07
+    4.412190285781337e-07
+    6.349551993991084e-08
+    1.193324290561307e-07
+    4.411843103086099e-07
+    3.429434115575728e-08
+     6.35241688285271e-08
+    1.842728023675597e-07
+    4.521296224509889e-07
+ 5.33e+10    
+    4.518336650885038e-07
+    1.842862149817274e-07
+    4.413206024494059e-07
+    6.350558758256285e-08
+    1.193869172324476e-07
+    4.412859669640869e-07
+    3.427046342644195e-08
+    6.353439886473877e-08
+    1.843606953234836e-07
+     4.52264444258441e-07
+ 5.34e+10    
+    4.519687973838515e-07
+    1.843740049010554e-07
+    4.414222953995823e-07
+    6.351552163475448e-08
+    1.194413933273386e-07
+    4.413877426321204e-07
+    3.424642105549496e-08
+    6.354449566169428e-08
+    1.844486295142134e-07
+    4.523994640785157e-07
+ 5.35e+10    
+    4.521041280837918e-07
+    1.844618353239165e-07
+    4.415241074077828e-07
+    6.352532202851064e-08
+    1.194958573411764e-07
+    4.414896372901049e-07
+    3.422221432753157e-08
+     6.35544591505429e-08
+     1.84536604629574e-07
+    4.525346818823152e-07
+ 5.36e+10    
+    4.522396571601321e-07
+    1.845497059393697e-07
+    4.416260384534308e-07
+    6.353498869793706e-08
+    1.195503092754732e-07
+    4.415916509157455e-07
+    3.419784353027112e-08
+    6.356428926450772e-08
+    1.846246203589602e-07
+    4.526700976407615e-07
+ 5.37e+10    
+    4.523753845845034e-07
+    1.846376164360494e-07
+    4.417280885162569e-07
+    6.354452157923651e-08
+    1.196047491328829e-07
+    4.416937834870623e-07
+    3.417330895455659e-08
+    6.357398593890144e-08
+    1.847126763913416e-07
+    4.528057113245995e-07
+ 5.38e+10    
+    4.525113103283652e-07
+    1.847255665021708e-07
+    4.418302575763017e-07
+    6.355392061072418e-08
+    1.196591769172033e-07
+    4.417960349823904e-07
+    3.414861089437403e-08
+    6.358354911114208e-08
+    1.848007724152684e-07
+    4.529415229044058e-07
+ 5.39e+10    
+    4.526474343630099e-07
+    1.848135558255345e-07
+    4.419325456139179e-07
+    6.356318573284349e-08
+    1.197135926333777e-07
+    4.418984053803856e-07
+    3.412374964687142e-08
+    6.359297872076848e-08
+    1.848889081188762e-07
+    4.530775323505903e-07
+ 5.4e+10     
+    4.527837566595693e-07
+    1.849015840935327e-07
+    4.420349526097732e-07
+    6.357231688818112e-08
+    1.197679962874977e-07
+    4.420008946600236e-07
+     3.40987255123774e-08
+    6.360227470945553e-08
+     1.84977083189892e-07
+    4.532137396334047e-07
+ 5.41e+10    
+    4.529202771890194e-07
+    1.849896509931538e-07
+    4.421374785448522e-07
+    6.358131402148227e-08
+    1.198223878868043e-07
+    4.421035028006052e-07
+    3.407353879441929e-08
+    6.361143702102907e-08
+    1.850652973156379e-07
+    4.533501447229441e-07
+ 5.42e+10    
+    4.530569959221839e-07
+    1.850777562109875e-07
+    4.422401234004603e-07
+    6.359017707966534e-08
+    1.198767674396905e-07
+    4.422062297817576e-07
+    3.404818979974112e-08
+    6.362046560148084e-08
+    1.851535501830383e-07
+    4.534867475891556e-07
+ 5.43e+10    
+    4.531939128297412e-07
+    1.851658994332299e-07
+    4.423428871582238e-07
+    6.359890601183661e-08
+    1.199311349557028e-07
+    4.423090755834383e-07
+    3.402267883832099e-08
+    6.362936039898295e-08
+    1.852418414786228e-07
+    4.536235482018408e-07
+ 5.44e+10    
+     4.53331027882228e-07
+    1.852540803456886e-07
+    4.424457698000949e-07
+    6.360750076930471e-08
+    1.199854904455432e-07
+    4.424120401859349e-07
+    3.399700622338822e-08
+     6.36381213639023e-08
+    1.853301708885323e-07
+    4.537605465306621e-07
+ 5.45e+10    
+     4.53468341050044e-07
+    1.853422986337875e-07
+    4.425487713083524e-07
+    6.361596130559462e-08
+    1.200398339210711e-07
+    4.425151235698705e-07
+    3.397117227143997e-08
+    6.364674844881466e-08
+     1.85418538098524e-07
+    4.538977425451468e-07
+ 5.46e+10    
+    4.536058523034569e-07
+    1.854305539825711e-07
+    4.426518916656041e-07
+     6.36242875764616e-08
+    1.200941653953048e-07
+    4.426183257162027e-07
+     3.39451773022576e-08
+    6.365524160851851e-08
+    1.855069427939752e-07
+    4.540351362146917e-07
+ 5.47e+10    
+     4.53743561612608e-07
+    1.855188460767102e-07
+    4.427551308547904e-07
+    6.363247953990513e-08
+    1.201484848824235e-07
+    4.427216466062293e-07
+    3.391902163892263e-08
+    6.366360080004881e-08
+    1.855953846598886e-07
+    4.541727275085679e-07
+ 5.48e+10    
+    4.538814689475148e-07
+    1.856071746005059e-07
+    4.428584888591847e-07
+    6.364053715618219e-08
+    1.202027923977687e-07
+    4.428250862215894e-07
+    3.389270560783219e-08
+    6.367182598269039e-08
+    1.856838633808978e-07
+    4.543105163959256e-07
+ 5.49e+10    
+    4.540195742780773e-07
+    1.856955392378942e-07
+    4.429619656623972e-07
+    6.364846038782048e-08
+    1.202570879578461e-07
+    4.429286445442641e-07
+    3.386622953871426e-08
+    6.367991711799125e-08
+    1.857723786412704e-07
+    4.544485028457993e-07
+ 5.5e+10     
+     4.54157877574081e-07
+    1.857839396724512e-07
+    4.430655612483761e-07
+     6.36562491996317e-08
+    1.203113715803272e-07
+    4.430323215565811e-07
+    3.383959376464229e-08
+    6.368787416977542e-08
+    1.858609301249131e-07
+    4.545866868271114e-07
+ 5.51e+10    
+    4.542963788052029e-07
+    1.858723755873966e-07
+    4.431692756014102e-07
+    6.366390355872405e-08
+    1.203656432840507e-07
+    4.431361172412145e-07
+    3.381279862204964e-08
+    6.369569710415582e-08
+    1.859495175153768e-07
+    4.547250683086766e-07
+ 5.52e+10    
+    4.544350779410158e-07
+    1.859608466655991e-07
+    4.432731087061317e-07
+    6.367142343451503e-08
+     1.20419903089024e-07
+    4.432400315811894e-07
+    3.378584445074351e-08
+    6.370338588954685e-08
+    1.860381404958603e-07
+    4.548636472592066e-07
+ 5.53e+10    
+    4.545739749509889e-07
+    1.860493525895802e-07
+    4.433770605475161e-07
+    6.367880879874367e-08
+     1.20474151016425e-07
+    4.433440645598834e-07
+    3.375873159391837e-08
+    6.371094049667647e-08
+    1.861267987492146e-07
+    4.550024236473137e-07
+ 5.54e+10    
+    4.547130698044972e-07
+    1.861378930415183e-07
+     4.43481131110887e-07
+    6.368605962548262e-08
+    1.205283870886029e-07
+    4.434482161610257e-07
+    3.373146039816926e-08
+    6.371836089859862e-08
+    1.862154919579478e-07
+    4.551413974415172e-07
+ 5.55e+10    
+    4.548523624708225e-07
+    1.862264677032536e-07
+    4.435853203819163e-07
+    6.369317589115018e-08
+    1.205826113290807e-07
+    4.435524863687038e-07
+    3.370403121350434e-08
+    6.372564707070487e-08
+    1.863042198042286e-07
+    4.552805686102442e-07
+ 5.56e+10    
+    4.549918529191579e-07
+    1.863150762562918e-07
+    4.436896283466268e-07
+    6.370015757452184e-08
+    1.206368237625551e-07
+    4.436568751673627e-07
+    3.367644439335727e-08
+    6.373279899073597e-08
+    1.863929819698906e-07
+    4.554199371218361e-07
+ 5.57e+10    
+    4.551315411186126e-07
+    1.864037183818082e-07
+    4.437940549913946e-07
+    6.370700465674171e-08
+    1.206910244148992e-07
+    4.437613825418062e-07
+    3.364870029459913e-08
+    6.373981663879347e-08
+    1.864817781364373e-07
+    4.555595029445527e-07
+ 5.58e+10    
+    4.552714270382151e-07
+    1.864923937606518e-07
+    4.438986003029491e-07
+    6.371371712133373e-08
+     1.20745213313163e-07
+    4.438660084772021e-07
+    3.362079927754983e-08
+    6.374669999735067e-08
+    1.865706079850445e-07
+     4.55699266046574e-07
+ 5.59e+10    
+    4.554115106469171e-07
+    1.865811020733497e-07
+    4.440032642683781e-07
+    6.372029495421267e-08
+    1.207993904855747e-07
+    4.439707529590802e-07
+    3.359274170598921e-08
+    6.375344905126381e-08
+    1.866594711965655e-07
+    4.558392263960069e-07
+ 5.6e+10     
+    4.555517919135984e-07
+    1.866698430001104e-07
+    4.441080468751266e-07
+    6.372673814369483e-08
+    1.208535559615421e-07
+    4.440756159733374e-07
+    3.356452794716763e-08
+    6.376006378778241e-08
+    1.867483674515347e-07
+    4.559793839608862e-07
+ 5.61e+10    
+    4.556922708070686e-07
+     1.86758616220828e-07
+    4.442129481110013e-07
+     6.37330466805086e-08
+    1.209077097716538e-07
+    4.441805975062377e-07
+    3.353615837181628e-08
+    6.376654419656026e-08
+    1.868372964301716e-07
+    4.561197387091821e-07
+ 5.62e+10    
+    4.558329472960722e-07
+    1.868474214150858e-07
+    4.443179679641687e-07
+    6.373922055780462e-08
+    1.209618519476804e-07
+    4.442856975444147e-07
+     3.35076333541568e-08
+    6.377289026966507e-08
+    1.869262578123839e-07
+    4.562602906087987e-07
+ 5.63e+10    
+    4.559738213492935e-07
+    1.869362582621605e-07
+    4.444231064231616e-07
+    6.374525977116587e-08
+    1.210159825225747e-07
+     4.44390916074872e-07
+    3.347895327191083e-08
+    6.377910200158889e-08
+    1.870152512777717e-07
+    4.564010396275821e-07
+ 5.64e+10    
+    4.561148929353569e-07
+    1.870251264410253e-07
+    4.445283634768771e-07
+    6.375116431861749e-08
+    1.210701015304742e-07
+    4.444962530849874e-07
+    3.345011850630882e-08
+    6.378517938925796e-08
+    1.871042765056317e-07
+    4.565419857333241e-07
+ 5.65e+10    
+    4.562561620228329e-07
+    1.871140256303542e-07
+    4.446337391145804e-07
+    6.375693420063647e-08
+    1.211242090067011e-07
+    4.446017085625135e-07
+     3.34211294420985e-08
+    6.379112243204179e-08
+    1.871933331749598e-07
+    4.566831288937605e-07
+ 5.66e+10    
+    4.563976285802407e-07
+    1.872029555085248e-07
+    4.447392333259051e-07
+    6.376256942016075e-08
+    1.211783049877635e-07
+    4.447072824955782e-07
+    3.339198646755316e-08
+    6.379693113176312e-08
+    1.872824209644555e-07
+    4.568244690765817e-07
+ 5.67e+10    
+    4.565392925760522e-07
+    1.872919157536223e-07
+    4.448448461008555e-07
+    6.376806998259852e-08
+    1.212323895113564e-07
+    4.448129748726882e-07
+      3.3362689974479e-08
+    6.380260549270638e-08
+    1.873715395525248e-07
+    4.569660062494301e-07
+ 5.68e+10    
+    4.566811539786949e-07
+    1.873809060434431e-07
+    4.449505774298086e-07
+    6.377343589583695e-08
+    1.212864626163623e-07
+    4.449187856827285e-07
+    3.333324035822253e-08
+    6.380814552162697e-08
+    1.874606886172839e-07
+    4.571077403799073e-07
+ 5.69e+10    
+    4.568232127565544e-07
+    1.874699260554982e-07
+    4.450564273035154e-07
+     6.37786671702511e-08
+    1.213405243428528e-07
+     4.45024714914967e-07
+    3.330363801767733e-08
+    6.381355122775984e-08
+    1.875498678365629e-07
+    4.572496714355755e-07
+ 5.7e+10     
+    4.569654688779797e-07
+    1.875589754670158e-07
+    4.451623957131016e-07
+    6.378376381871194e-08
+    1.213945747320884e-07
+    4.451307625590523e-07
+     3.32738833552902e-08
+    6.381882262282765e-08
+    1.876390768879082e-07
+    4.573917993839609e-07
+ 5.71e+10    
+    4.571079223112838e-07
+    1.876480539549458e-07
+    4.452684826500709e-07
+    6.378872585659494e-08
+    1.214486138265203e-07
+    4.452369286050192e-07
+    3.324397677706728e-08
+    6.382395972104924e-08
+    1.877283154485872e-07
+    4.575341241925587e-07
+ 5.72e+10    
+    4.572505730247493e-07
+    1.877371611959618e-07
+    4.453746881063037e-07
+    6.379355330178769e-08
+    1.215026416697899e-07
+    4.453432130432872e-07
+    3.321391869257934e-08
+    6.382896253914717e-08
+      1.8781758319559e-07
+    4.576766458288322e-07
+ 5.73e+10    
+    4.573934209866295e-07
+    1.878262968664655e-07
+    4.454810120740623e-07
+    6.379824617469778e-08
+     1.21556658306731e-07
+    4.454496158646625e-07
+    3.318370951496681e-08
+    6.383383109635594e-08
+    1.879068798056336e-07
+    4.578193642602213e-07
+ 5.74e+10    
+    4.575364661651528e-07
+    1.879154606425892e-07
+    4.455874545459896e-07
+    6.380280449826031e-08
+    1.216106637833691e-07
+    4.455561370603413e-07
+    3.315334966094444e-08
+    6.383856541442907e-08
+    1.879962049551652e-07
+    4.579622794541409e-07
+ 5.75e+10    
+    4.576797085285241e-07
+    1.880046522001985e-07
+     4.45694015515111e-07
+    6.380722829794497e-08
+     1.21664658146923e-07
+    4.456627766219084e-07
+    3.312283955080523e-08
+    6.384316551764636e-08
+    1.880855583203638e-07
+    4.581053913779859e-07
+ 5.76e+10    
+    4.578231480449304e-07
+    1.880938712148965e-07
+    4.458006949748366e-07
+    6.381151760176324e-08
+    1.217186414458045e-07
+    4.457695345413401e-07
+    3.309217960842427e-08
+    6.384763143282107e-08
+    1.881749395771452e-07
+    4.582486999991338e-07
+ 5.77e+10    
+      4.5796678468254e-07
+     1.88183117362026e-07
+     4.45907492918962e-07
+    6.381567244027502e-08
+      1.2177261372962e-07
+    4.458764108110069e-07
+    3.306137026126184e-08
+    6.385196318930652e-08
+    1.882643484011634e-07
+    4.583922052849475e-07
+ 5.78e+10    
+    4.581106184095083e-07
+    1.882723903166719e-07
+    4.460144093416684e-07
+    6.381969284659532e-08
+    1.218265750491699e-07
+    4.459834054236716e-07
+    3.303041194036625e-08
+    6.385616081900273e-08
+    1.883537844678144e-07
+    4.585359072027779e-07
+ 5.79e+10    
+    4.582546491939798e-07
+    1.883616897536659e-07
+    4.461214442375274e-07
+    6.382357885640053e-08
+      1.2188052545645e-07
+    4.460905183724935e-07
+    3.299930508037624e-08
+    6.386022435636273e-08
+    1.884432474522388e-07
+    4.586798057199676e-07
+ 5.8e+10     
+    4.583988770040892e-07
+    1.884510153475872e-07
+    4.462285976014989e-07
+    6.382733050793434e-08
+    1.219344650046512e-07
+    4.461977496510279e-07
+    3.296805011952259e-08
+    6.386415383839853e-08
+    1.885327370293241e-07
+    4.588239008038518e-07
+ 5.81e+10    
+     4.58543301807966e-07
+    1.885403667727671e-07
+    4.463358694289328e-07
+    6.383094784201386e-08
+    1.219883937481602e-07
+    4.463050992532276e-07
+    3.293664749962987e-08
+    6.386794930468711e-08
+     1.88622252873709e-07
+    4.589681924217627e-07
+ 5.82e+10    
+    4.586879235737375e-07
+    1.886297437032906e-07
+    4.464432597155724e-07
+    6.383443090203514e-08
+    1.220423117425602e-07
+    4.464125671734453e-07
+     3.29050976661172e-08
+    6.387161079737594e-08
+    1.887117946597842e-07
+    4.591126805410313e-07
+ 5.83e+10    
+    4.588327422695279e-07
+    1.887191458129993e-07
+    4.465507684575524e-07
+    6.383777973397839e-08
+    1.220962190446307e-07
+    4.465201534064339e-07
+    3.287340106799884e-08
+     6.38751383611883e-08
+    1.888013620616965e-07
+    4.592573651289895e-07
+ 5.84e+10    
+    4.589777578634655e-07
+    1.888085727754949e-07
+     4.46658395651404e-07
+    6.384099438641337e-08
+    1.221501157123478e-07
+    4.466278579473467e-07
+    3.284155815788423e-08
+    6.387853204342862e-08
+    1.888909547533506e-07
+    4.594022461529732e-07
+ 5.85e+10    
+    4.591229703236807e-07
+    1.888980242641404e-07
+    4.467661412940515e-07
+    6.384407491050421e-08
+    1.222040018048848e-07
+    4.467356807917402e-07
+    3.280956939197767e-08
+    6.388179189398726e-08
+    1.889805724084124e-07
+    4.595473235803247e-07
+ 5.86e+10    
+    4.592683796183121e-07
+    1.889874999520641e-07
+    4.468740053828175e-07
+    6.384702136001411e-08
+     1.22257877382612e-07
+    4.468436219355747e-07
+     3.27774352300774e-08
+     6.38849179653452e-08
+    1.890702147003111e-07
+     4.59692597378395e-07
+ 5.87e+10    
+    4.594139857155071e-07
+    1.890769995121612e-07
+    4.469819879154212e-07
+    6.384983379130976e-08
+    1.223117425070974e-07
+    4.469516813752141e-07
+    3.274515613557434e-08
+    6.388791031257846e-08
+    1.891598813022412e-07
+    4.598380675145461e-07
+ 5.88e+10    
+    4.595597885834228e-07
+    1.891665226170965e-07
+    4.470900888899819e-07
+    6.385251226336561e-08
+    1.223655972411061e-07
+    4.470598591074298e-07
+    3.271273257545037e-08
+    6.389076899336253e-08
+    1.892495718871662e-07
+    4.599837339561522e-07
+ 5.89e+10    
+    4.597057881902317e-07
+    1.892560689393071e-07
+    4.471983083050172e-07
+    6.385505683776798e-08
+    1.224194416486012e-07
+    4.471681551293979e-07
+    3.268016502027617e-08
+    6.389349406797624e-08
+    1.893392861278205e-07
+    4.601295966706058e-07
+ 5.9e+10     
+    4.598519845041212e-07
+    1.893456381510043e-07
+    4.473066461594462e-07
+    6.385746757871861e-08
+     1.22473275794743e-07
+    4.472765694387042e-07
+    3.264745394420836e-08
+    6.389608559930536e-08
+    1.894290236967108e-07
+    4.602756556253134e-07
+ 5.91e+10    
+    4.599983774932968e-07
+    1.894352299241765e-07
+    4.474151024525899e-07
+     6.38597445530383e-08
+    1.225270997458899e-07
+    4.473851020333416e-07
+    3.261459982498668e-08
+    6.389854365284644e-08
+    1.895187842661197e-07
+    4.604219107877043e-07
+ 5.92e+10    
+    4.601449671259826e-07
+     1.89524843930591e-07
+     4.47523677184171e-07
+    6.386188783017021e-08
+    1.225809135695975e-07
+    4.474937529117127e-07
+    3.258160314393019e-08
+    6.390086829670988e-08
+    1.896085675081076e-07
+    4.605683621252281e-07
+ 5.93e+10    
+    4.602917533704271e-07
+    1.896144798417968e-07
+    4.476323703543178e-07
+    6.386389748218305e-08
+    1.226347173346193e-07
+    4.476025220726323e-07
+    3.254846438593335e-08
+    6.390305960162321e-08
+    1.896983730945147e-07
+    4.607150096053583e-07
+ 5.94e+10    
+    4.604387361949016e-07
+    1.897041373291266e-07
+    4.477411819635618e-07
+    6.386577358377378e-08
+    1.226885111109063e-07
+     4.47711409515325e-07
+    3.251518403946159e-08
+    6.390511764093379e-08
+    1.897882006969634e-07
+    4.608618531955959e-07
+ 5.95e+10    
+     4.60585915567704e-07
+    1.897938160636985e-07
+    4.478501120128407e-07
+    6.386751621227027e-08
+    1.227422949696066e-07
+    4.478204152394287e-07
+     3.24817625965463e-08
+    6.390704249061155e-08
+    1.898780499868604e-07
+    4.610088928634682e-07
+ 5.96e+10    
+    4.607332914571591e-07
+     1.89883515716419e-07
+    4.479591605034981e-07
+    6.386912544763364e-08
+    1.227960689830657e-07
+    4.479295392449933e-07
+    3.244820055277944e-08
+    6.390883422925128e-08
+    1.899679206353987e-07
+    4.611561285765332e-07
+ 5.97e+10    
+    4.608808638316231e-07
+    1.899732359579849e-07
+     4.48068327437286e-07
+    6.387060137246071e-08
+    1.228498332248261e-07
+    4.480387815324848e-07
+    3.241449840730781e-08
+    6.391049293807486e-08
+    1.900578123135605e-07
+      4.6130356030238e-07
+ 5.98e+10    
+    4.610286326594841e-07
+    1.900629764588847e-07
+    4.481776128163628e-07
+    6.387194407198551e-08
+    1.229035877696269e-07
+    4.481481421027822e-07
+    3.238065666282667e-08
+    6.391201870093329e-08
+    1.901477246921176e-07
+    4.614511880086322e-07
+ 5.99e+10    
+    4.611765979091621e-07
+    1.901527368894015e-07
+    4.482870166432978e-07
+    6.387315363408133e-08
+     1.22957332693404e-07
+     4.48257620957181e-07
+    3.234667582557303e-08
+    6.391341160430826e-08
+    1.902376574416353e-07
+    4.615990116629483e-07
+ 6e+10       
+     4.61324759549114e-07
+    1.902425169196141e-07
+    4.483965389210681e-07
+    6.387423014926197e-08
+    1.230110680732889e-07
+    4.483672180973917e-07
+    3.231255640531838e-08
+    6.391467173731363e-08
+    1.903276102324727e-07
+    4.617470312330227e-07
+ 6.01e+10    
+    4.614731175478342e-07
+    1.903323162194004e-07
+     4.48506179653063e-07
+    6.387517371068327e-08
+    1.230647939876096e-07
+    4.484769335255447e-07
+    3.227829891536125e-08
+    6.391579919169699e-08
+    1.904175827347859e-07
+    4.618952466865907e-07
+ 6.02e+10    
+    4.616216718738547e-07
+    1.904221344584375e-07
+    4.486159388430821e-07
+    6.387598441414379e-08
+    1.231185105158889e-07
+     4.48586767244185e-07
+    3.224390387251886e-08
+    6.391679406184032e-08
+    1.905075746185292e-07
+    4.620436579914267e-07
+ 6.03e+10    
+    4.617704224957486e-07
+    1.905119713062052e-07
+     4.48725816495337e-07
+    6.387666235808601e-08
+    1.231722177388452e-07
+    4.486967192562786e-07
+    3.220937179711875e-08
+    6.391765644476115e-08
+    1.905975855534574e-07
+     4.62192265115348e-07
+ 6.04e+10    
+    4.619193693821324e-07
+    1.906018264319868e-07
+    4.488358126144526e-07
+    6.387720764359667e-08
+    1.232259157383912e-07
+    4.488067895652096e-07
+    3.217470321298971e-08
+    6.391838644011288e-08
+     1.90687615209127e-07
+    4.623410680262145e-07
+ 6.05e+10    
+    4.620685125016642e-07
+    1.906916995048716e-07
+    4.489459272054667e-07
+    6.387762037440709e-08
+    1.232796045976334e-07
+     4.48916978174782e-07
+    3.213989864745236e-08
+    6.391898415018539e-08
+    1.907776632548986e-07
+    4.624900666919323e-07
+ 6.06e+10    
+    4.622178518230494e-07
+     1.90781590193756e-07
+    4.490561602738312e-07
+    6.387790065689358e-08
+    1.233332844008722e-07
+    4.490272850892201e-07
+    3.210495863130922e-08
+    6.391944967990497e-08
+    1.908677293599385e-07
+    4.626392610804532e-07
+ 6.07e+10    
+     4.62367387315039e-07
+     1.90871498167346e-07
+    4.491665118254125e-07
+    6.387804860007706e-08
+     1.23386955233601e-07
+    4.491377103131702e-07
+    3.206988369883448e-08
+    6.391978313683456e-08
+    1.909578131932204e-07
+    4.627886511597793e-07
+ 6.08e+10    
+    4.625171189464332e-07
+    1.909614230941585e-07
+    4.492769818664932e-07
+    6.387806431562298e-08
+    1.234406171825055e-07
+    4.492482538516994e-07
+    3.203467438776304e-08
+    6.391998463117311e-08
+    1.910479144235269e-07
+    4.629382368979598e-07
+ 6.09e+10    
+    4.626670466860811e-07
+     1.91051364642523e-07
+    4.493875704037709e-07
+    6.387794791784063e-08
+     1.23494270335463e-07
+    4.493589157102963e-07
+    3.199933123927947e-08
+     6.39200542757554e-08
+    1.911380327194512e-07
+    4.630880182630969e-07
+ 6.1e+10     
+    4.628171705028841e-07
+    1.911413224805834e-07
+      4.4949827744436e-07
+    6.387769952368254e-08
+    1.235479147815422e-07
+    4.494696958948746e-07
+    3.196385479800616e-08
+    6.391999218605111e-08
+    1.912281677493995e-07
+    4.632379952233441e-07
+ 6.11e+10    
+    4.629674903657958e-07
+    1.912312962762996e-07
+    4.496091029957919e-07
+    6.387731925274352e-08
+    1.236015506110019e-07
+    4.495805944117694e-07
+    3.192824561199143e-08
+    6.391979848016392e-08
+    1.913183191815916e-07
+    4.633881677469096e-07
+ 6.12e+10    
+    4.631180062438228e-07
+    1.913212856974491e-07
+    4.497200470660164e-07
+    6.387680722725928e-08
+    1.236551779152909e-07
+     4.49691611267741e-07
+    3.189250423269673e-08
+    6.391947327883046e-08
+    1.914084866840626e-07
+    4.635385358020559e-07
+ 6.13e+10    
+    4.632687181060292e-07
+    1.914112904116286e-07
+    4.498311096634005e-07
+    6.387616357210531e-08
+    1.237087967870465e-07
+    4.498027464699727e-07
+    3.185663121498384e-08
+    6.391901670541875e-08
+    1.914986699246652e-07
+    4.636890993571018e-07
+ 6.14e+10    
+    4.634196259215327e-07
+    1.915013100862548e-07
+    4.499422907967297e-07
+    6.387538841479491e-08
+    1.237624073200942e-07
+    4.499140000260729e-07
+    3.182062711710131e-08
+    6.391842888592675e-08
+    1.915888685710702e-07
+    4.638398583804246e-07
+ 6.15e+10    
+    4.635707296595119e-07
+    1.915913443885681e-07
+    4.500535904752102e-07
+    6.387448188547796e-08
+     1.23816009609447e-07
+    4.500253719440761e-07
+    3.178449250067079e-08
+    6.391770994898061e-08
+     1.91679082290769e-07
+    4.639908128404598e-07
+ 6.16e+10    
+     4.63722029289203e-07
+    1.916813929856314e-07
+    4.501650087084663e-07
+    6.387344411693815e-08
+    1.238696037513039e-07
+    4.501368622324421e-07
+    3.174822793067246e-08
+    6.391686002583241e-08
+    1.917693107510742e-07
+    4.641419627057019e-07
+ 6.17e+10    
+    4.638735247799012e-07
+     1.91771455544333e-07
+    4.502765455065439e-07
+    6.387227524459123e-08
+    1.239231898430497e-07
+    4.502484709000564e-07
+    3.171183397543055e-08
+    6.391587925035823e-08
+    1.918595536191217e-07
+     4.64293307944709e-07
+ 6.18e+10    
+    4.640252161009655e-07
+     1.91861531731388e-07
+    4.503882008799075e-07
+    6.387097540648236e-08
+    1.239767679832533e-07
+    4.503601979562314e-07
+    3.167531120659803e-08
+    6.391476775905541e-08
+    1.919498105618714e-07
+    4.644448485260987e-07
+ 6.19e+10    
+    4.641771032218161e-07
+    1.919516212133396e-07
+    4.504999748394449e-07
+    6.386954474328348e-08
+    1.240303382716675e-07
+    4.504720434107068e-07
+    3.163866019914112e-08
+    6.391352569104017e-08
+    1.920400812461094e-07
+    4.645965844185537e-07
+ 6.2e+10     
+    4.643291861119373e-07
+    1.920417236565601e-07
+    4.506118673964633e-07
+    6.386798339829039e-08
+    1.240839008092276e-07
+    4.505840072736494e-07
+    3.160188153132324e-08
+    6.391215318804455e-08
+    1.921303653384488e-07
+    4.647485155908205e-07
+ 6.21e+10    
+    4.644814647408775e-07
+    1.921318387272529e-07
+    4.507238785626929e-07
+    6.386629151741952e-08
+    1.241374556980502e-07
+    4.506960895556526e-07
+     3.15649757846885e-08
+    6.391065039441333e-08
+    1.922206625053308e-07
+      4.6490064201171e-07
+ 6.22e+10    
+    4.646339390782523e-07
+    1.922219660914536e-07
+    4.508360083502866e-07
+    6.386446924920493e-08
+    1.241910030414324e-07
+    4.508082902677395e-07
+    3.152794354404502e-08
+    6.390901745710099e-08
+    1.923109724130272e-07
+    4.650529636501011e-07
+ 6.23e+10    
+    4.647866090937427e-07
+    1.923121054150306e-07
+     4.50948256771818e-07
+    6.386251674479443e-08
+    1.242445429438505e-07
+    4.509206094213598e-07
+    3.149078539744749e-08
+    6.390725452566789e-08
+    1.924012947276403e-07
+    4.652054804749392e-07
+ 6.24e+10    
+     4.64939474757098e-07
+    1.924022563636875e-07
+    4.510606238402848e-07
+     6.38604341579461e-08
+    1.242980755109593e-07
+    4.510330470283935e-07
+    3.145350193617957e-08
+    6.390536175227682e-08
+    1.924916291151047e-07
+    4.653581924552382e-07
+ 6.25e+10    
+    4.650925360381369e-07
+    1.924924186029641e-07
+    4.511731095691089e-07
+    6.385822164502424e-08
+    1.243516008495901e-07
+    4.511456031011482e-07
+    3.141609375473571e-08
+    6.390333929168895e-08
+    1.925819752411886e-07
+     4.65511099560081e-07
+ 6.26e+10    
+    4.652457929067472e-07
+    1.925825917982371e-07
+    4.512857139721343e-07
+    6.385587936499534e-08
+    1.244051190677505e-07
+    4.512582776523615e-07
+    3.137856145080273e-08
+    6.390118730125982e-08
+    1.926723327714952e-07
+    4.656642017586199e-07
+ 6.27e+10    
+    4.653992453328875e-07
+    1.926727756147216e-07
+     4.51398437063629e-07
+     6.38534074794235e-08
+     1.24458630274622e-07
+    4.513710706952001e-07
+    3.134090562524077e-08
+     6.38989059409349e-08
+    1.927627013714639e-07
+      4.6581749902008e-07
+ 6.28e+10    
+    4.655528932865886e-07
+    1.927629697174726e-07
+     4.51511278858286e-07
+    6.385080615246615e-08
+    1.245121345805599e-07
+    4.514839822432602e-07
+    3.130312688206407e-08
+    6.389649537324535e-08
+    1.928530807063705e-07
+    4.659709913137569e-07
+ 6.29e+10    
+    4.657067367379536e-07
+     1.92853173771386e-07
+    4.516242393712222e-07
+    6.384807555086911e-08
+    1.245656320970911e-07
+    4.515970123105676e-07
+    3.126522582842115e-08
+    6.389395576330289e-08
+    1.929434704413298e-07
+    4.661246786090188e-07
+ 6.3e+10     
+    4.658607756571581e-07
+    1.929433874411995e-07
+    4.517373186179786e-07
+    6.384521584396184e-08
+    1.246191229369134e-07
+    4.517101609115798e-07
+    3.122720307457462e-08
+    6.389128727879524e-08
+    1.930338702412957e-07
+    4.662785608753075e-07
+ 6.31e+10    
+     4.66015010014453e-07
+    1.930336103914943e-07
+    4.518505166145228e-07
+    6.384222720365199e-08
+    1.246726072138935e-07
+    4.518234280611831e-07
+     3.11890592338808e-08
+    6.388849008998081e-08
+     1.93124279771063e-07
+    4.664326380821386e-07
+ 6.32e+10    
+     4.66169439780164e-07
+    1.931238422866958e-07
+    4.519638333772465e-07
+    6.383910980442038e-08
+    1.247260850430662e-07
+    4.519368137746951e-07
+    3.115079492276866e-08
+     6.38855643696836e-08
+     1.93214698695268e-07
+    4.665869101991042e-07
+ 6.33e+10    
+    4.663240649246922e-07
+    1.932140827910746e-07
+    4.520772689229664e-07
+    6.383586382331505e-08
+    1.247795565406325e-07
+    4.520503180678627e-07
+    3.111241076071844e-08
+    6.388251029328734e-08
+    1.933051266783895e-07
+    4.667413771958702e-07
+ 6.34e+10    
+    4.664788854185168e-07
+    1.933043315687484e-07
+    4.521908232689267e-07
+    6.383248943994611e-08
+    1.248330218239585e-07
+    4.521639409568659e-07
+    3.107390737024008e-08
+    6.387932803873025e-08
+    1.933955633847509e-07
+    4.668960390421804e-07
+ 6.35e+10    
+    4.666339012321919e-07
+    1.933945882836818e-07
+    4.523044964327947e-07
+    6.382898683647914e-08
+    1.248864810115737e-07
+    4.522776824583154e-07
+    3.103528537685097e-08
+    6.387601778649858e-08
+    1.934860084785199e-07
+     4.67050895707854e-07
+ 6.36e+10    
+    4.667891123363519e-07
+    1.934848525996889e-07
+    4.524182884326661e-07
+    6.382535619762946e-08
+    1.249399342231692e-07
+    4.523915425892505e-07
+    3.099654540905349e-08
+    6.387257971962107e-08
+      1.9357646162371e-07
+    4.672059471627898e-07
+ 6.37e+10    
+    4.669445187017088e-07
+    1.935751241804328e-07
+    4.525321992870618e-07
+    6.382159771065573e-08
+    1.249933815795968e-07
+    4.525055213671442e-07
+    3.095768809831218e-08
+    6.386901402366239e-08
+    1.936669224841821e-07
+    4.673611933769639e-07
+ 6.38e+10    
+    4.671001202990557e-07
+     1.93665402689428e-07
+    4.526462290149293e-07
+    6.381771156535344e-08
+    1.250468232028671e-07
+    4.526196188099011e-07
+    3.091871407903047e-08
+    6.386532088671662e-08
+    1.937573907236451e-07
+    4.675166343204316e-07
+ 6.39e+10    
+    4.672559170992643e-07
+    1.937556877900403e-07
+    4.527603776356421e-07
+    6.381369795404811e-08
+    1.251002592161474e-07
+    4.527338349358561e-07
+    3.087962398852696e-08
+    6.386150049940071e-08
+    1.938478660056565e-07
+    4.676722699633284e-07
+ 6.4e+10     
+     4.67411909073288e-07
+    1.938459791454886e-07
+    4.528746451690013e-07
+    6.380955707158849e-08
+    1.251536897437608e-07
+    4.528481697637758e-07
+    3.084041846701152e-08
+    6.385755305484758e-08
+    1.939383479936238e-07
+    4.678281002758697e-07
+ 6.41e+10    
+    4.675680961921622e-07
+    1.939362764188457e-07
+     4.52989031635234e-07
+    6.380528911533934e-08
+    1.252071149111839e-07
+    4.529626233128585e-07
+     3.08010981575609e-08
+    6.385347874869906e-08
+    1.940288363508056e-07
+     4.67984125228351e-07
+ 6.42e+10    
+    4.677244784270041e-07
+    1.940265792730392e-07
+    4.531035370549945e-07
+    6.380089428517445e-08
+    1.252605348450457e-07
+    4.530771956027351e-07
+    3.076166370609393e-08
+    6.384927777909878e-08
+    1.941193307403123e-07
+    4.681403447911511e-07
+ 6.43e+10    
+    4.678810557490148e-07
+    1.941168873708526e-07
+    4.532181614493649e-07
+    6.379637278346889e-08
+    1.253139496731254e-07
+    4.531918866534677e-07
+    3.072211576134655e-08
+    6.384495034668463e-08
+    1.942098308251071e-07
+    4.682967589347295e-07
+ 6.44e+10    
+    4.680378281294762e-07
+    1.942072003749254e-07
+    4.533329048398522e-07
+    6.379172481509144e-08
+    1.253673595243507e-07
+    4.533066964855504e-07
+    3.068245497484619e-08
+    6.384049665458126e-08
+    1.943003362680071e-07
+    4.684533676296282e-07
+ 6.45e+10    
+    4.681947955397583e-07
+    1.942975179477558e-07
+     4.53447767248393e-07
+    6.378695058739692e-08
+    1.254207645287959e-07
+    4.534216251199092e-07
+     3.06426820008861e-08
+    6.383591690839218e-08
+    1.943908467316838e-07
+    4.686101708464733e-07
+ 6.46e+10    
+    4.683519579513134e-07
+    1.943878397517003e-07
+    4.535627486973505e-07
+    6.378205031021801e-08
+    1.254741648176804e-07
+    4.535366725779019e-07
+    3.060279749649917e-08
+    6.383121131619201e-08
+    1.944813618786646e-07
+    4.687671685559739e-07
+ 6.47e+10    
+    4.685093153356795e-07
+     1.94478165448975e-07
+    4.536778492095146e-07
+    6.377702419585714e-08
+    1.255275605233666e-07
+    4.536518388813184e-07
+    3.056280212143133e-08
+    6.382638008851822e-08
+    1.945718813713332e-07
+     4.68924360728923e-07
+ 6.48e+10    
+    4.686668676644804e-07
+    1.945684947016561e-07
+    4.537930688081032e-07
+     6.37718724590781e-08
+    1.255809517793582e-07
+    4.537671240523804e-07
+    3.052269653811479e-08
+    6.382142343836279e-08
+    1.946624048719308e-07
+    4.690817473361982e-07
+ 6.49e+10    
+    4.688246149094271e-07
+    1.946588271716821e-07
+    4.539084075167616e-07
+    6.376659531709764e-08
+    1.256343387202978e-07
+     4.53882528113742e-07
+    3.048248141164087e-08
+    6.381634158116382e-08
+    1.947529320425568e-07
+    4.692393283487627e-07
+ 6.5e+10     
+    4.689825570423173e-07
+    1.947491625208532e-07
+    4.540238653595624e-07
+    6.376119298957662e-08
+    1.256877214819654e-07
+    4.539980510884887e-07
+    3.044215740973242e-08
+    6.381113473479687e-08
+    1.948434625451699e-07
+    4.693971037376652e-07
+ 6.51e+10    
+    4.691406940350365e-07
+    1.948395004108333e-07
+    4.541394423610063e-07
+    6.375566569861106e-08
+    1.257411002012763e-07
+    4.541136930001381e-07
+    3.040172520271602e-08
+    6.380580311956615e-08
+     1.94933996041589e-07
+     4.69555073474041e-07
+ 6.52e+10    
+    4.692990258595581e-07
+    1.949298405031503e-07
+    4.542551385460215e-07
+    6.375001366872335e-08
+    1.257944750162793e-07
+    4.542294538726402e-07
+    3.036118546349369e-08
+     6.38003469581953e-08
+    1.950245321934935e-07
+    4.697132375291101e-07
+ 6.53e+10    
+    4.694575524879443e-07
+     1.95020182459197e-07
+    4.543709539399631e-07
+    6.374423712685281e-08
+    1.258478460661542e-07
+     4.54345333730377e-07
+     3.03205388675146e-08
+    6.379476647581857e-08
+    1.951150706624252e-07
+    4.698715958741817e-07
+ 6.54e+10    
+    4.696162738923464e-07
+    1.951105259402325e-07
+    4.544868885686146e-07
+    6.373833630234633e-08
+      1.2590121349121e-07
+    4.544613325981616e-07
+    3.027978609274601e-08
+    6.378906189997124e-08
+    1.952056111097879e-07
+    4.700301484806506e-07
+ 6.55e+10    
+    4.697751900450054e-07
+    1.952008706073827e-07
+    4.546029424581869e-07
+    6.373231142694883e-08
+    1.259545774328828e-07
+    4.545774505012386e-07
+    3.023892781964436e-08
+    6.378323346058018e-08
+    1.952961531968494e-07
+    4.701888953200003e-07
+ 6.56e+10    
+     4.69934300918253e-07
+     1.95291216121641e-07
+    4.547191156353187e-07
+    6.372616273479359e-08
+    1.260079380337338e-07
+    4.546936874652866e-07
+    3.019796473112561e-08
+    6.377728138995419e-08
+    1.953866965847419e-07
+    4.703478363638027e-07
+ 6.57e+10    
+    4.700936064845114e-07
+    1.953815621438699e-07
+    4.548354081270768e-07
+    6.371989046239223e-08
+     1.26061295437447e-07
+    4.548100435164127e-07
+    3.015689751253572e-08
+    6.377120592277423e-08
+    1.954772409344625e-07
+    4.705069715837186e-07
+ 6.58e+10    
+    4.702531067162938e-07
+     1.95471908334801e-07
+    4.549518199609541e-07
+    6.371349484862489e-08
+    1.261146497888269e-07
+    4.549265186811591e-07
+    3.011572685162037e-08
+    6.376500729608324e-08
+    1.955677859068748e-07
+    4.706663009514971e-07
+ 6.59e+10    
+     4.70412801586206e-07
+    1.955622543550361e-07
+    4.550683511648722e-07
+    6.370697613472958e-08
+    1.261680012337965e-07
+    4.550431129864968e-07
+    3.007445343849479e-08
+    6.375868574927616e-08
+     1.95658331162709e-07
+    4.708258244389769e-07
+ 6.6e+10     
+    4.705726910669444e-07
+    1.956525998650492e-07
+    4.551850017671808e-07
+     6.37003345642924e-08
+    1.262213499193951e-07
+    4.551598264598299e-07
+    3.003307796561304e-08
+    6.375224152408963e-08
+    1.957488763625631e-07
+    4.709855420180875e-07
+ 6.61e+10    
+       4.707327751313e-07
+    1.957429445251853e-07
+    4.553017717966561e-07
+    6.369357038323646e-08
+     1.26274695993776e-07
+    4.552766591289932e-07
+    2.999160112773708e-08
+    6.374567486459132e-08
+     1.95839421166904e-07
+    4.711454536608481e-07
+ 6.62e+10    
+    4.708930537521562e-07
+    1.958332879956633e-07
+    4.554186612825031e-07
+    6.368668383981155e-08
+    1.263280396062042e-07
+    4.553936110222536e-07
+    2.995002362190559e-08
+    6.373898601716962e-08
+    1.959299652360679e-07
+    4.713055593393684e-07
+ 6.63e+10    
+    4.710535269024903e-07
+    1.959236299365752e-07
+    4.555356702543525e-07
+     6.36796751845831e-08
+    1.263813809070536e-07
+     4.55510682168308e-07
+    2.990834614740246e-08
+    6.373217523052242e-08
+    1.960205082302613e-07
+    4.714658590258498e-07
+ 6.64e+10    
+    4.712141945553729e-07
+    1.960139700078887e-07
+    4.556527987422636e-07
+    6.367254467042121e-08
+    1.264347200478058e-07
+    4.556278725962856e-07
+    2.986656940572502e-08
+     6.37252427556466e-08
+    1.961110498095618e-07
+    4.716263526925852e-07
+ 6.65e+10    
+    4.713750566839708e-07
+    1.961043078694465e-07
+    4.557700467767239e-07
+    6.366529255248974e-08
+    1.264880571810468e-07
+    4.557451823357465e-07
+    2.982469410055205e-08
+    6.371818884582683e-08
+    1.962015896339192e-07
+    4.717870403119587e-07
+ 6.66e+10    
+    4.715361132615449e-07
+    1.961946431809678e-07
+    4.558874143886465e-07
+    6.365791908823464e-08
+    1.265413924604648e-07
+    4.558626114166817e-07
+    2.978272093771138e-08
+    6.371101375662408e-08
+    1.962921273631561e-07
+    4.719479218564472e-07
+ 6.67e+10    
+    4.716973642614525e-07
+    1.962849756020497e-07
+    4.560049016093732e-07
+    6.365042453737272e-08
+    1.265947260408482e-07
+    4.559801598695124e-07
+    2.974065062514747e-08
+    6.370371774586465e-08
+    1.963826626569687e-07
+    4.721089972986205e-07
+ 6.68e+10    
+    4.718588096571463e-07
+     1.96375304792167e-07
+    4.561225084706717e-07
+    6.364280916188002e-08
+    1.266480580780823e-07
+    4.560978277250914e-07
+    2.969848387288847e-08
+     6.36963010736283e-08
+    1.964731951749281e-07
+    4.722702666111416e-07
+ 6.69e+10    
+    4.720204494221759e-07
+    1.964656304106743e-07
+    4.562402350047383e-07
+    6.363507322598013e-08
+    1.267013887291479e-07
+    4.562156150147023e-07
+    2.965622139301323e-08
+    6.368876400223675e-08
+    1.965637245764807e-07
+    4.724317297667661e-07
+ 6.7e+10     
+    4.721822835301881e-07
+    1.965559521168057e-07
+    4.563580812441961e-07
+    6.362721699613221e-08
+    1.267547181521183e-07
+    4.563335217700579e-07
+    2.961386389961796e-08
+     6.36811067962419e-08
+    1.966542505209488e-07
+    4.725933867383441e-07
+ 6.71e+10    
+    4.723443119549277e-07
+    1.966462695696767e-07
+    4.564760472220944e-07
+    6.361924074101901e-08
+    1.268080465061563e-07
+    4.564515480233024e-07
+    2.957141210878269e-08
+    6.367332972241376e-08
+    1.967447726675325e-07
+      4.7275523749882e-07
+ 6.72e+10    
+    4.725065346702366e-07
+    1.967365824282845e-07
+      4.5659413297191e-07
+    6.361114473153472e-08
+    1.268613739515126e-07
+    4.565696938070101e-07
+    2.952886673853746e-08
+    6.366543304972838e-08
+    1.968352906753096e-07
+     4.72917282021233e-07
+ 6.73e+10    
+    4.726689516500561e-07
+    1.968268903515093e-07
+    4.567123385275467e-07
+    6.360292924077271e-08
+    1.269147006495229e-07
+    4.566879591541863e-07
+    2.948622850882832e-08
+     6.36574170493557e-08
+    1.969258042032371e-07
+    4.730795202787168e-07
+ 6.74e+10    
+    4.728315628684266e-07
+    1.969171929981146e-07
+    4.568306639233353e-07
+    6.359459454401304e-08
+    1.269680267626048e-07
+    4.568063440982641e-07
+     2.94434981414831e-08
+     6.36492819946472e-08
+    1.970163129101515e-07
+    4.732419522445013e-07
+ 6.75e+10    
+     4.72994368299487e-07
+    1.970074900267492e-07
+    4.569491091940326e-07
+    6.358614091870983e-08
+    1.270213524542557e-07
+    4.569248486731084e-07
+    2.940067636017692e-08
+    6.364102816112318e-08
+    1.971068164547702e-07
+    4.734045778919113e-07
+ 6.76e+10    
+     4.73157367917478e-07
+    1.970977810959467e-07
+     4.57067674374823e-07
+    6.357756864447873e-08
+    1.270746778890505e-07
+    4.570434729130133e-07
+     2.93577638903975e-08
+    6.363265582646041e-08
+    1.971973144956924e-07
+     4.73567397194369e-07
+ 6.77e+10    
+    4.733205616967398e-07
+    1.971880658641277e-07
+     4.57186359501317e-07
+    6.356887800308397e-08
+    1.271280032326381e-07
+    4.571622168527023e-07
+    2.931476145941029e-08
+    6.362416527047928e-08
+    1.972878066913995e-07
+    4.737304101253929e-07
+ 6.78e+10    
+    4.734839496117134e-07
+    1.972783439896001e-07
+    4.573051646095511e-07
+    6.356006927842543e-08
+    1.271813286517394e-07
+    4.572810805273286e-07
+    2.927166979622335e-08
+    6.361555677513075e-08
+    1.973782927002565e-07
+    4.738936166585976e-07
+ 6.79e+10    
+    4.736475316369421e-07
+    1.973686151305603e-07
+    4.574240897359889e-07
+    6.355114275652549e-08
+    1.272346543141441e-07
+    4.574000639724747e-07
+     2.92284896315521e-08
+    6.360683062448362e-08
+     1.97468772180513e-07
+    4.740570167676974e-07
+ 6.8e+10     
+    4.738113077470716e-07
+    1.974588789450942e-07
+    4.575431349175204e-07
+      6.3542098725516e-08
+    1.272879803887086e-07
+    4.575191672241519e-07
+    2.918522169778378e-08
+    6.359798710471112e-08
+    1.975592447903036e-07
+     4.74220610426502e-07
+ 6.81e+10    
+    4.739752779168498e-07
+    1.975491350911777e-07
+    4.576623001914616e-07
+    6.353293747562476e-08
+    1.273413070453527e-07
+    4.576383903188012e-07
+    2.914186672894176e-08
+    6.358902650407785e-08
+    1.976497101876493e-07
+     4.74384397608922e-07
+ 6.82e+10    
+    4.741394421211282e-07
+    1.976393832266784e-07
+    4.577815855955544e-07
+     6.35236592991621e-08
+    1.273946344550572e-07
+    4.577577332932923e-07
+    2.909842546064971e-08
+    6.357994911292626e-08
+    1.977401680304585e-07
+    4.745483782889645e-07
+ 6.83e+10    
+    4.743038003348604e-07
+    1.977296230093556e-07
+    4.579009911679668e-07
+    6.351426449050726e-08
+    1.274479627898605e-07
+    4.578771961849234e-07
+    2.905489863009549e-08
+    6.357075522366324e-08
+    1.978306179765276e-07
+     4.74712552440738e-07
+ 6.84e+10    
+    4.744683525331077e-07
+    1.978198540968631e-07
+    4.580205169472939e-07
+    6.350475334609508e-08
+     1.27501292222857e-07
+    4.579967790314214e-07
+    2.901128697599505e-08
+    6.356144513074651e-08
+    1.979210596835423e-07
+    4.748769200384505e-07
+ 6.85e+10    
+    4.746330986910336e-07
+    1.979100761467482e-07
+    4.581401629725551e-07
+    6.349512616440145e-08
+    1.275546229281929e-07
+    4.581164818709424e-07
+    2.896759123855585e-08
+    6.355201913067068e-08
+    1.980114928090784e-07
+    4.750414810564081e-07
+ 6.86e+10    
+     4.74798038783908e-07
+    1.980002888164536e-07
+    4.582599292831957e-07
+    6.348538324593013e-08
+    1.276079550810642e-07
+    4.582363047420694e-07
+    2.892381215944052e-08
+    6.354247752195369e-08
+     1.98101917010603e-07
+    4.752062354690204e-07
+ 6.87e+10    
+    4.749631727871072e-07
+     1.98090491763319e-07
+    4.583798159190885e-07
+    6.347552489319823e-08
+    1.276612888577139e-07
+    4.583562476838162e-07
+    2.887995048172992e-08
+    6.353282060512272e-08
+    1.981923319454756e-07
+    4.753711832507965e-07
+ 6.88e+10    
+    4.751285006761134e-07
+     1.98180684644581e-07
+      4.5849982292053e-07
+    6.346555141072229e-08
+    1.277146244354282e-07
+     4.58476310735621e-07
+    2.883600694988648e-08
+    6.352304868270001e-08
+    1.982827372709484e-07
+    4.755363243763478e-07
+ 6.89e+10    
+    4.752940224265166e-07
+    1.982708671173756e-07
+    4.586199503282438e-07
+    6.345546310500397e-08
+    1.277679619925349e-07
+    4.585964939373537e-07
+    2.879198230971705e-08
+    6.351316205918892e-08
+    1.983731326441685e-07
+    4.757016588203881e-07
+ 6.9e+10     
+    4.754597380140151e-07
+    1.983610388387374e-07
+    4.587401981833774e-07
+    6.344526028451552e-08
+    1.278213017083991e-07
+    4.587167973293089e-07
+    2.874787730833578e-08
+    6.350316104105938e-08
+    1.984635177221779e-07
+    4.758671865577336e-07
+ 6.91e+10    
+     4.75625647414415e-07
+    1.984511994656028e-07
+     4.58860566527505e-07
+    6.343494325968569e-08
+    1.278746437634216e-07
+    4.588372209522109e-07
+    2.870369269412683e-08
+    6.349304593673371e-08
+    1.985538921619155e-07
+    4.760329075633039e-07
+ 6.92e+10    
+    4.757917506036318e-07
+    1.985413486548095e-07
+    4.589810554026256e-07
+    6.342451234288482e-08
+    1.279279883390349e-07
+    4.589577648472116e-07
+    2.865942921670694e-08
+    6.348281705657198e-08
+    1.986442556202173e-07
+    4.761988218121222e-07
+ 6.93e+10    
+    4.759580475576911e-07
+    1.986314860630985e-07
+    4.591016648511632e-07
+    6.341396784841024e-08
+    1.279813356177007e-07
+    4.590784290558889e-07
+    2.861508762688791e-08
+    6.347247471285755e-08
+    1.987346077538182e-07
+    4.763649292793171e-07
+ 6.94e+10    
+    4.761245382527288e-07
+    1.987216113471149e-07
+    4.592223949159673e-07
+    6.340331009247158e-08
+    1.280346857829067e-07
+    4.591992136202488e-07
+    2.857066867663884e-08
+    6.346201921978226e-08
+    1.988249482193529e-07
+    4.765312299401204e-07
+ 6.95e+10    
+    4.762912226649922e-07
+    1.988117241634093e-07
+    4.593432456403132e-07
+    6.339253939317591e-08
+    1.280880390191638e-07
+     4.59320118582726e-07
+    2.852617311904842e-08
+    6.345145089343167e-08
+     1.98915276673357e-07
+    4.766977237698714e-07
+ 6.96e+10    
+    4.764581007708409e-07
+    1.989018241684388e-07
+    4.594642170678997e-07
+    6.338165607051262e-08
+    1.281413955120027e-07
+    4.594411439861784e-07
+    2.848160170828701e-08
+     6.34407700517702e-08
+    1.990055927722681e-07
+    4.768644107440131e-07
+ 6.97e+10    
+    4.766251725467452e-07
+    1.989919110185678e-07
+     4.59585309242851e-07
+     6.33706604463385e-08
+    1.281947554479713e-07
+     4.59562289873895e-07
+    2.843695519956859e-08
+     6.34299770146261e-08
+    1.990958961724268e-07
+    4.770312908380978e-07
+ 6.98e+10    
+    4.767924379692911e-07
+    1.990819843700705e-07
+    4.597065222097181e-07
+    6.335955284436253e-08
+    1.282481190146313e-07
+    4.596835562895891e-07
+    2.839223434911274e-08
+    6.341907210367652e-08
+    1.991861865300789e-07
+    4.771983640277836e-07
+ 6.99e+10    
+    4.769598970151775e-07
+    1.991720438791309e-07
+    4.598278560134738e-07
+    6.334833359013072e-08
+    1.283014864005552e-07
+    4.598049432774023e-07
+     2.83474399141064e-08
+    6.340805564243213e-08
+    1.992764635013754e-07
+    4.773656302888371e-07
+ 7e+10       
+    4.771275496612187e-07
+    1.992620892018445e-07
+    4.599493106995181e-07
+    6.333700301101069e-08
+    1.283548577953231e-07
+    4.599264508819013e-07
+    2.830257265266555e-08
+    6.339692795622215e-08
+    1.993667267423742e-07
+    4.775330895971331e-07
* NOTE: Solution at 1e+08 Hz used as DC point.

.model g_m4lines_HFSS_W_1 sp N=4 SPACING=nonuniform VALTYPE=real
+ INTERPOLATION=spline
+ DATA = 700
+ 0           
+    0.0008510784137774075
+   -0.0001574885068096611
+    0.0008545778793345019
+   -1.126766962080041e-06
+   -6.750040879516493e-05
+    0.0008550095139155642
+    1.916452937783147e-07
+   -1.124233049329695e-06
+   -0.0001577728606750277
+    0.0008493537729414312
+ 2e+08       
+     0.001771925943544663
+   -0.0003422192817968613
+     0.001783399601946027
+   -1.914479231735113e-06
+   -0.0001439836006190334
+     0.001784884906339565
+   -6.883795793363981e-07
+   -1.813070534314566e-06
+   -0.0003453609017088446
+     0.001767794398634545
+ 3e+08       
+     0.002589167663714148
+   -0.0004862325620218706
+     0.002602172368458493
+    -4.24264201150778e-06
+   -0.0002051949894804335
+     0.002603649703392652
+   -1.940403693732582e-07
+   -4.204261684875072e-06
+   -0.0004883451826726586
+     0.002583267608278901
+ 4e+08       
+     0.003410105892792772
+   -0.0006320826667550488
+     0.003424593582586204
+     -5.1603471438556e-06
+   -0.0002692968407564275
+     0.003426344206001315
+    5.596352698386012e-07
+   -5.145223856449713e-06
+   -0.0006336447058186832
+     0.003402965625411628
+ 5e+08       
+     0.004251253720891197
+   -0.0007859891797900177
+     0.004268388482517638
+   -5.531784450129825e-06
+   -0.0003363604182242495
+     0.004270538996314664
+    1.186565496963342e-06
+   -5.519217064341381e-06
+   -0.0007874793443164447
+     0.004242635950122304
+ 6e+08       
+     0.005100762312396182
+   -0.0009430014308700359
+     0.005121210927044995
+   -6.066091067623449e-06
+   -0.0004039347148926231
+     0.005123776599907521
+     1.67805249550687e-06
+   -6.051272278310955e-06
+   -0.0009446545702791783
+     0.005090428624025207
+ 7e+08       
+     0.005949399036259124
+     -0.00109962973832101
+     0.005973202478298719
+   -6.900387855348104e-06
+   -0.0004708633623819473
+     0.005976190203725119
+     2.12850066081404e-06
+   -6.883330585852565e-06
+    -0.001101564261166545
+     0.005937328260258257
+ 8e+08       
+     0.006794944394096883
+    -0.001255145629963329
+     0.006821879978445718
+   -7.853925401216596e-06
+   -0.0005371624762598283
+     0.006825307379807402
+    2.624896992374523e-06
+   -7.835220263012374e-06
+    -0.001257412333507148
+     0.006781220521678108
+ 9e+08       
+     0.007639961161126815
+    -0.001410465549404944
+     0.007669958032171864
+   -8.650914985511579e-06
+   -0.0006034038777395368
+     0.007673828728046199
+    3.223908515412809e-06
+   -8.630619741544247e-06
+    -0.001413048983927965
+     0.007624599633091086
+ 1e+09       
+     0.008489164179541578
+    -0.001567089680793842
+     0.008522596763779127
+    -9.03333658169665e-06
+   -0.0006702837516171617
+     0.008526868098619748
+    3.958713626491957e-06
+   -9.010999740784024e-06
+    -0.001569901800190448
+     0.008471994312932428
+ 1.1e+09     
+     0.009365240377547138
+    -0.001722266892223308
+     0.009404256167478054
+   -9.423266663160531e-06
+   -0.0007857177301352359
+     0.009410139247021816
+    1.205728962055263e-05
+   -8.863825249618031e-06
+    -0.001727516837899321
+     0.009350418670556184
+ 1.2e+09     
+      0.01027358581207574
+    -0.001893766827112009
+      0.01031918129761795
+   -1.098712930394506e-05
+   -0.0009043907792473753
+       0.0103266333565252
+    2.188845267251413e-05
+   -9.851738114845894e-06
+    -0.001901318689218514
+      0.01026077554425189
+ 1.3e+09     
+      0.01120508314273132
+    -0.002077491652537177
+      0.01125805886864822
+   -1.358148729716694e-05
+     -0.00102445548700732
+      0.01126701656795569
+    3.312220396494996e-05
+   -1.186571235826012e-05
+    -0.002087187188230752
+      0.01119391251952879
+ 1.4e+09     
+      0.01215177503188965
+     -0.00226975982073262
+      0.01221275621035362
+   -1.701266719404887e-05
+    -0.001144423134243082
+      0.01222314154416545
+    4.542182774441917e-05
+   -1.473678286565219e-05
+    -0.002281429018654841
+      0.01214185436760519
+ 1.5e+09     
+      0.01310689786897508
+    -0.002467384346829484
+      0.01317634824390623
+   -2.106901166756732e-05
+    -0.001263102881715434
+      0.01318807342383928
+    5.846253322731964e-05
+    -1.82699682389388e-05
+    -0.002480853150292131
+      0.01309783379920386
+ 1.6e+09     
+      0.01406484794301911
+    -0.002667687929676103
+      0.01414308072944281
+   -2.554112832261454e-05
+    -0.001379554788594624
+        0.014156052147932
+     7.19426945193532e-05
+   -2.226632781937273e-05
+    -0.002682783689278925
+      0.01405625463486187
+ 1.7e+09     
+      0.01502110336915699
+     -0.00286848094739762
+       0.0151082914484777
+    -3.02337158262647e-05
+    -0.001493051502216864
+      0.01512241284049648
+    8.559001087671191e-05
+    -2.65364066837319e-05
+    -0.002885036121207663
+      0.01501261090348283
+ 1.8e+09     
+       0.0159721199600859
+    -0.003068019440043474
+      0.01606830642232875
+   -3.497173732576632e-05
+    -0.001603045708648557
+      0.01608348134049752
+    9.916426663530168e-05
+   -3.090772712410484e-05
+    -0.003085873970501822
+      0.01596338019202186
+ 1.9e+09     
+      0.01691521466932164
+    -0.003264953975040904
+         0.01702032410361
+   -3.960295056036582e-05
+    -0.001709141791717847
+      0.01703645781122268
+     0.000112457862774526
+   -3.522833235378051e-05
+    -0.003283956684190661
+      0.01690590494409298
+ 2e+09       
+      0.01784844637676117
+    -0.003458276126291491
+      0.01796229690213946
+   -4.399819143089473e-05
+    -0.001811070899646675
+      0.01797929777804945
+    0.0001252949242323399
+   -3.936782032214778e-05
+    -0.003478285396460204
+      0.01783827150068856
+ 2.1e+09     
+      0.01877050065594481
+     -0.00364726656306578
+      0.01889281646706835
+    -4.80503512050122e-05
+    -0.001908668996931689
+      0.01891059700671141
+    0.0001375295312901009
+   -4.321686100640197e-05
+    -0.003668150510027718
+      0.01875919350964359
+ 2.2e+09     
+      0.01968058271073447
+    -0.003831446971078448
+      0.01981100682162004
+   -5.167266269621122e-05
+    -0.002001857646109308
+       0.0198294843094085
+    0.0001490434485531878
+   -4.668586288669578e-05
+    -0.003853083268935076
+      0.01966790385551422
+ 2.3e+09     
+      0.02057832081937954
+     -0.00401053689133327
+      0.02071642767609169
+   -5.479668664406901e-05
+    -0.002090627321437817
+      0.02073552459560022
+    0.0001597436058387994
+   -4.970322194290514e-05
+    -0.004032812370404358
+      0.02056405739895874
+ 2.4e+09     
+       0.0214636812838417
+    -0.004184415846709998
+      0.02160898895021911
+   -5.737023836009596e-05
+    -0.002175023064360656
+      0.02162863318985807
+    0.0001695595033189767
+   -5.221342618520947e-05
+    -0.004207225955553296
+      0.02144764546992921
+ 2.5e+09     
+      0.02233689495635542
+    -0.004353090689305508
+      0.02248887663271251
+    -5.93553946562198e-05
+    -0.002255132281685338
+      0.02250900153604074
+     0.000178440656178024
+   -5.417518049834463e-05
+    -0.004376338888019506
+      0.02231892213416952
+ 2.6e+09     
+      0.02319839481315557
+    -0.004516667848678325
+      0.02335648951129803
+   -6.072665607595494e-05
+    -0.002331074477905164
+      0.02337703381296798
+    0.0001863541537430118
+   -5.555964494840214e-05
+    -0.004540264981725635
+      0.02317834165517049
+ 2.7e+09     
+      0.02404876368700916
+    -0.004675330029038036
+       0.0242123859466545
+   -6.146929811250018e-05
+    -0.002402992709637334
+      0.02423329362742856
+    0.0001932823793092931
+   -5.634883327072261e-05
+    -0.004699193711053706
+      0.02402650622203943
+ 2.8e+09     
+      0.02488869108829252
+    -0.004829316849272676
+      0.02505723967499358
+   -6.157791953034413e-05
+    -0.002471046554295416
+       0.0250784597624932
+    0.0001992209163112054
+    -5.65341889054642e-05
+    -0.004853370885958032
+      0.02486412283909217
+ 2.9e+09     
+      0.02571893798471482
+     -0.00497890891448334
+      0.02589180355534933
+   -6.105518071652474e-05
+    -0.002535406395985167
+      0.02591328989129596
+    0.0002041766518207992
+   -5.611533800633508e-05
+    -0.005003082772111882
+      0.02569196822040123
+ 3e+09       
+      0.02654030843057249
+    -0.005124414831741709
+      0.02671688018888572
+   -5.991071653041316e-05
+    -0.002596248847434945
+      0.02673859117859712
+    0.0002081660780411611
+   -5.509900842038426e-05
+    -0.005148643162484806
+      0.02651086055970409
+ 3.1e+09     
+      0.02735362700647446
+    -0.005266160722923767
+      0.02753329839861923
+   -5.816020395380855e-05
+    -0.002653753145652403
+      0.02755519675440199
+    0.0002112137853879599
+   -5.349809807284262e-05
+    -0.005290382948681832
+       0.0273216371216105
+ 3.2e+09     
+      0.02815972112745218
+     -0.00540448183502547
+      0.02834189464708476
+   -5.582456334206602e-05
+    -0.002708098379288795
+      0.02836394713384759
+    0.0002133511361060742
+   -5.133087370685159e-05
+    -0.005428641789331289
+      0.02812513670151764
+ 3.3e+09     
+      0.02895940738582068
+    -0.005539715897779149
+      0.02914349857143562
+   -5.292927217311518e-05
+    -0.002759461426106182
+      0.02916567576024055
+    0.0002146151045286214
+   -4.862028033594562e-05
+    -0.005563761523296067
+      0.02892218611365642
+ 3.4e+09     
+      0.02975348120491277
+    -0.005672197926265376
+      0.02993892192008673
+   -4.950377119089478e-05
+    -0.002808015498559527
+      0.02996119795335504
+    0.0002150472685775968
+   -4.539334228734866e-05
+    -0.005696081024162277
+      0.02971358997917103
+ 3.5e+09     
+      0.03054270918454387
+    -0.005802256210619414
+      0.03072895027584877
+   -4.558094430274699e-05
+    -0.002853929213707344
+      0.03075130264644053
+    0.0002146929365604516
+    -4.16806378442724e-05
+    -0.005825932237447606
+      0.03050012319287979
+ 3.6e+09     
+      0.03132782361519434
+    -0.005930209274906457
+       0.0315143370437994
+    -4.11966552474558e-05
+    -0.002897366120062069
+      0.03153674638909023
+    0.0002136003934513309
+   -3.751583092252968e-05
+    -0.005953637182357517
+       0.0312825255449273
+ 3.7e+09     
+      0.03210951872371821
+    -0.006056363622458887
+      0.03229579926598097
+   -3.638932574895624e-05
+    -0.002938484628346175
+      0.03231824917728614
+    0.0002118202514428352
+   -3.293524475659194e-05
+    -0.006079505735412627
+      0.03206149806032708
+ 3.8e+09     
+      0.03288844828842345
+    -0.006181012115497719
+      0.03307401489873355
+   -3.119954153644479e-05
+    -0.002977438305277276
+      0.03309649174589871
+    0.0002094048904512994
+   -2.797746412765189e-05
+    -0.006203834043973792
+      0.03283770069505192
+ 3.9e+09     
+      0.03366522432593198
+    -0.006304432862993208
+      0.03384962125216794
+   -2.566967422656713e-05
+    -0.003014376499337106
+      0.03387211402279833
+    0.0002064079753370875
+    -2.26829542073325e-05
+    -0.006326903443923064
+       0.0336117510922465
+ 4e+09       
+      0.03444041660705933
+    -0.006426888512868241
+      0.03462321434552248
+   -1.984350864853157e-05
+    -0.003049445274841402
+      0.03464571449810941
+     0.000202884037777293
+    -1.70936856262586e-05
+    -0.006448979777951346
+      0.03438422415713679
+ 4.1e+09     
+      0.03521455280503739
+    -0.006548625863273356
+      0.03539534897773616
+   -1.376586679868424e-05
+    -0.003082788635327055
+      0.03541785030781897
+     0.000198888111945822
+    -1.12527569492496e-05
+    -0.006570313029535196
+      0.03515565225533099
+ 4.2e+09     
+      0.03598811911779282
+    -0.006669875723224587
+      0.03616653935039939
+    -7.48222130944132e-06
+    -0.003114550019050932
+      0.03618903786884654
+    0.0001944754143812919
+   -5.204007415423499e-06
+    -0.006691137203228396
+      0.03592652587754672
+ 4.3e+09     
+      0.03676156123773796
+    -0.006790852965834956
+      0.03693726011121552
+   -1.038293196122897e-06
+    -0.003144874047921431
+      0.03695975393369288
+    0.0001897010596396189
+    1.008385333896994e-06
+    -0.006811670394798404
+      0.03669729464543964
+ 4.4e+09     
+      0.03753528556861304
+    -0.006911756728085977
+      0.03770794771105323
+    5.520369198262689e-06
+    -0.003173908506072943
+      0.03773043695775746
+     0.000184619804531333
+    7.340325669106694e-06
+    -0.006932115005408823
+      0.03746836855915953
+ 4.5e+09     
+      0.03830966061023246
+     -0.00703277071993447
+      0.03847900198736422
+    1.214883060730594e-05
+    -0.003201806515140816
+      0.03850148869211994
+    0.0001792858149376997
+    1.374823913048782e-05
+    -0.007052658062849524
+      0.03824011940842812
+ 4.6e+09     
+      0.03908501844931703
+    -0.007154063612841361
+      0.03925078790185312
+    1.880322614403114e-05
+    -0.003228728859742837
+      0.03927327592969865
+    0.0001737524503931347
+    2.018952793903699e-05
+    -0.007173471620058344
+      0.03901288228611935
+ 4.7e+09     
+      0.03986165630862881
+    -0.007275789483810718
+      0.04002363737144016
+    2.544122952743343e-05
+    -0.003254846398518356
+      0.04004613234384806
+    0.0001680720628227935
+    2.662303694660152e-05
+    -0.007294713207131516
+      0.03978695715721735
+ 4.8e+09     
+      0.04063983811794344
+    -0.007398088295963741
+      0.04079785113931124
+    3.202252219415577e-05
+      -0.0032803424734062
+      0.04082036036620797
+    0.0001622958070374384
+    3.300952005008293e-05
+    -0.007416526317911974
+      0.04056261044722113
+ 4.9e+09     
+      0.04141979607948782
+    -0.007521086400731428
+      0.04157370063777268
+    3.850924871641906e-05
+     -0.00330541520322601
+      0.04159623305553259
+    0.0001564734618064254
+    3.931209255591574e-05
+     -0.00753904091626189
+      0.04134007662304314
+ 5e+09       
+      0.04220173220775175
+    -0.007644897050086832
+      0.04235142979731701
+    4.486643910290691e-05
+    -0.003330279518324451
+      0.04237399591190392
+     0.000150653261531544
+    4.549665013841523e-05
+    -0.007662373950425647
+      0.04211955974663219
+ 5.1e+09     
+      0.04298581982937297
+    -0.007769620909974465
+      0.04313125675743106
+    5.106237372474253e-05
+    -0.003355168763232237
+      0.04315386859185737
+    0.0001448817396854025
+     5.15322302033455e-05
+    -0.007786629866593876
+      0.04290123498725861
+ 5.2e+09     
+      0.04377220503337659
+    -0.007895346568330398
+       0.0439133754350427
+    5.706886226780619e-05
+    -0.003380335667221548
+      0.04393604648029603
+    0.0001392035861875824
+    5.739128712945645e-05
+    -0.007911901114984384
+      0.04368525008290714
+ 5.3e+09     
+      0.04456100806562334
+    -0.008022151032891903
+      0.04469795690702939
+    6.286140492985345e-05
+    -0.003406052462803893
+      0.04472070207559622
+    0.0001336615216707136
+    6.304984968105829e-05
+     -0.00803826864353803
+      0.04447172674474176
+ 5.4e+09     
+      0.04535232466405426
+    -0.008150100215423931
+      0.04548515056496469
+    6.841920288400431e-05
+    -0.003432609925074866
+      0.04550798614604779
+    0.0001282961920121089
+     6.84875276910728e-05
+    -0.008165802375732863
+      0.04526076200128947
+ 5.5e+09     
+      0.04614622733333946
+    -0.008279249400077742
+      0.04627508500438419
+    7.372498674901377e-05
+    -0.003460315116567516
+      0.04629802861987575
+    0.0001231460864333892
+    7.368733683640427e-05
+    -0.008294561670091606
+      0.04605242948097246
+ 5.6e+09     
+      0.04694276655893637
+    -0.008409643694368458
+      0.04706786861839184
+    7.876463735368022e-05
+    -0.003489487658979101
+      0.04709093917862448
+    0.0001182474817617296
+    7.863531587858378e-05
+    -0.008424595759713877
+      0.04684678063298782
+ 5.7e+09     
+      0.04774197196142031
+    -0.008541318461735488
+      0.04786358987726221
+    8.352658317844751e-05
+     -0.00352045441957497
+      0.04788680753551447
+    0.0001136344139931951
+    8.331992084240764e-05
+    -0.008555944170630318
+      0.04764384588736566
+ 5.8e+09     
+      0.04854385339233939
+    -0.008674299734854809
+      0.04866231729221764
+    8.800097380111589e-05
+    -0.003553542598275248
+      0.04868570339690814
+    0.0001093386760579192
+    8.773119555407225e-05
+    -0.008688637117973273
+      0.04844363575541112
+ 5.9e+09     
+      0.04934840197284134
+    -0.008808604608839707
+      0.04946409908247976
+    9.217864810670328e-05
+    -0.003589071329085415
+       0.0494876761259367
+    0.0001053898377191126
+    9.185973739849352e-05
+    -0.008822695878919772
+      0.04924614187171852
+ 6e+09       
+      0.05015559107601822
+    -0.008944241613248539
+      0.05026896258880111
+    9.604993872756683e-05
+    -0.003627342058692736
+      0.05029275415144966
+    0.0001018152800377145
+    9.569549986763798e-05
+    -0.008958133141141555
+      0.05005133797863487
+ 6.1e+09     
+      0.05096537725342531
+    -0.009081211061485156
+      0.05107691350178677
+    9.960337800514658e-05
+    -0.003668628121597061
+      0.05110094419055325
+    9.864023314378747e-05
+    9.922649730407141e-05
+    -0.009094953325161605
+      0.05085918085355693
+ 6.2e+09     
+      0.05177770110568441
+    -0.009219505375819991
+      0.05188793499636234
+    0.0001028243927309124
+    -0.003713164075518574
+      0.05191223037605126
+    9.588780264572854e-05
+    0.0001024374992187409
+    -0.009233152878658973
+      0.05166961117889519
+ 6.3e+09     
+      0.05259248809662359
+    -0.009359109385981772
+      0.05270198688116731
+    0.0001056940915753068
+    -0.003761135470312672
+      0.05272657339752819
+     9.35789674241965e-05
+    0.0001053088182237027
+    -0.009372720540484497
+      0.05248255435407902
+ 6.4e+09     
+      0.05340964931015848
+    -0.009500000599164407
+      0.05351900487999077
+    0.0001081882570927563
+    -0.003812669776132892
+      0.05354390977315068
+    9.173253032921085e-05
+    0.0001078153036125941
+    -0.009513637572045786
+      0.05329792124873011
+ 6.5e+09     
+      0.05422908214919382
+    -0.009642149439444652
+      0.05433890015898076
+    0.0001102766509483789
+    -0.003867829175314569
+      0.05436415136588001
+    9.036500382729852e-05
+    0.0001099256493942086
+    -0.009655877953869362
+       0.0541156088962049
+ 6.6e+09     
+       0.0550506709762635
+    -0.009785519455046344
+      0.05516155919716047
+    0.0001119227254883009
+    -0.003926605820384631
+      0.05518718524158849
+    8.949041509812602e-05
+    0.0001116021100783138
+    -0.009799408545587456
+      0.05493550112714396
+ 6.7e+09     
+      0.05587428769641289
+    -0.009930067492608019
+      0.05598684406970772
+    0.0001130838078587801
+    -0.003988919983514335
+      0.05601287393849481
+    8.912001931632722e-05
+    0.0001128006906155675
+    -0.009944189208317907
+      0.05575746914345731
+ 6.8e+09     
+      0.05669979228387809
+     -0.01007574383854498
+      0.05681459317650969
+    0.0001137117874660383
+    -0.004054621289616338
+      0.05684105618038499
+    8.926191541864365e-05
+    0.0001134718415010281
+     -0.01009017288933805
+      0.05658137203422099
+ 6.9e+09     
+      0.05752703325529138
+     -0.01022249232863571
+       0.0576446224073737
+    0.0001137542981576765
+    -0.004123492965688367
+      0.05767154802495507
+     8.99205648409679e-05
+    0.0001135616506616668
+     -0.01023730566999354
+      0.05740705723613764
+ 7e+09       
+      0.05835584809326538
+     -0.01037025042797262
+      0.05847672669546109
+    0.0001131563483854286
+    -0.004195258787687191
+      0.05850414439879372
+    9.109621968326391e-05
+    0.0001130134856492482
+     -0.01038552677879577
+      0.05823436094234004
+ 7.1e+09     
+      0.05918606362513353
+     -0.01051894928426954
+      0.05931068187727106
+     0.000111862320834393
+    -0.004269592196449753
+       0.0593386209372835
+    9.278427172779873e-05
+    0.0001117700079071833
+      -0.0105347685725194
+      0.05906310846424067
+ 7.2e+09     
+      0.06001749636220865
+     -0.01066851375811188
+      0.06014624675485599
+    0.0001098182414366729
+    -0.004346126911401301
+      0.06017473602505715
+    9.497453709194433e-05
+    0.0001097754593339557
+     -0.01068495648871345
+      0.05989311455172049
+ 7.3e+09     
+      0.06084995280511461
+     -0.01081886243401343
+      0.06098316524599482
+    0.0001069742083346579
+    -0.004424468308269198
+      0.06101223292269104
+    9.765049272682409e-05
+    0.0001069781120337258
+     -0.01083600897333137
+      0.06072418367714527
+ 7.4e+09     
+      0.06168322972054284
+     -0.01096990761610606
+      0.06182116851073617
+     0.000103286874169359
+    -0.004504204844482509
+      0.06185084186801239
+    0.0001007884804871547
+    0.0001033327749747617
+     -0.01098783738716352
+      0.06155611028850152
+ 7.5e+09     
+      0.06251711439424903
+     -0.01112155531197719
+      0.06265997695612448
+    9.872188818187388e-05
+     -0.00458491890121797
+      0.06269028205380203
+    0.0001043568923901829
+    9.880326440903347e-05
+     -0.01114034589446468
+      0.06238867903641124
+ 7.6e+09     
+      0.06335138486433239
+     -0.01127370520766319
+      0.06349930204184366
+    9.325622495431169e-05
+    -0.004666196543958371
+      0.06353026340461151
+    0.0001083153474377395
+    9.336476526450093e-05
+     -0.01129343133668754
+      0.06322166497902189
+ 7.7e+09     
+      0.06418581013795863
+     -0.01142625063619657
+      0.06433884783425589
+    8.688035061374063e-05
+    -0.004747635860539773
+       0.0643704881001588
+    0.0001126138665573382
+    8.700603473960284e-05
+      -0.0114469830936475
+      0.06405483376788973
+ 7.8e+09     
+      0.06502015039378924
+     -0.01157907854147542
+      0.06517831228137018
+    7.960020160914765e-05
+    -0.004828853694820438
+      0.06521065181784455
+    0.0001171920483561233
+    7.973142363722555e-05
+     -0.01160088293384654
+      0.06488794181708933
+ 7.9e+09     
+      0.06585415717157481
+     -0.01173206943865094
+      0.06601738820386296
+    7.143897306065294e-05
+    -0.004909490737639595
+      0.06605044468952292
+    0.0001219782448985403
+    7.156271288723953e-05
+     -0.01175500485514074
+         0.06572073645698
+ 8e+09       
+       0.0666875735496964
+     -0.01188509737175428
+      0.06685576401556297
+    6.243873142236219e-05
+    -0.004989215053119181
+      0.06688955198597121
+    0.0001268887338896306
+     6.25407804722266e-05
+     -0.01190921491649779
+      0.06655295607340019
+ 8.1e+09     
+      0.06752013431093691
+     -0.01203802986893642
+      0.06769312419998215
+     5.26618789935172e-05
+    -0.005067724202307853
+      0.06772765455567858
+    0.0001318268815974095
+    5.272712678841118e-05
+     -0.01206337106127721
+      0.06738433023256341
+ 8.2e+09     
+      0.06835156609642565
+     -0.01219072789547175
+      0.06852914957751499
+    4.219250565831105e-05
+    -0.005144746177665587
+      0.06856442905263356
+    0.0001366822895791837
+     4.22052943444837e-05
+     -0.01221732293228379
+      0.06821457979160576
+ 8.3e+09     
+      0.06918158754751333
+     -0.01234304580456699
+       0.0693635174014342
+    3.113766670129279e-05
+    -0.005220039384664501
+      0.06939954799130822
+    0.0001413299176990295
+    3.108222119228106e-05
+     -0.01237091167877495
+      0.06904341699455294
+ 8.4e+09     
+      0.07000990943526032
+     -0.01249483128599927
+      0.07019590132070823
+    1.962862551864751e-05
+    -0.005293391906663178
+        0.070232679666949
+    0.0001456291758976692
+    1.948956748174706e-05
+     -0.01252396975563034
+      0.06987054555341771
+ 8.5e+09     
+      0.07083623477724274
+     -0.01264592531265572
+      0.07102597124497613
+    7.822097515599918e-06
+    -0.005364620272708447
+      0.07106348797661048
+    0.0001494229775465432
+    7.585052026513363e-06
+     -0.01267632071498615
+      0.07069566071416773
+ 8.6e+09     
+      0.07166025894144809
+     -0.01279616208513739
+      0.07185339314271851
+   -4.098472617140533e-06
+    -0.005433567921199902
+      0.07189163217208995
+    0.0001525367478384888
+   -4.446168307189764e-06
+     -0.01282777899077784
+      0.07151844930738668
+ 8.7e+09     
+       0.0724816697371387
+     -0.01294536897470282
+      0.07267782879858722
+   -1.592157292931419e-05
+    -0.005500103520631428
+      0.07271676657085868
+    0.0001547773814144153
+   -1.639004842824386e-05
+     -0.01297814967679944
+       0.0723385897835693
+ 8.8e+09     
+      0.07330014749266985
+     -0.01309336646494316
+      0.07349893555061932
+   -2.740620326969849e-05
+    -0.005564119275885217
+      0.07353854024587266
+    0.0001559321442053503
+   -2.800211113330748e-05
+     -0.01312722829906113
+      0.07315575223311499
+ 8.9e+09     
+      0.07411536512035602
+     -0.01323996809269175
+       0.0743163660231092
+   -3.828035391473256e-05
+    -0.005625529317560036
+      0.07435659671021014
+    0.0001557675152174239
+   -3.900579136176035e-05
+      -0.0132748005833965
+      0.07396959839120701
+ 9e+09       
+      0.07492698816857342
+      -0.0133849803887681
+      0.07512976786650874
+   -4.823937061988325e-05
+    -0.005684268244238754
+      0.07517057360809958
+    0.0001540279646660985
+   -4.909065475012554e-05
+     -0.01342064221942946
+      0.07477978162787444
+ 9.1e+09     
+      0.07573467486136153
+      -0.0135282028192344
+      0.07593878351198866
+   -5.694419665038013e-05
+    -0.005740289864259162
+      0.07598010242019369
+    0.0001504346654577647
+    -5.79104803341661e-05
+     -0.01356451862215576
+      0.07558594692362579
+ 9.2e+09     
+       0.0765380761258443
+     -0.01366942772790385
+      0.07674304994527163
+   -6.401948541650925e-05
+    -0.005793566164633837
+      0.07678480818793591
+    0.0001446841355194086
+   -6.508120030677836e-05
+     -0.01370618469251933
+      0.07638773083111923
+ 9.3e+09     
+      0.07733683560783229
+     -0.01380844028087824
+       0.0775421985019821
+   -6.905157981164204e-05
+    -0.005844086520048032
+      0.07758430925953401
+    0.0001364468088985602
+   -7.017869220700889e-05
+     -0.01384538457847529
+      0.07718476142339242
+ 9.4e+09     
+      0.07813058967598839
+     -0.01394501841391585
+      0.07833585468500061
+   -7.158635630386646e-05
+    -0.005891857143884822
+      0.07837821705831416
+    0.0001253655339099895
+    -7.27364208683379e-05
+     -0.01398185143812279
+       0.0779766582292182
+ 9.5e+09     
+       0.0789189674149563
+      -0.0140789327834338
+      0.07912363800304285
+   -7.112693335917068e-05
+      -0.0059369007754087
+      0.07916613587299422
+    0.0001110539969093097
+   -7.224292898544383e-05
+     -0.01411530720656916
+       0.0787630321561832
+ 9.6e+09     
+      0.07970159060784765
+     -0.01420994672193901
+      0.07990516182884204
+   -6.713124497152359e-05
+    -0.005979256591989042
+      0.07994766266859411
+    9.309507054471684e-05
+   -6.813917636707204e-05
+     -0.01424546236824982
+      0.07954348540211048
+ 9.7e+09     
+       0.0804780737084855
+     -0.01433781619865664
+        0.080680033274781
+   -5.900948103674321e-05
+    -0.006018980331996954
+      0.08072238691619553
+    7.103908559336286e-05
+   -5.981572892117858e-05
+     -0.01437201573647566
+       0.0803176113554622
+ 9.8e+09     
+      0.08124802380378797
+     -0.01446228978608608
+      0.08144785308353972
+   -4.612139711545482e-05
+    -0.006056144612268973
+      0.08148989043951198
+    4.440202574462477e-05
+    -4.66097992518357e-05
+     -0.01449465424201697
+      0.08108499448537031
+ 9.9e+09     
+      0.08201104056667137
+     -0.01458310863316487
+      0.08220821553121899
+   -2.777349685838151e-05
+    -0.006090839423373145
+      0.08224974727614504
+    1.266364496297018e-05
+   -2.780214150908695e-05
+     -0.01461305273255238
+      0.08184521022195509
+ 1e+10       
+      0.08276671619984004
+      -0.0147000064456568
+      0.08296070834041837
+   -3.216091076274673e-06
+    -0.006123172785997904
+      0.08300152355145053
+   -2.473449263825115e-05
+   -2.613803885043002e-06
+     -0.01472687378482095
+      0.08259782482760331
+ 1.01e+10    
+      0.08358103488630225
+     -0.01483754692766492
+       0.0837868708752173
+   -5.131704652226775e-06
+     -0.00619975142264406
+      0.08381973709464782
+   -3.078811604518899e-05
+   -4.901673887094428e-06
+     -0.01486324361076061
+      0.08341116781724983
+ 1.02e+10    
+       0.0843951054542099
+     -0.01497498698539517
+      0.08461123386058836
+    -7.19015564050495e-06
+    -0.006275369116238049
+      0.08463685285560454
+   -3.693712015043638e-05
+   -7.307883775140543e-06
+     -0.01499964398118805
+      0.08422425136508603
+ 1.03e+10    
+      0.08520888641009869
+     -0.01511233074322629
+      0.08543385084343005
+   -9.392881922643415e-06
+    -0.006350057796906667
+      0.08545288295870682
+    -4.31852493535073e-05
+   -9.835105329059415e-06
+     -0.01513607083991632
+      0.08503703304518799
+ 1.04e+10    
+      0.08602233850201152
+     -0.01524958213112529
+       0.0862547739355793
+   -1.174139443390536e-05
+     -0.00642384849193948
+      0.08626784018330433
+   -4.953619126085045e-05
+   -1.248602227462044e-05
+     -0.01527252035821899
+      0.08584947276288489
+ 1.05e+10    
+      0.08683542463776751
+     -0.01538674489166767
+      0.08707405381700487
+   -1.423726730757544e-05
+    -0.006496771351633519
+      0.08708173787273572
+   -5.599357279717021e-05
+   -1.526332322794501e-05
+     -0.01540898892283817
+      0.08666153266843797
+ 1.06e+10    
+      0.08764810980501586
+     -0.01552382258721446
+      0.08789173974280388
+   -1.688212860654465e-05
+    -0.006568855674316229
+      0.08789458985059012
+   -6.256095647759388e-05
+   -1.816969512547255e-05
+     -0.01554547312482846
+      0.08747317707266003
+ 1.07e+10    
+      0.08846036099309927
+     -0.01566081860718187
+      0.08870787955353784
+   -1.967765161712328e-05
+    -0.006640129930578985
+      0.08870641034370982
+    -6.92418368443172e-05
+   -2.120781711309385e-05
+     -0.01568196974916722
+      0.08828437236449665
+ 1.08e+10    
+      0.08927214711674922
+     -0.01579773617534824
+      0.08952251968848646
+   -2.262554667381783e-05
+    -0.006710621786753763
+      0.08951721391146596
+   -7.603963707297203e-05
+   -2.438035486605544e-05
+     -0.01581847576506778
+      0.08909508693059248
+ 1.09e+10    
+      0.09008343894162638
+     -0.01593457835714943
+      0.09033570520144067
+   -2.572755349147294e-05
+    -0.006780358127662104
+      0.09032701538087343
+   -8.295770575074456e-05
+   -2.768995531635902e-05
+     -0.01595498831693756
+      0.08990529107685323
+ 1.1e+10     
+      0.09089420901171812
+     -0.01607134806692177
+      0.09114747977869091
+    -2.89854339768083e-05
+    -0.006849365078664941
+      0.09113582978713305
+   -8.999931382892195e-05
+   -3.113924176423874e-05
+     -0.01609150471592748
+      0.09071495695201523
+ 1.11e+10    
+      0.09170443157859663
+      -0.0162080480750561
+      0.09195788575890072
+   -3.240096549963762e-05
+    -0.006917668027039294
+      0.09194367231922046
+   -9.716765175056498e-05
+   -3.473080935258513e-05
+     -0.01622802243202356
+      0.09152405847322248
+ 1.12e+10    
+       0.0925140825325423
+     -0.01634468101503398
+      0.09276696415458724
+   -3.597593459819988e-05
+    -0.006985291642708011
+      0.09275055827016328
+   -0.0001044658267540569
+   -3.846722088346683e-05
+     -0.01636453908663621
+       0.0923325712536134
+ 1.13e+10    
+      0.09332313933552726
+     -0.01648124939032047
+      0.09357475467495818
+   -3.971213109773956e-05
+    -0.007052259898345823
+      0.09355650299167081
+   -0.0001118968603523486
+   -4.235100295893425e-05
+     -0.01650105244564599
+      0.09314047253191043
+ 1.14e+10    
+      0.09413158095605376
+     -0.01661775558109191
+      0.09438129574987687
+   -4.361134262386075e-05
+     -0.00711859608888459
+      0.09436152185280482
+   -0.0001194636859868413
+   -4.638464242735264e-05
+     -0.01663756041286831
+      0.09394774110400252
+ 1.15e+10    
+      0.09493938780583816
+     -0.01675420185078275
+      0.09518662455475679
+   -4.767534948993358e-05
+    -0.007184322850439458
+      0.09516563020239811
+   -0.0001271691468543749
+   -5.057058312003164e-05
+     -0.01677406102390307
+      0.09475435725650974
+ 1.16e+10    
+        0.095746541678328
+     -0.01689059035243737
+      0.09599077703620072
+   -5.190591993933682e-05
+    -0.007249462178676808
+      0.09596884333494964
+   -0.0001350159939061688
+    -5.49112228608057e-05
+     -0.01691055244033802
+      0.09556030270231293
+ 1.17e+10    
+      0.09655302568903512
+     -0.01702692313485601
+      0.09679378793822488
+   -5.630480572751191e-05
+    -0.007314035446643008
+      0.09677117645974019
+   -0.0001430068840153256
+   -5.940891073529615e-05
+     -0.01704703294427736
+      0.09636556051802829
+ 1.18e+10    
+       0.0973588242176687
+      -0.0171632021485275
+      0.09759569082892074
+   -6.087373802548884e-05
+    -0.007378063422072929
+      0.09757264467293246
+   -0.0001511443783107297
+    -6.40659446057134e-05
+     -0.01718350093316957
+       0.0971701150834067
+ 1.19e+10    
+      0.09816392285204502
+     -0.01729942925134241
+      0.09839651812742853
+   -6.561442362942264e-05
+    -0.007441566284196315
+      0.09837326293243516
+   -0.0001594309406742172
+   -6.888456885762763e-05
+     -0.01731995491491146
+       0.0979739520226325
+ 1.2e+10     
+      0.09896830833375389
+     -0.01743560621408423
+      0.09919630113110406
+    -7.05285414605468e-05
+    -0.007504563640058938
+      0.09917304603532186
+   -0.0001678689363977474
+   -7.386697236610009e-05
+     -0.01745639350320616
+      0.09877705814749599
+ 1.21e+10    
+      0.09977196850555484
+     -0.01757173472569586
+      0.09999507004278171
+   -7.561773934189472e-05
+    -0.007567074540374497
+       0.0999720085976171
+   -0.0001764606309963505
+   -7.901528667121713e-05
+     -0.01759281541315658
+      0.09957942140240954
+ 1.22e+10    
+       0.1005748922604767
+      -0.0177078163983212
+       0.1007928539980386
+   -8.088363103917623e-05
+    -0.007629117494922978
+       0.1007701650362671
+   -0.0001852081891732141
+   -8.433158434985669e-05
+     -0.01772921945707569
+       0.1003810308112388
+ 1.23e+10    
+       0.1013770694925932
+     -0.01784385277212413
+       0.1015896810923852
+   -8.632779354794315e-05
+    -0.007690710487511326
+       0.1015675295531309
+   -0.0001941136739337167
+   -8.981787757348508e-05
+     -0.01786560454049863
+       0.1011818764259167
+ 1.24e+10    
+       0.1021784910494454
+     -0.01797984531988565
+       0.1023855784083101
+   -9.195176462178207e-05
+    -0.007751870990508991
+       0.1023641161208369
+   -0.0002031790458421607
+   -9.547611684396131e-05
+     -0.01800196965838101
+        0.101981949276806
+ 1.25e+10    
+       0.1029791486860778
+     -0.01811579545138379
+       0.1031805720421203
+    -9.77570405217373e-05
+    -0.007812615978973722
+       0.1031599384703594
+   -0.0002124061624190709
+   -0.0001013081898954367
+     -0.01813831389147089
+       0.1027812413247771
+ 1.26e+10    
+       0.1037790350206597
+     -0.01825170451755939
+       0.1039746871305202
+   -0.0001037450739833116
+    -0.007872961944379522
+       0.1039550100801824
+   -0.0002217967776725538
+   -0.0001073159207545978
+     -0.01827463640284244
+       0.1035797454149661
+ 1.27e+10    
+       0.1045781434916561
+      -0.0183875738144731
+       0.1047679478768887
+   -0.0001099172723819837
+    -0.007932924907960557
+       0.1047493441669272
+   -0.0002313525417609289
+   -0.0001135010689505174
+     -0.01841093643458006
+       0.1043774552321749
+ 1.28e+10    
+       0.1053764683165167
+     -0.01852340458705903
+       0.1055603775772109
+   -0.0001162749960941698
+     -0.00799252043368206
+       0.1055429536773246
+   -0.0002410750007803917
+   -0.0001198653288659963
+     -0.01854721330460327
+       0.1051743652578795
+ 1.29e+10    
+       0.1061740044518487
+     -0.01865919803268007
+       0.1063519986456318
+   -0.0001228195570386959
+    -0.008051763640850569
+       0.1063358512814278
+   -0.0002509655966743988
+   -0.0001264103292213476
+     -0.01868346640362361
+       0.1059704707288056
+ 1.3e+10     
+       0.1069707475550361
+     -0.01879495530449191
+       0.1071428326396036
+   -0.0001295522173907068
+    -0.008110669216374588
+       0.1071280493669642
+   -0.0002610256672590282
+   -0.0001331376326858084
+     -0.01881969519222513
+       0.1067657675970374
+ 1.31e+10    
+        0.107766693947277
+     -0.01893067751462213
+       0.1079329002846038
+   -0.0001364741884601434
+    -0.008169251426686194
+       0.1079195600347336
+   -0.0002712564463600931
+   -0.0001400487356071692
+     -0.01895589919806144
+       0.1075602524916172
+ 1.32e+10    
+       0.1085618405779956
+     -0.01906636573717004
+       0.1087222214984012
+   -0.0001435866297233887
+     -0.00822752412933433
+        0.108710395094967
+   -0.0002816590640575289
+   -0.0001471450678531177
+     -0.01909207801316241
+       0.1083539226816031
+ 1.33e+10    
+       0.1093561849905995
+      -0.0192020210110352
+       0.1095108154148574
+   -0.0001508906480017115
+    -0.008285500784259438
+       0.1095005660645657
+   -0.0002922345470317638
+   -0.0001544279927598122
+     -0.01922823129134415
+       0.1091467760405393
+ 1.34e+10    
+       0.1101497252895464
+     -0.01933764434258111
+        0.110298700407249
+   -0.0001583872967779287
+    -0.008343194464759531
+       0.1102900841651466
+   -0.0003029838190081479
+   -0.0001618988071775285
+     -0.01936435874571767
+       0.1099388110123079
+ 1.35e+10    
+       0.1109424601086815
+     -0.01947323670814014
+          0.1110858941111
+   -0.0001660775756431601
+    -0.008400617868156197
+       0.1110789603218253
+   -0.0003139077012941399
+   -0.0001695587416125459
+     -0.01950046014629034
+       0.1107300265783195
+ 1.36e+10    
+       0.1117343885808127
+     -0.01960879905636782
+       0.1118724134465194
+   -0.0001739624298658702
+    -0.008457783326170466
+       0.1118672051626726
+   -0.0003250069134056155
+   -0.0001774089604547353
+     -0.01963653531765568
+       0.1115204222260046
+ 1.37e+10    
+       0.1125255103084904
+     -0.01974433231045257
+       0.1126582746400377
+   -0.0001820427500783156
+    -0.008514702815016102
+       0.1126548290187848
+   -0.0003362820737767202
+   -0.0001854505622892605
+     -0.01977258413676752
+       0.1123099979185712
+ 1.38e+10    
+       0.1133158253359525
+     -0.01987983737018746
+       0.1134434932459395
+    -0.000190319372070502
+     -0.00857138796521967
+       0.1134418419249149
+   -0.0003477337005500835
+   -0.0001936845802836791
+     -0.01990860653079487
+       0.1130987540659874
+ 1.39e+10    
+       0.1141053341222048
+     -0.02001531511391094
+       0.1142280841670929
+   -0.0001987930766875055
+    -0.008627850071174458
+       0.1142282536206114
+    -0.000359362212442088
+   -0.0002021119826496366
+     -0.02004460247505331
+       0.1138866914971555
+ 1.4e+10     
+       0.1148940375151994
+     -0.02015076640032307
+        0.115012061675273
+   -0.0002074645898229798
+    -0.008684100100436569
+        0.115014073551819
+   -0.0003711679296796414
+   -0.0002107336731697563
+     -0.02018057199101037
+       0.1146738114332366
+ 1.41e+10    
+       0.1156819367270789
+     -0.02028619207018322
+       0.1157954394309853
+   -0.0002163345825029083
+    -0.008740148702770742
+       0.1157993108728979
+    -0.000383151075004085
+   -0.0002195504917886096
+      -0.0203165151443616
+       0.1154601154620958
+ 1.42e+10    
+       0.1164690333104523
+      -0.0204215929478954
+       0.1165782305027911
+   -0.0002254036710538638
+    -0.008796006218952381
+       0.1165839744490196
+   -0.0003953117747381436
+   -0.0002285632152622631
+     -0.02045243204317437
+       0.1162456055138253
+ 1.43e+10    
+       0.1172553291356725
+     -0.02055696984298778
+       0.1173604473861366
+   -0.0002346724173510873
+    -0.008851682689333741
+       0.1173680728589041
+   -0.0004076500599121922
+   -0.0002377725578612188
+     -0.02058832283609773
+       0.1170302838373171
+ 1.44e+10    
+       0.1180408263690783
+     -0.02069232355149143
+       0.1181421020216955
+   -0.0002441413291395452
+    -0.008907187862180019
+       0.1181516143978609
+   -0.0004201658674457495
+   -0.0002471791721250704
+     -0.02072418771063428
+        0.117814152977845
+ 1.45e+10    
+       0.1188255274521732
+     -0.02082765485722391
+       0.1189232058132279
+   -0.0002538108604249057
+    -0.008962531201782841
+       0.1189346070811069
+   -0.0004328590413808552
+   -0.0002567836496621539
+     -0.02086002689147417
+       0.1185972157556279
+ 1.46e+10    
+       0.1196094350817097
+       -0.020962964532984
+       0.1197037696449628
+   -0.0002636814119276705
+    -0.009017721896356556
+       0.1197170586473241
+   -0.0004457293341634566
+   -0.0002665865219924372
+      -0.0209958406388868
+       0.1193794752453355
+ 1.47e+10    
+       0.1203925521906458
+      -0.0210982533416615
+       0.1204838038985138
+   -0.0002737533315974683
+    -0.009072768865723967
+       0.1204989765624381
+   -0.0004587764079691681
+   -0.0002765882614306509
+     -0.02113162924717015
+       0.1201609347565095
+ 1.48e+10    
+       0.1211748819299467
+     -0.02123352203726759
+       0.1212633184693315
+   -0.0002840269151832628
+    -0.009127680768797008
+       0.1212803680235845
+    -0.000471999836070392
+   -0.0002867892820031534
+     -0.02126739304315473
+       0.1209415978148645
+ 1.49e+10    
+        0.121956427651202
+      -0.0213687713658912
+       0.1220423227827065
+   -0.0002945024068515162
+    -0.009182466010858877
+       0.1220612399632462
+   -0.0004853991042416332
+   -0.0002971899403992175
+     -0.02140313238476115
+         0.12172146814444
+ 1.5e+10     
+       0.1227371928900283
+     -0.02150400206658442
+       0.1228208258093245
+    -0.000305179999855903
+    -0.009237132750651349
+       0.1228415990535352
+   -0.0004989736121986613
+   -0.0003077905369512201
+     -0.02153884765960895
+        0.122500549650571
+ 1.51e+10    
+       0.1235171813502309
+     -0.02163921487218269
+       0.1235988360803905
+   -0.0003160598372460977
+    -0.009291688907275025
+       0.1236214517106031
+    -0.000512722675070288
+   -0.0003185913166410363
+     -0.02167453928367622
+       0.1232788464036519
+ 1.52e+10    
+       0.1242963968886966
+     -0.02177441051006321
+       0.1243763617023235
+   -0.0003271420126176752
+     -0.00934614216690555
+       0.1244008040991578
+   -0.0005266455248983852
+    -0.000329592470130622
+     -0.02181020770000738
+       0.1240563626236587
+ 1.53e+10    
+        0.125074843500992
+     -0.02190958970284546
+       0.1251534103710349
+   -0.0003384265708990192
+    -0.009400499989331609
+       0.1251796621370731
+   -0.0005407413121635068
+   -0.0003407941348139223
+     -0.02194585337746817
+       0.1248331026654076
+ 1.54e+10    
+         0.12585252530764
+     -0.02204475316903805
+       0.1259299893858002
+   -0.0003499135091683374
+    -0.009454769614320497
+       0.1259580315000742
+   -0.0005550091073344781
+   -0.0003521963958855612
+     -0.02208147680954705
+       0.1256090710045185
+ 1.55e+10    
+       0.1266294465410508
+     -0.02217990162363518
+       0.1267061056627316
+   -0.0003616027775028184
+    -0.009508958067813758
+       0.1267359176264849
+   -0.0005694479024373664
+   -0.0003637992874282415
+     -0.02221707851320065
+       0.1263842722240594
+ 1.56e+10    
+       0.1274056115330811
+     -0.02231503577866563
+       0.1274817657478599
+   -0.0003734942798519685
+    -0.009563072167959612
+       0.1275133257220221
+   -0.0005840566126433353
+   -0.0003756027935116124
+     -0.02235265902774268
+       0.1271587110018436
+ 1.57e+10    
+       0.1281810247032011
+     -0.02245015634369844
+       0.1282569758298386
+   -0.0003855878749366865
+     -0.00961711853098525
+       0.1282902607646288
+   -0.0005988340778714722
+     -0.00038760684930279
+     -0.02248821891377521
+       0.1279323920983571
+ 1.58e+10    
+       0.1289556905472415
+     -0.02258526402630752
+       0.1290317417522761
+   -0.0003978833771672202
+    -0.009671103576913651
+       0.1290667275093305
+   -0.0006137790644049224
+   -0.0003998113421880348
+     -0.02262375875216005
+       0.1287053203452896
+ 1.59e+10    
+        0.129729613626702
+      -0.0227203595324982
+       0.1298060690257063
+   -0.0004103805575803865
+    -0.009725033535129301
+        0.129842730493108
+   -0.0006288902665182263
+   -0.0004122161128991171
+     -0.02275927914303084
+       0.1294775006346477
+ 1.6e+10     
+        0.130502798558598
+     -0.02285544356709859
+       0.1305799628392073
+   -0.0004230791447929084
+    -0.009778914449796233
+       0.1306182740397761
+   -0.0006441663081129916
+   -0.0004248209566471662
+     -0.02289478070484317
+       0.1302489379084248
+ 1.61e+10    
+       0.1312752500058235
+      -0.0229905168341184
+       0.1313534280716769
+   -0.0004359788259667794
+    -0.009832752185133069
+       0.1313933622648584
+   -0.0006596057443608591
+    -0.000437625624258974
+      -0.0230302640734622
+       0.1310196371488086
+ 1.62e+10    
+       0.1320469726680117
+     -0.02312558003707689
+       0.1321264693027719
+   -0.0004490792477871562
+    -0.009886552430547878
+       0.1321679990804527
+   -0.0006752070633510325
+   -0.0004506298233152633
+     -0.02316572990128683
+       0.1317896033689016
+ 1.63e+10    
+        0.132817971272872
+     -0.02326063387930329
+       0.1328990908235248
+   -0.0004623800174484071
+    -0.009940320705637443
+       0.1329421882000791
+   -0.0006909686877407035
+   -0.0004638332192900196
+     -0.02330117885640925
+       0.1325588416039355
+ 1.64e+10    
+       0.1335882505679848
+     -0.02339567906421065
+         0.13367129664664
+   -0.0004758807036481907
+     -0.00999406236505398
+       0.1337159331435035
+   -0.0007068889764069728
+   -0.0004772354366869291
+     -0.02343661162180873
+       0.1333273569029602
+ 1.65e+10    
+        0.134357815313035
+     -0.02353071629554585
+       0.1344430905164833
+   -0.0004895808375853046
+      -0.0100477826032427
+       0.1344892372415308
+   -0.0007229662260980312
+   -0.0004908360601745014
+     -0.02357202889457884
+       0.1340951543209859
+ 1.66e+10    
+       0.1351266702724668
+     -0.02366574627761761
+       0.1352144759187707
+   -0.0005034799139619871
+     -0.01010148645905391
+       0.1352621036407638
+   -0.0007391986730824534
+   -0.0005046346357161892
+     -0.02370743138518704
+       0.1348622389115605
+ 1.67e+10    
+       0.1358948202085431
+     -0.02380076971550374
+        0.135985456089965
+    -0.000517577391987732
+     -0.01015517882023253
+       0.1360345353083213
+   -0.0007555844947946398
+   -0.0005186306716955099
+     -0.02384281981676531
+       0.1356286157197636
+ 1.68e+10    
+       0.1366622698747908
+     -0.02393578731523963
+       0.1367560340263875
+   -0.0005318726963826803
+     -0.01020886442778865
+        0.136806535036512
+   -0.0007721218114755523
+   -0.0005328236400339338
+     -0.02397819492443163
+       0.1363942897756022
+ 1.69e+10    
+       0.1374290240098167
+     -0.02407079978398943
+       0.1375262124930547
+   -0.0005463652183801733
+     -0.01026254788025156
+       0.1375781054474602
+   -0.0007888086878067857
+   -0.0005472129773014586
+     -0.02411355745464068
+       0.1371592660877856
+ 1.7e+10     
+       0.1381950873314802
+     -0.02420580783020119
+       0.1382959940322446
+   -0.0005610543167255189
+     -0.01031623363781111
+       0.1383492489976796
+   -0.0008056431345370985
+   -0.0005617980858177796
+     -0.02424890816456331
+       0.1379235496378698
+ 1.71e+10    
+       0.1389604645314044
+     -0.02434081216374754
+       0.1390653809718031
+   -0.0005759393186719472
+     -0.01036992602634816
+       0.1391199679825905
+   -0.0008226231100999649
+   -0.0005765783347439803
+     -0.02438424782149316
+       0.1386871453747499
+ 1.72e+10    
+       0.1397251602698134
+     -0.02447581349605272
+       0.1398343754331949
+   -0.0005910195209705481
+     -0.01042362924135802
+       0.1398902645409821
+   -0.0008397465222208444
+    -0.000591553061163169
+     -0.02451957720228071
+       0.1394500582094884
+ 1.73e+10    
+       0.1404891791706809
+     -0.02461081254020753
+       0.1406029793393094
+   -0.0006062941908521795
+     -0.01047734735176924
+       0.1406601406594115
+   -0.0008570112295139057
+   -0.0006067215711493485
+     -0.02465489709279282
+       0.1402122930104661
+ 1.74e+10    
+       0.1412525258171771
+      -0.0247458100110729
+       0.1413711944220248
+   -0.0006217625670045927
+     -0.01053108430365983
+       0.1414295981765418
+   -0.0008744150430658711
+   -0.0006220831408235332
+     -0.02479020828739738
+       0.1409738545988357
+ 1.75e+10    
+          0.1420152047474
+     -0.02488080662537336
+       0.1421390222295396
+   -0.0006374238605386357
+      -0.0105848439238746
+       0.1421986387874145
+    -0.000891955728007098
+    -0.000637637017397023
+     -0.02492551158847205
+       0.1417347477442714
+ 1.76e+10    
+       0.1427772204503793
+     -0.02501580310178106
+       0.1429064641334777
+   -0.0006532772559447556
+     -0.01063862992354531
+       0.1429672640476572
+    -0.000909631005068821
+   -0.0006533824202003434
+     -0.02506080780593679
+       0.1424949771609978
+ 1.77e+10    
+       0.1435385773623411
+     -0.02515080016099116
+       0.1436735213357739
+   -0.0006693219120410369
+     -0.01069244590151628
+       0.1437354753776218
+   -0.0009274385521250129
+   -0.0006693185416973765
+     -0.02519609775680833
+       0.1432545475040838
+ 1.78e+10    
+       0.1442992798632199
+     -0.02528579852578967
+       0.1444401948753426
+   -0.0006855569629071978
+     -0.01074629534767807
+       0.1445032740664556
+   -0.0009453760057191512
+   -0.0006854445484846469
+     -0.02533138226477705
+       0.1440134633659949
+ 1.79e+10    
+       0.1450593322734096
+      -0.0254207989211142
+       0.1452064856345436
+   -0.0007019815188088654
+     -0.01080018164621139
+       0.1452706612761015
+   -0.0009634409625741622
+   -0.0007017595822745373
+     -0.02546666215980452
+       0.1447717292733872
+ 1.8e+10     
+       0.1458187388507403
+     -0.02555580207410801
+       0.1459723943454398
+   -0.0007185946671071651
+     -0.01085410807874332
+       0.1460376380452271
+   -0.0009816309810857134
+   -0.0007182627608623548
+     -0.02560193827774103
+       0.1455293496841321
+ 1.81e+10    
+       0.1465775037876711
+     -0.02569080871416855
+        0.146737921595864
+   -0.0007353954731566963
+     -0.01090807782741842
+       0.1468042052930836
+   -0.0009999435827974493
+   -0.0007349531790765348
+     -0.02573721145996338
+       0.1462863289845672
+ 1.82e+10    
+       0.1473356312086908
+     -0.02582581957299079
+       0.1475030678352915
+   -0.0007523829811876184
+      -0.0109620939778868
+       0.1475703638232921
+    -0.001018376253858422
+   -0.0007518299097116479
+     -0.02587248255303059
+       0.1470426714869526
+ 1.83e+10    
+        0.148093125167914
+      -0.0259608353846057
+       0.1482678333805303
+   -0.0007695562151748131
+     -0.01101615952221085
+       0.1483361143275566
+    -0.001036926446461278
+   -0.0007688920044444337
+      -0.0260077524083582
+        0.147798381427133
+ 1.84e+10    
+       0.1488499896468655
+      -0.0260958568854141
+       0.1490322184212284
+   -0.0007869141796908357
+     -0.01107027736169316
+       0.1491014573893077
+    -0.001055591580261596
+   -0.0007861384947310734
+     -0.02614302188190989
+       0.1485534629623891
+ 1.85e+10    
+       0.1496062285524438
+     -0.02623088481421729
+       0.1497962230252093
+   -0.0008044558607445346
+     -0.01112445030962724
+       0.1498663934872689
+    -0.001074369043777072
+   -0.0008035683926880411
+     -0.02627829183390529
+       0.1493079201694732
+ 1.86e+10    
+       0.1503618457150537
+     -0.02636591991224328
+       0.1505598471436355
+   -0.0008221802266032442
+     -0.01117868109397336
+       0.1506309229989546
+    -0.001093256195767047
+   -0.0008211806919521201
+     -0.02641356312854457
+       0.1500617570428162
+ 1.87e+10    
+       0.1511168448869035
+      -0.0265009629231709
+       0.1513230906160086
+    -0.000840086228598145
+     -0.01123297235996109
+       0.1513950462040927
+    -0.001112250366591329
+   -0.0008389743685243605
+     -0.02654883663374769
+       0.1508149774929034
+ 1.88e+10    
+       0.1518712297404546
+     -0.02663601459315007
+        0.152085953175008
+   -0.0008581728019143462
+     -0.01128732667262036
+       0.1521587632879777
+    -0.001131348859548122
+   -0.0008569483815940287
+     -0.02668411322090879
+       0.1515675853448041
+ 1.89e+10    
+       0.1526250038670199
+     -0.02677107567082029
+        0.152848434451176
+   -0.0008764388663639552
+     -0.01134174651924298
+        0.152922074344748
+    -0.001150548952190962
+   -0.0008751016743440759
+     -0.02681939376466452
+       0.1523195843368536
+ 1.9e+10     
+       0.1533781707754996
+     -0.02690614690732584
+       0.1536105339774489
+    -0.000894883327141252
+      -0.0113962343117764
+       0.1536849793805945
+     -0.00116984789762441
+   -0.0008934331747373261
+     -0.02695467914267597
+       0.1530709781194759
+ 1.91e+10    
+       0.1541307338912539
+     -0.02704122905633032
+       0.1543722511935448
+   -0.0009135050755621379
+     -0.01145079238915136
+       0.1544474783168978
+    -0.001189242925777951
+   -0.0009119417962840997
+     -0.02708997023542327
+       0.1538217702541415
+ 1.92e+10    
+        0.154882696555097
+     -0.02717632287402733
+       0.1551335854502051
+   -0.0009323029897850699
+     -0.01150542301954466
+       0.1552095709932926
+    -0.001208731244658144
+   -0.0009306264387908495
+     -0.02722526792601301
+       0.1545719642124546
+ 1.93e+10    
+       0.1556340620224171
+     -0.02731142911915141
+       0.1558945360133018
+   -0.0009512759355151961
+     -0.01156012840257969
+       0.1559712571706635
+    -0.001228310041579051
+   -0.0009494859890890502
+     -0.02736057309999665
+       0.1553215633753601
+ 1.94e+10    
+       0.1563848334624055
+      -0.0274465485529859
+       0.1566551020678058
+   -0.0009704227666908509
+     -0.01161491067146515
+       0.1567325365340718
+    -0.001247976484370356
+    -0.000968519321745377
+     -0.02749588664520138
+       0.1560705710324685
+ 1.95e+10    
+       0.1571350139573965
+     -0.02758168193937025
+       0.1574152827216285
+   -0.0009897423261520585
+     -0.01166977189507432
+       0.1574934086956124
+    -0.001267727722563453
+   -0.0009877252997531009
+     -0.02763120945157036
+       0.1568189903814884
+ 1.96e+10    
+       0.1578846065023106
+      -0.0277168300447056
+       0.1581750770093348
+    -0.001009233446292438
+     -0.01172471407996586
+       0.1582538731972019
+    -0.001287560888555065
+    -0.001007102775204108
+      -0.0277665424110141
+       0.1575668245277638
+ 1.97e+10    
+       0.1586336140041933
+      -0.0278519936379592
+       0.1589344838957327
+    -0.001028894949692185
+     -0.01177973917234794
+       0.1590139295133011
+    -0.001307473098748783
+    -0.001026650589942095
+     -0.02790188641727111
+       0.1583140764839091
+ 1.98e+10    
+       0.1593820392818475
+     -0.02798717349066774
+       0.1596935022793435
+    -0.001048725649733874
+     -0.01183484905998721
+       0.1597735770535693
+    -0.001327461454674298
+    -0.001046367576196391
+     -0.02803724236577803
+       0.1590607491695389
+ 1.99e+10    
+       0.1601298850655537
+     -0.02812237037693963
+       0.1604521309957562
+    -0.001068724351201805
+     -0.01189004557406314
+       0.1605328151654547
+    -0.001347523044083734
+    -0.001066252557198342
+     -0.02817261115354851
+       0.1598068454110837
+ 2e+10       
+       0.1608771539968728
+      -0.0282575850734564
+       0.1612103688208695
+    -0.001088889850861427
+     -0.01194533049097082
+       0.1612916431367172
+    -0.001367654942026428
+    -0.001086304347777452
+        -0.02830799367906
+       0.1605523679416899
+ 2.01e+10    
+       0.1616238486285272
+     -0.02839281835947289
+       0.1619682144740229
+    -0.001109220938023891
+     -0.01200070553407121
+        0.162050060197889
+    -0.001387854211900626
+    -0.001106521754940405
+     -0.02844339084214884
+       0.1612973194011996
+ 2.02e+10    
+       0.1623699714243565
+      -0.0285280710168169
+       0.1627256666210223
+    -0.001129716395091232
+     -0.01205617237539261
+       0.1628080655246723
+    -0.001408117906483453
+    -0.001126903578430567
+     -0.02857880354391281
+       0.1620417023362034
+ 2.03e+10    
+       0.1631155247593441
+     -0.02866334382988743
+       0.1634827238770616
+    -0.001150374998085438
+     -0.01211173263728248
+       0.1635656582402737
+     -0.00142844306893835
+    -0.001147448611270302
+     -0.02871423268662055
+       0.1627855192001646
+ 2.04e+10    
+       0.1638605109197082
+     -0.02879863758565305
+       0.1642393848095461
+    -0.001171195517159874
+     -0.01216738789401233
+       0.1643228374176769
+    -0.001448826733800437
+    -0.001168155640285181
+     -0.02884967917362719
+       0.1635287723536081
+ 2.05e+10    
+       0.1646049321030578
+     -0.02893395307364808
+       0.1649956479408142
+    -0.001192176717094144
+     -0.01222313967333613
+       0.1650796020818576
+    -0.001469265927939937
+    -0.001189023446609343
+     -0.02898514390929744
+       0.1642714640643747
+ 2.06e+10    
+       0.1653487904186068
+     -0.02906929108596927
+       0.1657515117507695
+    -0.001213317357771439
+     -0.01227898945800353
+       0.1658359512119357
+    -0.001489757671503656
+    -0.001210050806174938
+     -0.02912062779893319
+       0.1650135965079308
+ 2.07e+10    
+       0.1660920878874441
+     -0.02920465241727112
+       0.1665069746794173
+    -0.001234616194639707
+     -0.01233493868722948
+       0.1665918837432712
+    -0.001510298978834601
+    -0.001231236490182833
+     -0.02925613174870759
+       0.1657551717677367
+ 2.08e+10    
+       0.1668348264428556
+     -0.02934003786476008
+       0.1672620351293135
+    -0.001256071979157067
+     -0.01239098875812033
+       0.1673473985695029
+    -0.001530886859369912
+    -0.001252579265557059
+     -0.02939165666560396
+       0.1664961918356644
+ 2.09e+10    
+       0.1675770079306959
+     -0.02947544822818837
+       0.1680166914679265
+    -0.001277683459218853
+     -0.01244714102705897
+       0.1681024945445286
+     -0.00155151831851753
+    -0.001274077895381867
+     -0.02952720345735929
+       0.1672366586124663
+ 2.1e+10     
+       0.1683186341098092
+     -0.02961088430984705
+       0.1687709420299155
+     -0.00129944937957118
+     -0.01250339681104868
+       0.1688571704844314
+    -0.001572190358511222
+    -0.001295731139322564
+     -0.02966277303241283
+       0.1679765739082895
+ 2.11e+10    
+       0.1690597066524897
+     -0.02974634691455806
+       0.1695247851193265
+    -0.001321368482206586
+     -0.01255975738901787
+       0.1696114251693525
+      -0.0015928999792448
+    -0.001317537754029234
+     -0.02979836629985861
+       0.1687159394432323
+ 2.12e+10    
+       0.1698002271449853
+     -0.02988183684966521
+       0.1702782190117094
+    -0.001343439506745219
+     -0.01261622400308554
+       0.1703652573453082
+    -0.001613644179084996
+    -0.001339496493525556
+     -0.02993398416940163
+       0.1694547568479419
+ 2.13e+10    
+       0.1705401970880418
+     -0.03001735492502466
+       0.1710312419561581
+    -0.001365661190800528
+     -0.01267279785978982
+       0.1711186657259555
+    -0.001634419955663863
+      -0.0013616061095804
+     -0.03006962755131828
+       0.1701930276642506
+ 2.14e+10    
+       0.1712796178974783
+     -0.03015290195299446
+       0.1717838521772755
+    -0.001388032270328693
+     -0.01272948013127929
+       0.1718716489943065
+    -0.001655224306650548
+    -0.001383865352065064
+     -0.03020529735641932
+       0.1709307533458455
+ 2.15e+10    
+       0.1720184909048031
+     -0.03028847874842311
+       0.1725360478770679
+    -0.001410551479964839
+     -0.01278627195646916
+       0.1726242058043928
+    -0.001676054230502693
+    -0.001406272969293817
+     -0.03034099449601699
+       0.1716679352589728
+ 2.16e+10    
+       0.1727568173578551
+     -0.03042408612863707
+       0.1732878272367658
+     -0.00143321755334381
+     -0.01284317444216196
+       0.1733763347828781
+    -0.001696906727197588
+    -0.001428827708351136
+     -0.03047671988189372
+       0.1724045746831727
+ 2.17e+10    
+        0.173494598421478
+     -0.03055972491342743
+        0.174039188418579
+    -0.001456029223405742
+     -0.01290018866413502
+       0.1741280345306258
+    -0.001717778798943742
+     -0.00145152831540242
+     -0.03061247442627476
+       0.1731406728120421
+ 2.18e+10    
+       0.1742318351782227
+     -0.03069539592503585
+       0.1747901295673852
+    -0.001478985222689004
+     -0.01295731566819459
+       0.1748793036242152
+    -0.001738667450872466
+    -0.001474373535991887
+     -0.03074825904180174
+       0.1738762307540243
+ 2.19e+10    
+       0.1749685286290734
+     -0.03083109998813888
+       0.1755406488123518
+    -0.001502084283608258
+       -0.013014556471198
+       0.1756301406174148
+    -0.001759569691710299
+    -0.001497362115324762
+      -0.0308840746415099
+       0.1746112495332239
+ 2.2e+10     
+       0.1757046796941981
+     -0.03096683792983204
+       0.1762907442685006
+    -0.001525325138719441
+      -0.0130719120620443
+       0.1763805440426065
+    -0.001780482534432045
+    -0.001520492798536888
+     -0.03101992213880586
+       0.1753457300902441
+ 2.21e+10    
+       0.1764402892137224
+     -0.03110261057961175
+       0.1770404140382043
+    -0.001548706520970897
+     -0.01312938340263476
+       0.1771305124121689
+    -0.001801402996895099
+    -0.001543764330949942
+     -0.03115580244744808
+       0.1760796732830442
+ 2.22e+10    
+       0.1771753579485238
+     -0.03123841876935781
+       0.1777896562126323
+    -0.001572227163941848
+     -0.01318697142880355
+       0.1778800442198127
+    -0.001822328102455068
+    -0.001567175458313605
+     -0.03129171648152825
+        0.176813079887819
+ 2.23e+10    
+       0.1779098865810427
+     -0.03137426333331279
+       0.1785384688731335
+    -0.001595885802068424
+     -0.01324467705121942
+       0.1786291379418782
+    -0.001843254880562796
+    -0.001590724927035023
+      -0.0314276651554545
+       0.1775459505998936
+ 2.24e+10    
+       0.1786438757161144
+     -0.03151014510806208
+       0.1792868500925671
+    -0.001619681170856295
+     -0.01330250115625949
+        0.179377792038585
+    -0.001864180367343594
+    -0.001614411484394964
+      -0.0315636493839351
+       0.1782782860346349
+ 2.25e+10    
+       0.1793773258818141
+     -0.03164606493251133
+       0.1800347979365777
+    -0.001643612007081693
+     -0.01336044460685563
+       0.1801260049552469
+    -0.001885101606158436
+     -0.00163823387875197
+     -0.03169967008196383
+       0.1790100867283799
+ 2.26e+10    
+       0.1801102375303194
+     -0.03178202364786374
+       0.1807823104648204
+    -0.001667677048981132
+     -0.01341850824331391
+       0.1808737751234429
+    -0.001906015648147394
+    -0.001662190859734765
+     -0.03183572816480593
+       0.1797413531393762
+ 2.27e+10    
+        0.180842611038784
+     -0.03191802209759589
+       0.1815293857321336
+    -0.001691875036427432
+     -0.01347669288410879
+       0.1816211009621503
+    -0.001926919552756225
+    -0.001686281178421933
+     -0.03197182454798436
+       0.1804720856487332
+ 2.28e+10    
+       0.1815744467102255
+     -0.03205406112743166
+       0.1822760217896652
+    -0.001716204711097263
+     -0.01353499932665135
+       0.1823679808788386
+    -0.001947810388245389
+    -0.001710503587510712
+     -0.03210796014726714
+       0.1812022845613891
+ 2.29e+10    
+       0.1823057447744233
+     -0.03219014158531593
+       0.1830222166859478
+    -0.001740664816624603
+     -0.01359342834803351
+       0.1831144132705287
+    -0.001968685232182739
+    -0.001734856841474808
+     -0.03224413587865459
+        0.181931950107082
+ 2.3e+10     
+       0.1830365053888268
+     -0.03232626432138615
+       0.1837679684679315
+    -0.001765254098746334
+     -0.01365198070574807
+       0.1838603965248124
+    -0.001989541171919401
+    -0.001759339696710461
+     -0.03238035265836731
+       0.1826610824413353
+ 2.31e+10    
+       0.1837667286394744
+     -0.03246243018794323
+       0.1845132751819703
+    -0.001789971305434464
+      -0.0137106571383858
+       0.1846059290208382
+    -0.002010375305049795
+    -0.001783950911672596
+     -0.03251661140283352
+       0.1833896816464468
+ 2.32e+10    
+       0.1844964145419171
+     -0.03259864003942053
+       0.1852581348747654
+    -0.001814815187020347
+     -0.01376945836630958
+       0.1853510091302613
+    -0.002031184739855412
+     -0.00180868924700012
+     -0.03265291302867719
+       0.1841177477324863
+ 2.33e+10    
+       0.1852255630421523
+     -0.03273489473235217
+       0.1860025455942674
+    -0.001839784496307766
+      -0.0138283850923071
+       0.1860956352181621
+    -0.002051966595733171
+    -0.001833553465631696
+     -0.03278925845270583
+       0.1848452806383012
+ 2.34e+10    
+       0.1859541740175633
+     -0.03287119512533939
+       0.1867465053905366
+    -0.001864877988676491
+     -0.01388743800222155
+       0.1868398056439266
+    -0.002072718003608358
+    -0.001858542332911146
+      -0.0329256485918973
+       0.1855722802325216
+ 2.35e+10    
+       0.1866822472778635
+     -0.03300754207901582
+       0.1874900123165653
+    -0.001890094422176965
+     -0.01394661776556193
+       0.1875835187620994
+    -0.002093436106332461
+    -0.001883654616683876
+      -0.0330620843633875
+       0.1862987463145764
+ 2.36e+10    
+       0.1874097825660458
+     -0.03314393645601155
+       0.1882330644290612
+    -0.001915432557614749
+     -0.01400592503609338
+       0.1883267729232038
+    -0.002114118059066373
+    -0.001908889087383386
+     -0.03319856668445685
+       0.1870246786157074
+ 2.37e+10    
+       0.1881367795593353
+     -0.03328037912091505
+        0.188975659789194
+    -0.001940891158627303
+     -0.01406536045240716
+        0.189069566474529
+    -0.002134761029648804
+    -0.001934244518109971
+     -0.03333509647251622
+       0.1877500767999892
+ 2.38e+10    
+       0.1888632378701473
+       -0.033416870940235
+       0.1897177964633071
+     -0.00196646899175121
+     -0.01412492463847238
+       0.1898118977608895
+    -0.002155362198950876
+    -0.001959719684699077
+     -0.03347167464509282
+       0.1884749404653501
+ 2.39e+10    
+        0.189589157047045
+     -0.03355341278235931
+       0.1904594725235928
+    -0.001992164826481523
+     -0.01418461820416838
+        0.190553765125355
+    -0.002175918761216323
+    -0.001985313365783399
+     -0.03360830211981465
+       0.1891992691445931
+ 2.4e+10     
+       0.1903145365757012
+     -0.03369000551751366
+       0.1912006860487361
+    -0.002017977435322765
+     -0.01424444174579996
+       0.1912951669099509
+     -0.00219642792438854
+    -0.002011024342844213
+     -0.03374497981439496
+       0.1899230623064208
+ 2.41e+10    
+       0.1910393758798607
+     -0.03382665001771813
+       0.1919414351245247
+    -0.002043905593832321
+     -0.01430439584659426
+        0.192036101456332
+    -0.002216886910423675
+     -0.00203685140025759
+     -0.03388170864661519
+        0.190646319356457
+ 2.42e+10    
+       0.1917636743223032
+     -0.03396334715674263
+       0.1926817178444282
+    -0.002069948080656085
+     -0.01436448107718103
+       0.1927765671064276
+    -0.002237292955591187
+    -0.002062793325330558
+     -0.03401848953430731
+       0.1913690396382692
+ 2.43e+10    
+       0.1924874312058074
+     -0.03410009781006061
+       0.1934215323101457
+    -0.002096103677556342
+     -0.01442469799605657
+       0.1935165622030629
+    -0.002257643310761199
+    -0.002088848908331645
+     -0.03415532339533535
+       0.1920912224343909
+ 2.44e+10    
+       0.1932106457741134
+     -0.03423690285480186
+       0.1941608766321263
+     -0.00212237116943361
+     -0.01448504715003121
+       0.1942560850905519
+    -0.002277935241679432
+    -0.002115016942513146
+      -0.0342922111475756
+       0.1928128669673409
+ 2.45e+10    
+       0.1939333172128858
+     -0.03437376316970327
+       0.1948997489300589
+     -0.00214874934434075
+      -0.0145455290746614
+       0.1949951341152669
+    -0.002298166029229778
+    -0.002141296224127299
+     -0.03442915370889603
+       0.1935339724006425
+ 2.46e+10    
+       0.1946554446506745
+     -0.03451067963505816
+       0.1956381473333353
+    -0.002175236993490173
+     -0.01460614429466677
+       0.1957337076261829
+    -0.002318332969685114
+    -0.002167685552435185
+      -0.0345661519971342
+       0.1942545378398381
+ 2.47e+10    
+       0.1953770271598753
+     -0.03464765313266498
+       0.1963760699814869
+    -0.002201832911255882
+     -0.01466689332433224
+       0.1964718039753991
+    -0.002338433374946019
+    -0.002194183729709646
+     -0.03470320693007445
+       0.1949745623335029
+ 2.48e+10    
+       0.1960980637576862
+     -0.03478468454577326
+       0.1971135150245956
+    -0.002228535895168366
+     -0.01472777666789616
+       0.1972094215186369
+    -0.002358464572768227
+    -0.002220789561231999
+     -0.03484031942542323
+        0.195694044874254
+ 2.49e+10    
+       0.1968185534070642
+     -0.03492177475902916
+       0.1978504806236791
+    -0.002255344745903426
+     -0.01478879481992454
+       0.1979465586157152
+    -0.002378423906978935
+    -0.002247501855282453
+     -0.03497749040078431
+       0.1964129843997573
+ 2.5e+10     
+       0.1975384950176771
+     -0.03505892465841923
+       0.1985869649510521
+    -0.002282258267266371
+     -0.01484994826567151
+       0.1986832136310039
+    -0.002398308737681912
+    -0.002274319423125368
+     -0.03511472077363103
+       0.1971313797937295
+ 2.51e+10    
+        0.198257887446853
+     -0.03519613513121248
+       0.1993229661906666
+    -0.002309275266169484
+     -0.01491123748142746
+        0.199419384933857
+    -0.002418116441452198
+    -0.002301241078988452
+       -0.035252011461279
+       0.1978492298869355
+ 2.52e+10    
+       0.1989767295005269
+     -0.03533340706590146
+       0.2000584825384262
+    -0.002336394552605205
+     -0.01497266293485376
+       0.2001550708990245
+    -0.002437844411520153
+    -0.002328265640037033
+     -0.03538936338085607
+       0.1985665334581832
+ 2.53e+10    
+       0.1996950199341829
+     -0.03547074135214122
+       0.2007935122024803
+    -0.002363614939613305
+     -0.01503422508530596
+        0.200890269907044
+    -0.002457490057945444
+    -0.002355391926343441
+      -0.0355267774492718
+       0.1992832892353114
+ 2.54e+10    
+       0.2004127574537928
+     -0.03560813888068799
+       0.2015280534034987
+    -0.002390935243243864
+     -0.01509592438414463
+       0.2016249803446122
+    -0.002477050807781152
+    -0.002382618760850767
+     -0.03566425458318466
+       0.1999994958961731
+ 2.55e+10    
+       0.2011299407167504
+     -0.03574560054333503
+       0.2022621043749232
+    -0.002418354282516025
+      -0.0151577612750347
+       0.2023592006049408
+    -0.002496524105227933
+    -0.002409944969332771
+     -0.03580179569896909
+       0.2007151520696149
+ 2.56e+10    
+       0.2018465683328014
+     -0.03588312723284826
+       0.2029956633632019
+    -0.002445870879370961
+      -0.0152197361942341
+       0.2030929290880887
+    -0.002515907411779037
+    -0.002437369380349247
+     -0.03593940171267952
+       0.2014302563364488
+ 2.57e+10    
+       0.2025626388649691
+      -0.0360207198428995
+        0.203728728628003
+     -0.00247348385862145
+      -0.0152818495708708
+       0.2038261642012807
+    -0.002535198206356058
+    -0.002464890825196651
+     -0.03607707354001424
+       0.2021448072304196
+ 2.58e+10    
+       0.2032781508304734
+     -0.03615837926799922
+       0.2044612984424119
+    -0.002501192047897489
+     -0.01534410182721036
+       0.2045589043592076
+    -0.002554393985435634
+    -0.002492508137854897
+     -0.03621481209627714
+       0.2028588032391654
+ 2.59e+10    
+       0.2039931027016477
+     -0.03629610640342756
+       0.2051933710931099
+    -0.002528994277587662
+     -0.01540649337891263
+       0.2052911479843081
+    -0.002573492263167504
+    -0.002520220154930421
+     -0.03635261829633818
+       0.2035722428051736
+ 2.6e+10     
+       0.2047074929068471
+     -0.03643390214516325
+       0.2059249448805354
+    -0.002556889380776767
+      -0.0154690246352785
+       0.2060228935070361
+    -0.002592490571484024
+    -0.002548025715595807
+     -0.03649049305459195
+       0.2042851243267281
+ 2.61e+10    
+       0.2054213198313545
+     -0.03657176738981255
+       0.2066560181190299
+    -0.002584876193180355
+     -0.01553169599948807
+       0.2067541393661117
+    -0.002611386460201576
+    -0.002575923661524652
+     -0.03662843728491569
+       0.2049974461588524
+ 2.62e+10    
+       0.2061345818182779
+      -0.0367097030345357
+       0.2073865891369682
+    -0.002612953553075485
+     -0.01559450786882851
+       0.2074848840087564
+    -0.002630177497113643
+    -0.002603912836825074
+     -0.03676645190062451
+       0.2057092066142434
+ 2.63e+10    
+       0.2068472771694446
+      -0.0368477099769725
+       0.2081166562768715
+    -0.002641120301228452
+      -0.0156574606349136
+       0.2082151258909127
+    -0.002648861268076408
+    -0.002631992087968396
+     -0.03690453781442593
+       0.2064204039642019
+ 2.64e+10    
+       0.2075594041462877
+     -0.03698578911516665
+       0.2088462178955094
+     -0.00266937528081938
+     -0.01572055468389483
+       0.2089448634774522
+    -0.002667435377086673
+    -0.002660160263715121
+     -0.03704269593837291
+       0.2071310364395526
+ 2.65e+10    
+       0.2082709609707269
+     -0.03712394134748835
+       0.2095752723639845
+    -0.002697717337364463
+     -0.01578379039666348
+       0.2096740952423654
+    -0.002685897446352114
+    -0.002688416215039284
+     -0.03718092718381501
+       0.2078411022315597
+ 2.66e+10    
+        0.208981945826045
+     -0.03726216757255638
+       0.2103038180678047
+    -0.002726145318634647
+     -0.01584716814904537
+       0.2104028196689418
+    -0.002704245116354961
+     -0.00271675879504807
+     -0.03731923246134801
+       0.2085505994928341
+ 2.67e+10    
+       0.2096923568577534
+     -0.03740046868915785
+       0.2110318534069431
+    -0.002754658074572643
+     -0.01591068831198738
+       0.2111310352499339
+    -0.002722476045908145
+    -0.002745186858900786
+     -0.03745761268076238
+       0.2092595263382327
+ 2.68e+10    
+       0.2104021921744578
+     -0.03753884559616758
+       0.2117593767958855
+    -0.002783254457207075
+     -0.01597435125173651
+       0.2118587404877109
+    -0.002740587912204969
+    -0.002773699263724764
+     -0.03759606875098987
+       0.2099678808457529
+ 2.69e+10    
+       0.2111114498487112
+      -0.0376772991924659
+        0.212486386663663
+    -0.002811933320564404
+     -0.01603815733001171
+       0.2125859338943976
+    -0.002758578410862374
+    -0.002802294868528456
+     -0.03773460158004874
+       0.2106756610574163
+ 2.7e+10     
+       0.2118201279178643
+     -0.03781583037685508
+       0.2132128814538772
+    -0.002840693520579067
+      -0.0161021069041687
+       0.2133126139920035
+     -0.00277644525595758
+    -0.002830972534113395
+     -0.03787321207498741
+       0.2113828649801481
+ 2.71e+10    
+       0.2125282243849076
+     -0.03795444004797491
+       0.2139388596247115
+    -0.002869533915001042
+     -0.01616620032735799
+       0.2140387793125394
+    -0.002794186180058842
+    -0.002859731122983628
+       -0.038011901141827
+        0.212089490586646
+ 2.72e+10    
+       0.2132357372193071
+     -0.03809312910421679
+       0.2146643196489324
+    -0.002898453363302539
+     -0.01623043794867618
+       0.2147644283981222
+    -0.002811798934250024
+    -0.002888569499253743
+     -0.03815066968550155
+       0.2127955358162444
+ 2.73e+10    
+       0.2139426643578326
+     -0.03823189844363634
+       0.2153892600138806
+    -0.002927450726582165
+      -0.0162948201133113
+         0.21548955980107
+    -0.002829281288149591
+    -0.002917486528554756
+     -0.03828951860979738
+       0.2135009985757673
+ 2.74e+10    
+       0.2146490037053809
+     -0.03837074896386623
+       0.2161136792214526
+    -0.002956524867467833
+     -0.01635934716268164
+       0.2162141720839867
+    -0.002846631029924045
+    -0.002946481077938721
+      -0.0384284488172915
+       0.2142058767403785
+ 2.75e+10    
+       0.2153547531357896
+     -0.03850968156202563
+       0.2168375757880715
+    -0.002985674650018364
+     -0.01642401943456884
+       0.2169382638198344
+    -0.002863845966295829
+     -0.00297555201578209
+     -0.03856746120928663
+        0.214910168154418
+ 2.76e+10    
+       0.2160599104926454
+     -0.03864869713463079
+        0.217560948244652
+    -0.003014898939623567
+      -0.0164888372632455
+       0.2176618335919995
+    -0.002880923922546119
+    -0.003004698211687635
+     -0.03870655668574717
+       0.2156138706322354
+ 2.77e+10    
+       0.2167644735900856
+     -0.03878779657750291
+       0.2182837951365516
+    -0.003044196602903241
+     -0.01655380097959712
+       0.2183848799943465
+    -0.002897862742512659
+    -0.003033918536384628
+     -0.03884573614523215
+       0.2163169819590132
+ 2.78e+10    
+       0.2174684402135914
+     -0.03892698078567594
+       0.2190061150235176
+    -0.003073566507605462
+      -0.0166189109112385
+       0.2191074016312633
+    -0.002914660288582455
+    -0.003063211861629346
+     -0.03898500048482734
+       0.2170194998915832
+ 2.79e+10    
+       0.2181718081207745
+     -0.03906625065330267
+       0.2197279064796268
+    -0.003103007522502723
+     -0.01668416738262587
+        0.219829397117699
+    -0.002931314441680269
+    -0.003092577060103123
+     -0.03912435060007557
+        0.217721422159233
+ 2.8e+10     
+       0.2188745750421578
+     -0.03920560707355994
+        0.220449168093212
+     -0.00313251851728922
+     -0.01674957071516308
+       0.2205508650791916
+    -0.002947823101252059
+    -0.003122013005310301
+     -0.03926378738490629
+       0.2184227464645072
+ 2.81e+10    
+       0.2195767386819459
+     -0.03934505093855321
+       0.2211698984667884
+    -0.003162098362475017
+     -0.01681512122730407
+       0.2212718041518881
+    -0.002964184185244483
+    -0.003151518571475709
+     -0.03940331173156317
+       0.2191234704839995
+ 2.82e+10    
+        0.220278296718792
+     -0.03948458313921958
+       0.2218900962169671
+    -0.003191745929281664
+     -0.01688081923464995
+       0.2219922129825571
+     -0.00298039563007997
+    -0.003181092633440796
+     -0.03954292453053066
+       0.2198235918691357
+ 2.83e+10    
+       0.2209792468065553
+     -0.03962420456523028
+       0.2226097599743667
+    -0.003221460089536213
+     -0.01694666505004253
+       0.2227120902285932
+    -0.002996455390627852
+    -0.003210734066559721
+     -0.03968262667045905
+       0.2205231082469508
+ 2.84e+10    
+       0.2216795865750511
+     -0.03976391610489172
+       0.2233288883835148
+    -0.003251239715564474
+     -0.01701265898365291
+        0.223431434558013
+    -0.003012361440171673
+    -0.003240441746594928
+     -0.03982241903808795
+       0.2212220172208562
+ 2.85e+10    
+       0.2223793136307945
+       -0.039903718645046
+       0.2240474801027452
+    -0.003281083680085182
+     -0.01707880134306665
+       0.2241502446494478
+     -0.00302811177037251
+     -0.00327021454961241
+     -0.03996230251816951
+       0.2219203163714002
+ 2.86e+10    
+       0.2230784255577362
+     -0.04004361307097034
+       0.2247655338040901
+      -0.0033109908561026
+     -0.01714509243336475
+       0.2248685191921248
+    -0.003043704391229112
+    -0.003300051351876443
+     -0.04010227799338911
+       0.2226180032570204
+ 2.87e+10    
+       0.2237769199179926
+     -0.04018360026627575
+       0.2254830481731652
+    -0.003340960116799758
+     -0.01721153255720088
+       0.2255862568858447
+    -0.003059137331034244
+    -0.003329951029744538
+     -0.04024234634428511
+       0.2233150754147868
+ 2.88e+10    
+       0.2244747942525649
+     -0.04032368111280458
+       0.2262000219090505
+    -0.003370990335431301
+     -0.01727812201487529
+       0.2263034564409516
+    -0.003074408636327919
+      -0.0033599124595622
+     -0.04038250844916813
+       0.2240115303611385
+ 2.89e+10    
+       0.2251720460820554
+     -0.04046385649052729
+       0.2269164537241665
+    -0.003401080385216163
+     -0.01734486110440535
+        0.227020116578298
+    -0.003089516371847562
+    -0.003389934517557145
+     -0.04052276518403811
+       0.2247073655926119
+ 2.9e+10     
+       0.2258686729073725
+     -0.04060412727743851
+       0.2276323423441452
+    -0.003431229139231025
+     -0.01741175012159225
+        0.227736236029203
+    -0.003104458620474772
+    -0.003420016079735034
+     -0.04066311742250046
+       0.2254025785865598
+ 2.91e+10    
+       0.2265646722104319
+     -0.04074449434945231
+       0.2283476865076956
+    -0.003461435470302955
+      -0.0174787893600852
+       0.2284518135354043
+    -0.003119233483179753
+    -0.003450156021773457
+     -0.04080356603568146
+       0.2260971668018653
+ 2.92e+10    
+       0.2272600414548466
+     -0.04088495858029596
+       0.2290624849664677
+    -0.003491698250903314
+     -0.01754597911144246
+       0.2291668478490083
+    -0.003133839078962434
+    -0.003480353218917702
+     -0.04094411189214207
+        0.226791127679643
+ 2.93e+10    
+       0.2279547780866137
+     -0.04102552084140455
+       0.2297767364849109
+    -0.003522016353040633
+     -0.01761331966518938
+       0.2298813377324296
+    -0.003148273544791537
+    -0.003510606545875983
+     -0.04108475585779044
+       0.2274844586439388
+ 2.94e+10    
+       0.2286488795347906
+     -0.04116618200181287
+       0.2304904398401272
+    -0.003552388648155571
+     -0.01768081130887354
+       0.2305952819583295
+    -0.003162535035540493
+    -0.003540914876715552
+     -0.04122549879579376
+       0.2281771571024149
+ 2.95e+10    
+       0.2293423432121661
+     -0.04130694292804772
+        0.231203593821724
+    -0.003582814007015057
+     -0.01774845432811769
+       0.2313086793095497
+     -0.00317662172392156
+     -0.00357127708475871
+     -0.04136634156648887
+       0.2288692204470315
+ 2.96e+10    
+       0.2300351665159215
+     -0.04144780448401987
+       0.2319161972316621
+    -0.003613291299606703
+     -0.01781624900667012
+       0.2320215285790383
+    -0.003190531800417389
+    -0.003601692042480023
+     -0.04150728502729152
+       0.2295606460547205
+ 2.97e+10    
+       0.2307273468282885
+     -0.04158876753091392
+       0.2326282488840989
+    -0.003643819395035385
+     -0.01788419562645192
+       0.2327338285697753
+    -0.003204263473210469
+    -0.003632158621403248
+     -0.04164833003260472
+       0.2302514312880471
+ 2.98e+10    
+        0.231418881517195
+      -0.0417298329270786
+       0.2333397476052321
+    -0.003674397161418922
+     -0.01795229446760306
+       0.2334455780946921
+    -0.003217814968110535
+    -0.003662675691999875
+     -0.04178947743372648
+        0.230941573495869
+ 2.99e+10    
+       0.2321097679369078
+     -0.04187100152791643
+       0.2340506922331373
+    -0.003705023465784531
+     -0.01802054580852548
+       0.2341567759765847
+    -0.003231184528480274
+    -0.003693242123587445
+      -0.0419307280787555
+       0.2316310700139841
+ 3e+10       
+       0.2328000034286648
+     -0.04201227418577188
+       0.2347610816176061
+    -0.003735697173967796
+     -0.01808894992592445
+       0.2348674210480295
+    -0.003244370415158716
+    -0.003723856784229198
+     -0.04207208281249732
+       0.2323199181657717
+ 3.01e+10    
+       0.2334895853213036
+     -0.04215365174982012
+       0.2354709146199793
+    -0.003766417150509667
+     -0.01815750709484773
+       0.2355775121512878
+    -0.003257370906383561
+     -0.00375451854063447
+     -0.04221354247636802
+       0.2330081152628259
+ 3.02e+10    
+       0.2341785109318782
+     -0.04229513506595401
+        0.236180190112979
+    -0.003797182258556627
+      -0.0182262175887233
+       0.2362870481382126
+    -0.003270184297711487
+    -0.003785226258059335
+     -0.04235510790829811
+       0.2336956586055809
+ 3.03e+10    
+       0.2348667775662722
+     -0.04243672497667119
+        0.236888906980539
+    -0.003827991359760753
+     -0.01829508167939466
+       0.2369960278701494
+    -0.003282808901936916
+    -0.003815978800209386
+     -0.04249677994263479
+       0.2343825454839291
+ 3.04e+10    
+       0.2355543825198027
+      -0.0425784223209606
+       0.2375970641176324
+    -0.003858843314180492
+     -0.01836409963715514
+       0.2377044502178342
+    -0.003295243049009767
+    -0.003846775029141925
+     -0.04263855941004383
+       0.2350687731778304
+ 3.05e+10    
+       0.2362413230778196
+     -0.04272022793418825
+       0.2383046604300981
+    -0.003889736980183732
+     -0.01843327173077991
+       0.2384123140612896
+    -0.003307485085951384
+    -0.003877613805170668
+     -0.04278044713740997
+        0.235754338957915
+ 3.06e+10    
+       0.2369275965162941
+     -0.04286214264798262
+       0.2390116948344659
+    -0.003920671214349931
+     -0.01850259822755721
+       0.2391196182897158
+     -0.00331953337676986
+    -0.003908493986769885
+     -0.04292244394773698
+       0.2364392400860782
+ 3.07e+10    
+       0.2376132001024016
+     -0.04300416729011954
+         0.23971816625778
+    -0.003951644871375088
+     -0.01857207939331734
+       0.2398263618013812
+    -0.003331386302373527
+    -0.003939414430481703
+     -0.04306455066004695
+       0.2371234738160676
+ 3.08e+10    
+       0.2382981310951004
+     -0.04314630268440633
+       0.2404240736374192
+    -0.003982656803977249
+     -0.01864171549246101
+       0.2405325435035104
+    -0.003343042260484097
+    -0.003970373990822094
+       -0.043206768089278
+       0.2378070373940615
+ 3.09e+10    
+        0.238982386745697
+     -0.04328854965056612
+         0.24112941592092
+    -0.004013705862802813
+     -0.01871150678798602
+        0.241238162312168
+    -0.003354499665548384
+    -0.004001371520190021
+     -0.04334909704618254
+       0.2384899280592426
+ 3.1e+10     
+       0.2396659642984113
+     -0.04343090900412126
+       0.2418341920657953
+    -0.004044790896334435
+     -0.01878145354151281
+       0.2419432171521408
+    -0.003365756948649415
+    -0.004032405868776808
+     -0.04349153833722309
+         0.23917214304436
+ 3.11e+10    
+       0.2403488609909288
+     -0.04357338155627623
+       0.2425384010393535
+    -0.004075910750800177
+     -0.01885155601330882
+       0.2426477069568183
+    -0.003376812557416602
+    -0.004063475884477316
+     -0.04363409276446882
+       0.2398536795762893
+ 3.12e+10    
+       0.2410310740549498
+     -0.04371596811380064
+       0.2432420418185166
+    -0.004107064270083954
+     -0.01892181446231218
+       0.2433516306680727
+    -0.003387664955935447
+    -0.004094580412801072
+     -0.04377676112549088
+       0.2405345348765783
+ 3.13e+10    
+       0.2417126007167293
+     -0.04385866947891128
+       0.2439451133896367
+    -0.004138250295636843
+     -0.01899222914615352
+       0.2440549872361324
+    -0.003398312624656312
+     -0.00412571829678699
+     -0.04391954421325637
+       0.2412147061619915
+ 3.14e+10    
+        0.242393438197611
+     -0.04400148644915438
+       0.2446476147483147
+    -0.004169467666390525
+     -0.01906280032117789
+       0.2447577756194595
+    -0.003408754060302891
+    -0.004156888376917215
+     -0.04406244281602281
+       0.2418941906450442
+ 3.15e+10    
+       0.2430735837145541
+     -0.04414441981728712
+       0.2453495448992142
+    -0.004200715218671749
+     -0.01913352824246508
+       0.2454599947846205
+    -0.003418987775780098
+    -0.004188089491033454
+     -0.04420545771723104
+       0.2425729855345286
+ 3.16e+10    
+       0.2437530344806523
+     -0.04428747037115907
+       0.2460509028558797
+    -0.004231991786117249
+     -0.01920441316384949
+       0.2461616437061591
+    -0.003429012300081714
+    -0.004219320474254704
+     -0.04434858969539818
+       0.2432510880360354
+ 3.17e+10    
+       0.2444317877056479
+     -0.04443063889359317
+       0.2467516876405501
+    -0.004263296199592227
+     -0.01927545533793878
+       0.2468627213664654
+    -0.003438826178197405
+    -0.004250580158895881
+      -0.0444918395240092
+       0.2439284953524637
+ 3.18e+10    
+       0.2451098405964362
+     -0.04457392616226663
+        0.247451898283977
+    -0.004294627287108336
+     -0.01934665501613273
+       0.2475632267556453
+    -0.003448427971019724
+    -0.004281867374388531
+     -0.04463520797140863
+       0.2446052046845291
+ 3.19e+10    
+       0.2457871903575654
+     -0.04471733294959106
+       0.2481515338252364
+     -0.00432598387374382
+     -0.01941801244864029
+       0.2482631588713868
+     -0.00345781625525097
+    -0.004313180947202323
+     -0.04477869580069158
+       0.2452812132312603
+ 3.2e+10     
+        0.246463834191728
+     -0.04486086002259339
+       0.2488505933115474
+    -0.004357364781565642
+     -0.01948952788449694
+       0.2489625167188265
+    -0.003466989623309635
+      -0.0043445197007687
+     -0.04492230376959368
+       0.2459565181904899
+ 3.21e+10    
+       0.2471397693002474
+     -0.04500450814279552
+       0.2495490757980862
+    -0.004388768829552246
+     -0.01956120157158105
+       0.2496612993104159
+     -0.00347594668323705
+    -0.004375882455405778
+     -0.04506603263038134
+       0.2466311167593372
+ 3.22e+10    
+       0.2478149928835547
+      -0.0451482780660943
+       0.2502469803478015
+    -0.004420194833518746
+     -0.01963303375662983
+       0.2503595056657835
+    -0.003484686058603925
+    -0.004407268028244482
+     -0.04520988312974067
+       0.2473050061346869
+ 3.23e+10    
+       0.2484895021416615
+     -0.04529217054264113
+       0.2509443060312305
+    -0.004451641606043076
+     -0.01970502468525484
+       0.2510571348115994
+    -0.003493206388416928
+    -0.004438675233156794
+     -0.04535385600866672
+       0.2479781835136564
+ 3.24e+10    
+       0.2491632942746247
+     -0.04543618631672168
+       0.2516410519263164
+    -0.004483107956393866
+     -0.01977717460195723
+       0.2517541857814379
+    -0.003501506327025446
+    -0.004470102880685108
+     -0.04549795200235186
+       0.2486506460940591
+ 3.25e+10    
+       0.2498363664830042
+     -0.04558032612663501
+       0.2523372171182222
+    -0.004514592690460537
+     -0.01984948375014211
+        0.252450657615638
+    -0.003509584544028285
+    -0.004501549777973681
+     -0.04564217184007355
+       0.2493223910748589
+ 3.26e+10    
+       0.2505087159683149
+     -0.04572459070457314
+       0.2530328006991509
+    -0.004546094610683596
+     -0.01992195237213319
+        0.253146549361166
+    -0.003517439724181059
+     -0.00453301472870107
+     -0.04578651624508225
+       0.2499934156566196
+ 3.27e+10    
+       0.2511803399334709
+     -0.04586898077650006
+       0.2537278017681611
+     -0.00457761251598823
+     -0.01999458070918685
+       0.2538418600714755
+    -0.003525070567303315
+     -0.00456449653301487
+     -0.04593098593448842
+       0.2506637170419452
+ 3.28e+10    
+       0.2518512355832251
+      -0.0460134970620306
+       0.2544222194309851
+    -0.004609145201718657
+     -0.02006736900150572
+       0.2545365888063662
+    -0.003532475788186358
+    -0.004595993987467335
+     -0.04607558161914958
+       0.2513332924359146
+ 3.29e+10    
+       0.2525214001245989
+     -0.04615814027430987
+       0.2551160527998484
+    -0.004640691459574148
+     -0.02014031748825252
+       0.2552307346318468
+    -0.003539654116501261
+    -0.004627505884953375
+     -0.04622030400355689
+       0.2520021390465092
+ 3.3e+10     
+       0.2531908307673083
+     -0.04630291111989171
+       0.2558093009932889
+    -0.004672250077546897
+     -0.02021342640756314
+       0.2559242966199901
+    -0.003546604296707358
+    -0.004659031014650155
+     -0.04636515378572102
+        0.252670254085033
+ 3.31e+10    
+       0.2538595247241824
+     -0.04644781029861799
+       0.2565019631359769
+    -0.004703819839861805
+     -0.02028669599656005
+       0.2566172738487957
+    -0.003553325087961295
+    -0.004690568161957448
+     -0.04651013165705866
+        0.253337634766527
+ 3.32e+10    
+       0.2545274792115743
+     -0.04659283850349697
+       0.2571940383585358
+    -0.004735399526917448
+     -0.02036012649136526
+        0.257309665402047
+     -0.00355981526402637
+    -0.004722116108441086
+     -0.04665523830227767
+       0.2540042783101764
+ 3.33e+10    
+       0.2551946914497674
+     -0.04673799642058316
+       0.2578855257973653
+    -0.004766987915229459
+     -0.02043371812711327
+       0.2580014703691695
+    -0.003566073613182583
+    -0.004753673631777111
+      -0.0468004743992627
+       0.2546701819397092
+ 3.34e+10    
+       0.2558611586633734
+     -0.04688328472885493
+       0.2585764245944628
+    -0.004798583777374788
+     -0.02050747113796403
+        0.258692687845091
+     -0.00357209893813743
+    -0.004785239505697743
+      -0.0469458406189607
+       0.2553353428837922
+ 3.35e+10    
+       0.2565268780817264
+      -0.0470287041000947
+       0.2592667338972474
+    -0.004830185881938654
+     -0.02058138575711548
+       0.2593833169300999
+    -0.003577890055936883
+    -0.004816812499939758
+     -0.04709133762526538
+       0.2559997583764149
+ 3.36e+10    
+       0.2571918469392663
+      -0.0471742551987668
+       0.2599564528583852
+    -0.004861792993462431
+     -0.02065546221681663
+       0.2600733567297013
+    -0.003583445797877606
+    -0.004848391380193488
+     -0.04723696607490224
+       0.2566634256572725
+ 3.37e+10    
+       0.2578560624759202
+     -0.04731993868189769
+       0.2606455806356144
+    -0.004893403872393729
+     -0.02072970074838005
+       0.2607628063544798
+    -0.003588765009419416
+    -0.004879974908054835
+     -0.04738272661731364
+        0.257326341972138
+ 3.38e+10    
+       0.2585195219374759
+     -0.04746575519895386
+       0.2613341163915723
+    -0.004925017275037974
+      -0.0208041015821947
+       0.2614516649199544
+    -0.003593846550098857
+    -0.004911561840977701
+     -0.04752861989454247
+       0.2579885045732292
+ 3.39e+10    
+       0.2591822225759467
+     -0.04761170539172192
+       0.2620220592936231
+    -0.004956631953512286
+     -0.02087866494773879
+       0.2621399315464411
+     -0.00359868929344327
+    -0.004943150932229273
+     -0.04767464654111733
+       0.2586499107195694
+ 3.4e+10     
+       0.2598441616499353
+     -0.04775778989418827
+       0.2627094085136876
+    -0.004988246655700356
+     -0.02095339107359238
+       0.2628276053589083
+    -0.003603292126885886
+    -0.004974740930846416
+     -0.04782080718393619
+       0.2593105576773409
+ 3.41e+10    
+       0.2605053364249839
+     -0.04790400933241714
+       0.2633961632280727
+    -0.005019860125209601
+     -0.02102828018745063
+       0.2635146854868406
+    -0.003607653951681707
+    -0.005006330581593988
+     -0.04796710244215147
+       0.2599704427202337
+ 3.42e+10    
+       0.2611657441739264
+     -0.04805036432443198
+        0.264082322617303
+    -0.005051471101330085
+     -0.02110333251613622
+       0.2642011710640954
+    -0.003611773682824305
+    -0.005037918624924982
+     -0.04811353292705299
+       0.2606295631297849
+ 3.43e+10    
+       0.2618253821772272
+     -0.04819685548009407
+       0.2647678858659537
+    -0.005083078318994834
+     -0.02117854828561295
+       0.2648870612287631
+    -0.003615650248963462
+    -0.005069503796942447
+     -0.04826009924195297
+       0.2612879161957143
+ 3.44e+10    
+       0.2624842477233185
+     -0.04834348340098341
+       0.2654528521624855
+    -0.005114680508742786
+     -0.02125392772099858
+        0.265572355123031
+    -0.003619282592323815
+    -0.005101084829362917
+     -0.04840680198207002
+       0.2619454992162529
+ 3.45e+10    
+       0.2631423381089287
+     -0.04849024868027803
+       0.2661372206990774
+     -0.00514627639668216
+     -0.02132947104657817
+       0.2662570518930412
+    -0.003622669668624549
+    -0.005132660449481857
+     -0.04855364173441305
+       0.2626023094984634
+ 3.46e+10    
+       0.2637996506394064
+     -0.04863715190263505
+       0.2668209906714651
+    -0.005177864704456997
+     -0.02140517848581743
+       0.2669411506887527
+    -0.003625810446999997
+    -0.005164229380140857
+     -0.04870061907766517
+       0.2632583443585579
+ 3.47e+10    
+       0.2644561826290379
+     -0.04878419364407163
+       0.2675041612787803
+    -0.005209444149214976
+     -0.02148105026137652
+       0.2676246506638059
+    -0.003628703909921181
+    -0.005195790339696601
+     -0.04884773458206866
+       0.2639136011222061
+ 3.48e+10    
+       0.2651119314013571
+     -0.04893137447184485
+       0.2681867317233858
+    -0.005241013443576244
+     -0.02155708659512337
+       0.2683075509753816
+    -0.003631349053118776
+    -0.005227342041991209
+     -0.04899498880930821
+       0.2645680771248377
+ 3.49e+10    
+       0.2657668942894523
+     -0.04907869494433408
+       0.2688687012107208
+    -0.005272571295605364
+     -0.02163328770814792
+       0.2689898507840673
+    -0.003633744885506741
+    -0.005258883196324903
+     -0.04914238231239611
+       0.2652217697119411
+ 3.5e+10     
+       0.2664210686362636
+     -0.04922615561092185
+       0.2695500689491406
+    -0.005304116408784183
+     -0.02170965382077595
+       0.2696715492537196
+    -0.003635890429107242
+    -0.005290412507430307
+     -0.04928991563555585
+       0.2658746762393534
+ 3.51e+10    
+       0.2670744517948772
+     -0.04937375701187559
+       0.2702308341497599
+    -0.005335647481986758
+     -0.02178618515258325
+       0.2703526455513295
+    -0.003637784718976762
+    -0.005321928675448003
+     -0.04943758931410751
+       0.2665267940735447
+ 3.52e+10    
+       0.2677270411288124
+      -0.0495214996782301
+       0.2709109960262999
+    -0.005367163209455886
+     -0.02186288192241042
+       0.2710331388468881
+    -0.003639426803133277
+    -0.005353430395904597
+     -0.04958540387435197
+       0.2671781205918974
+ 3.53e+10    
+       0.2683788340123019
+     -0.04966938413166969
+       0.2715905537949311
+    -0.005398662280781571
+     -0.02193974434837672
+       0.2717130283132501
+    -0.003640815742484604
+    -0.005384916359692059
+     -0.04973335983345537
+       0.2678286531829787
+ 3.54e+10    
+       0.2690298278305687
+     -0.04981741088441138
+       0.2722695066741266
+    -0.005430143380881232
+     -0.02201677264789583
+       0.2723923131260047
+     -0.00364195061075801
+     -0.00541638525304864
+     -0.04988145769933529
+       0.2684783892468068
+ 3.55e+10    
+       0.2696800199800942
+     -0.04996558043908736
+       0.2729478538845059
+    -0.005461605189981634
+     -0.02209396703768993
+       0.2730709924633397
+    -0.003642830494430979
+    -0.005447835757542215
+     -0.05002969797054495
+       0.2691273261951116
+ 3.56e+10    
+       0.2703294078688824
+     -0.05011389328862951
+       0.2736255946486904
+    -0.005493046383602753
+     -0.02217132773380561
+       0.2737490655059111
+    -0.003643454492663197
+    -0.005479266550054741
+     -0.05017808113615888
+       0.2697754614515901
+ 3.57e+10    
+       0.2709779889167178
+     -0.05026234991615233
+       0.2743027281911524
+    -0.005524465632543005
+     -0.02224885495162873
+       0.2744265314367125
+      -0.0036438217172298
+    -0.005510676302768821
+     -0.05032660767565926
+       0.2704227924521544
+ 3.58e+10    
+       0.2716257605554173
+     -0.05041095079483809
+       0.2749792537380724
+    -0.005555861602866813
+     -0.02232654890590043
+       0.2751033894409458
+    -0.003643931292455996
+     -0.00554206368315552
+     -0.05047527805882098
+       0.2710693166451748
+ 3.59e+10    
+       0.2722727202290762
+     -0.05055969638782138
+       0.2756551705171916
+    -0.005587232955893192
+     -0.02240440981073272
+       0.2757796387058893
+    -0.003643782355152766
+    -0.005573427353964683
+      -0.0506240927455983
+       0.2717150314917167
+ 3.6e+10     
+       0.2729188653943104
+     -0.05070858714807435
+       0.2763304777576714
+    -0.005618578348186791
+      -0.0224824378796248
+       0.2764552784207739
+    -0.003643374054554064
+    -0.005604765973216203
+     -0.05077305218601188
+       0.2723599344657732
+ 3.61e+10    
+       0.2735641935204891
+     -0.05085762351829223
+       0.2770051746899511
+    -0.005649896431550261
+     -0.02256063332547901
+       0.2771303077766523
+    -0.003642705552255181
+    -0.005636078194193339
+     -0.05092215682003452
+       0.2730040230544879
+ 3.62e+10    
+       0.2742087020899657
+     -0.05100680593077984
+       0.2776792605456078
+    -0.005681185853018397
+     -0.02263899636061734
+       0.2778047259662736
+    -0.003641776022152522
+    -0.005667362665437888
+     -0.05107140707747941
+       0.2736472947583782
+ 3.63e+10    
+       0.2748523885983005
+      -0.0511561348073382
+       0.2783527345572189
+    -0.005712445254854125
+      -0.0227175271967985
+       0.2784785321839595
+    -0.003640584650384691
+     -0.00569861803074664
+     -0.05122080337788727
+       0.2742897470915465
+ 3.64e+10    
+       0.2754952505544794
+     -0.05130561055915134
+       0.2790255959582253
+    -0.005743673274546069
+     -0.02279622604523426
+       0.2791517256254778
+    -0.003639130635274926
+     -0.00572984292917012
+     -0.05137034613041418
+       0.2749313775818907
+ 3.65e+10    
+       0.2761372854811267
+     -0.05145523358667479
+       0.2796978439827971
+    -0.005774868544808003
+     -0.02287509311660698
+       0.2798243054879202
+    -0.003637413187274888
+     -0.00576103599501228
+     -0.05152003573372001
+       0.2755721837713058
+ 3.66e+10    
+       0.2767784909147116
+     -0.05160500427952308
+       0.2803694778656982
+    -0.005806029693579583
+     -0.02295412862108659
+       0.2804962709695804
+    -0.003635431528909967
+    -0.005792195857832409
+     -0.05166987257585733
+       0.2762121632158823
+ 3.67e+10    
+       0.2774188644057494
+     -0.05175492301635912
+       0.2810404968421567
+     -0.00583715534402943
+     -0.02303333276834851
+       0.2811676212698312
+    -0.003633184894725664
+      -0.0058233211424485
+     -0.05181985703416007
+       0.2768513134860962
+ 3.68e+10    
+       0.2780584035189983
+     -0.05190499016478307
+       0.2817109001477341
+    -0.005868244114559397
+     -0.02311270576759105
+       0.2818383555890059
+    -0.003630672531235724
+    -0.005854410468942351
+      -0.0519699894751341
+       0.2774896321669981
+ 3.69e+10    
+       0.2786971058336498
+     -0.05205520608122297
+       0.2823806870181969
+    -0.005899294618810464
+     -0.02319224782755351
+       0.2825084731282783
+    -0.003627893696871397
+    -0.005885462452666319
+     -0.05212027025434614
+       0.2781271168583911
+ 3.7e+10     
+       0.2793349689435138
+     -0.05220557111082462
+       0.2830498566893879
+    -0.005930305465670857
+     -0.02327195915653407
+       0.2831779730895443
+    -0.003624847661932296
+     -0.00591647570425155
+     -0.05227069971631523
+        0.278763765175008
+ 3.71e+10    
+       0.2799719904571986
+     -0.05235608558734339
+       0.2837184083971031
+    -0.005961275259284877
+     -0.02335183996240843
+       0.2838468546753057
+    -0.003621533708538638
+    -0.005947448829617903
+     -0.05242127819440326
+       0.2793995747466808
+ 3.72e+10    
+       0.2806081679982859
+     -0.05250674983303573
+       0.2843863413769664
+    -0.005992202599064515
+     -0.02343189045264802
+       0.2845151170885538
+    -0.003617951130584789
+    -0.005978380429985695
+     -0.05257200601070723
+       0.2800345432185057
+ 3.73e+10    
+       0.2812434992054988
+      -0.0526575641585517
+       0.2850536548643097
+     -0.00602308607970165
+     -0.02351211083433892
+       0.2851827595326537
+    -0.003614099233694428
+    -0.006009269101888759
+     -0.05272288347595058
+       0.2806686682510004
+ 3.74e+10    
+       0.2818779817328678
+     -0.05280852886282836
+       0.2857203480940492
+    -0.006053924291182667
+     -0.02359250131420045
+       0.2858497812112323
+    -0.003609977335177056
+    -0.006040113437189314
+     -0.05287391088937659
+       0.2813019475202618
+ 3.75e+10    
+       0.2825116132498869
+     -0.05295964423298317
+       0.2863864203005689
+    -0.006084715818803996
+      -0.0236730620986044
+       0.2865161813280644
+    -0.003605584763985981
+    -0.006070912023094292
+     -0.05302508853864125
+       0.2819343787181117
+ 3.76e+10    
+         0.28314439144167
+     -0.05311091054420895
+       0.2870518707176019
+    -0.006115459243189892
+     -0.02375379339359415
+       0.2871819590869615
+    -0.003600920860677754
+    -0.006101663442173184
+     -0.05317641669970725
+       0.2825659595522408
+ 3.77e+10    
+       0.2837763140090969
+     -0.05326232805966882
+       0.2877166985781159
+    -0.006146153140311375
+     -0.02383469540490397
+       0.2878471136916625
+    -0.003595984977373065
+    -0.006132366272377671
+     -0.05332789563673892
+       0.2831966877463489
+ 3.78e+10    
+       0.2844073786689585
+     -0.05341389703039277
+       0.2883809031141985
+    -0.006176796081506749
+     -0.02391576833797872
+       0.2885116443457229
+    -0.003590776477719113
+    -0.006163019087062597
+     -0.05347952560199647
+       0.2838265610402764
+ 3.79e+10    
+       0.2850375831540937
+     -0.05356561769517325
+       0.2890444835569436
+    -0.006207386633504058
+     -0.02399701239799307
+       0.2891755502524079
+    -0.003585294736853481
+    -0.006193620455008538
+     -0.05363130683573265
+       0.2844555771901323
+ 3.8e+10     
+       0.2856669252135217
+     -0.05371749028046391
+       0.2897074391363444
+    -0.006237923358444651
+     -0.02407842778987184
+       0.2898388306145856
+    -0.003579539141369313
+    -0.006224168940446053
+     -0.05378323956608888
+       0.2850837339684191
+ 3.81e+10    
+       0.2862954026125732
+       -0.053869515000277
+       0.2903697690811783
+    -0.006268404813908473
+     -0.02416001471830937
+       0.2905014846346201
+    -0.003573509089282338
+    -0.006254663103081004
+     -0.05393532400899207
+        0.285711029164149
+ 3.82e+10    
+       0.2869230131330092
+     -0.05402169205608259
+       0.2910314726189044
+    -0.006298829552941031
+     -0.02424177338778998
+       0.2911635115142694
+    -0.003567203989998869
+    -0.006285101498121995
+     -0.05408756036805308
+       0.2863374605829577
+ 3.83e+10    
+       0.2875497545731432
+     -0.05417402163670897
+        0.291692548975555
+    -0.006329196124081474
+     -0.02432370400260797
+       0.2918249104545808
+    -0.003560623264285803
+    -0.006315482676308732
+     -0.05423994883446522
+       0.2869630260472134
+ 3.84e+10    
+       0.2881756247479513
+     -0.05432650391824229
+        0.292352997375631
+    -0.006359503071392685
+     -0.02440580676688765
+       0.2924856806557876
+    -0.003553766344241697
+    -0.006345805183942175
+     -0.05439248958690263
+       0.2875877233961169
+ 3.85e+10    
+       0.2888006214891812
+     -0.05447913906392913
+       0.2930128170419997
+    -0.006389748934492222
+     -0.02448808188460416
+       0.2931458213172109
+    -0.003546632673269558
+    -0.006376067562916109
+     -0.05454518279142178
+       0.2882115504858047
+ 3.86e+10    
+       0.2894247426454565
+     -0.05463192722407806
+       0.2936720071957942
+    -0.006419932248585566
+      -0.0245705295596036
+       0.2938053316371589
+    -0.003539221706051004
+    -0.006406268350750057
+      -0.0546980286013614
+       0.2888345051894375
+ 3.87e+10    
+       0.2900479860823743
+     -0.05478486853596332
+       0.2943305670563117
+     -0.00645005154449986
+     -0.02465314999562353
+       0.2944642108128273
+    -0.003531532908522054
+    -0.006436406080623749
+     -0.05485102715724446
+       0.2894565853972932
+ 3.88e+10    
+        0.290670349682599
+     -0.05493796312372847
+        0.294988495840917
+    -0.006480105348719938
+      -0.0247359433963138
+       0.2951224580402029
+    -0.003523565757850242
+    -0.006466479281412809
+     -0.05500417858668026
+       0.2900777890168473
+ 3.89e+10    
+       0.2912918313459518
+     -0.05509121109829226
+       0.2956457927649459
+     -0.00651009218342524
+     -0.02481890996525717
+       0.2957800725139699
+    -0.003515319742413275
+    -0.006496486477726205
+     -0.05515748300426842
+       0.2906981139728541
+ 3.9e+10     
+        0.291912428989493
+     -0.05524461255725303
+       0.2963024570416083
+    -0.006540010566528397
+     -0.02490204990598984
+       0.2964370534274114
+    -0.003506794361779266
+    -0.006526426189944609
+     -0.05531094051150237
+       0.2913175582074201
+ 3.91e+10    
+       0.2925321405476048
+     -0.05539816758479723
+       0.2969584878818976
+    -0.006569859011715194
+      -0.0249853634220225
+       0.2970933999723181
+    -0.003497989126688333
+    -0.006556296934260604
+      -0.0554645511966748
+       0.2919361196800753
+ 3.92e+10    
+       0.2931509639720631
+     -0.05555187625160617
+       0.2976138844944968
+    -0.006599636028485575
+     -0.02506885071686093
+       0.2977491113388953
+    -0.003488903559035751
+    -0.006586097222719869
+     -0.05561831513478272
+       0.2925537963678355
+ 3.93e+10    
+       0.2937688972321089
+     -0.05570573861476498
+        0.298268646085689
+    -0.006629340122196772
+     -0.02515251199402714
+       0.2984041867156739
+    -0.003479537191856571
+    -0.006615825563263945
+      -0.0557722323874359
+       0.2931705862652663
+ 3.94e+10    
+       0.2943859383145137
+     -0.05585975471767216
+       0.2989227718592682
+    -0.006658969794106967
+        -0.02523634745708
+       0.2990586252894173
+    -0.003469889569311683
+    -0.006645480459774304
+     -0.05592630300276275
+       0.2937864873845366
+ 3.95e+10    
+        0.295002085223641
+     -0.05601392458995077
+       0.2995762610164514
+    -0.006688523541420675
+     -0.02532035730963604
+       0.2997124262450354
+    -0.003459960246675465
+    -0.006675060412117548
+     -0.05608052701532006
+       0.2944014977554711
+ 3.96e+10    
+       0.2956173359815016
+     -0.05616824824735949
+       0.3002291127557953
+    -0.006717999857335645
+     -0.02540454175539082
+       0.3003655887654963
+    -0.003449748790324767
+    -0.006704563916192089
+     -0.05623490444600227
+       0.2950156154255968
+ 3.97e+10    
+       0.2962316886278073
+     -0.05632272569170571
+       0.3008813262731095
+    -0.006747397231090637
+     -0.02548890099813923
+       0.3010181120317403
+    -0.003439254777729511
+    -0.006733989463976187
+     -0.05638943530195205
+       0.2956288384601874
+ 3.98e+10    
+       0.2968451412200167
+     -0.05647735691075939
+        0.301532900761375
+    -0.006776714148014746
+     -0.02557343524179682
+       0.3016699952225964
+    -0.003428477797444613
+    -0.006763335543576911
+     -0.05654411957647196
+       0.2962411649422984
+ 3.99e+10    
+       0.2974576918333782
+      -0.0566321418781671
+       0.3021838354106629
+    -0.006805949089578022
+     -0.02565814469042037
+       0.3023212375146965
+    -0.003417417449103476
+    -0.006792600639280838
+     -0.05669895724893667
+       0.2968525929728029
+ 4e+10       
+       0.2980693385609714
+     -0.05678708055336922
+       0.3028341294080551
+    -0.006835100533443137
+     -0.02574302954822888
+       0.3029718380823944
+     -0.00340607334341298
+     -0.00682178323160545
+     -0.05685394828470679
+       0.2974631206704215
+ 4.01e+10    
+       0.2986800795137375
+     -0.05694217288151528
+       0.3034837819375654
+    -0.006864166953518647
+     -0.02582809001962429
+       0.3036217960976869
+     -0.00339444510214978
+    -0.006850881797352127
+     -0.05700909263504381
+        0.298072746171746
+ 4.02e+10    
+       0.2992899128205121
+      -0.0570974187933834
+       0.3041327921800632
+    -0.006893146820013072
+     -0.02591332630921209
+        0.304271110730129
+     -0.00338253235815818
+    -0.006879894809660368
+     -0.05716439023702488
+       0.2986814676312616
+ 4.03e+10    
+       0.2998988366280498
+     -0.05725281820529833
+       0.3047811593131994
+     -0.00692203859949054
+     -0.02599873862182232
+       0.3049197811467607
+     -0.00337033475534947
+    -0.006908820738062755
+     -0.05731984101346055
+       0.2992892832213628
+ 4.04e+10    
+       0.3005068491010457
+     -0.05740837101905246
+       0.3054288825113312
+    -0.006950840754927284
+     -0.02608432716252965
+       0.3055678065120261
+    -0.003357851948702576
+    -0.006937658048541778
+     -0.05747544487281166
+       0.2998961911323664
+ 4.05e+10    
+       0.3011139484221531
+     -0.05756407712182685
+       0.3060759609454494
+    -0.006979551745769749
+     -0.02617009213667434
+       0.3062151859876996
+    -0.003345083604266285
+     -0.00696640520358705
+     -0.05763120170910912
+       0.3005021895725197
+ 4.06e+10    
+       0.3017201327919953
+      -0.0577199363861138
+       0.3067223937831108
+    -0.007008170027993431
+     -0.02625603374988253
+       0.3068619187328103
+    -0.003332029399162838
+    -0.006995060662254391
+      -0.0577871114018734
+       0.3011072767680047
+ 4.07e+10    
+        0.302325400429177
+      -0.0578759486696409
+       0.3073681801883662
+    -0.007036694054163035
+     -0.02634215220808647
+       0.3075080039035679
+    -0.003318689021592955
+    -0.007023622880225445
+     -0.05794317381603574
+       0.3017114509629393
+ 4.08e+10    
+       0.3029297495702846
+     -0.05803211381529525
+        0.308013319321693
+    -0.007065122273493808
+     -0.02642844771754493
+       0.3081534406532923
+    -0.003305062170842286
+    -0.007052090309868624
+     -0.05809938880186107
+       0.3023147104193719
+ 4.09e+10    
+       0.3035331784698916
+     -0.05818843165105037
+       0.3086578103399295
+    -0.007093453131914017
+     -0.02651492048486306
+       0.3087982281323408
+    -0.003291148557289262
+    -0.007080461400301327
+     -0.05825575619487065
+       0.3029170534172742
+ 4.1e+10     
+       0.3041356854005529
+     -0.05834490198989295
+       0.3093016523962103
+    -0.007121685072128302
+     -0.02660157071701268
+       0.3094423654880402
+    -0.003276947902414372
+    -0.007108734597452829
+     -0.05841227581576759
+         0.30351847825453
+ 4.11e+10    
+       0.3047372686527967
+     -0.05850152462975149
+       0.3099448446399015
+    -0.007149816533682261
+     -0.02668839862135185
+       0.3100858518646161
+    -0.003262459938810854
+    -0.007136908344128636
+      -0.0585689474703623
+         0.30411898324692
+ 4.12e+10    
+        0.305337926535115
+     -0.05865829935342647
+       0.3105873862165398
+    -0.007177845953028065
+     -0.02677540440564465
+       0.3107286864031283
+    -0.003247684410196702
+    -0.007164981080075503
+      -0.0587257709494997
+          0.3047185667281
+ 4.13e+10    
+       0.3059376573739464
+     -0.05881522592852076
+       0.3112292762677718
+      -0.0072057717635912
+     -0.02686258827808095
+        0.311370868241404
+    -0.003232621071428139
+    -0.007192951242047775
+     -0.05888274602898818
+       0.3053172270495803
+ 4.14e+10    
+       0.3065364595136587
+     -0.05897230410737266
+       0.3118705139312948
+    -0.007233592395837964
+     -0.02694995044729551
+       0.3120123965139713
+    -0.003217269688514407
+    -0.007220817263874437
+     -0.05903987246952783
+       0.3059149625806954
+ 4.15e+10    
+       0.3071343313165241
+     -0.05912953362698894
+        0.312511098340799
+    -0.007261306277344215
+     -0.02703749112238746
+       0.3126532703519988
+    -0.003201630038634019
+    -0.007248577576527471
+       -0.059197150016643
+       0.3065117717085769
+ 4.16e+10    
+        0.307731271162694
+     -0.05928691420897998
+       0.3131510286259109
+    -0.007288911832865146
+     -0.02712521051293904
+       0.3132934888832316
+    -0.003185701910152181
+     -0.00727623060819085
+     -0.05935457840061348
+        0.307107652838115
+ 4.17e+10    
+       0.3083272774501656
+     -0.05944444555949621
+       0.3137903039121374
+    -0.007316407484405721
+     -0.02721310882903488
+       0.3139330512319315
+    -0.003169485102639776
+    -0.007303774784330638
+     -0.05951215733640857
+       0.3077026043919225
+ 4.18e+10    
+       0.3089223485947497
+     -0.05960212736916522
+       0.3144289233208156
+    -0.007343791651292298
+     -0.02730118628128029
+       0.3145719565188157
+    -0.003152979426893551
+    -0.007331208527766132
+     -0.05966988652362128
+       0.3082966248102916
+ 4.19e+10    
+       0.3095164830300327
+     -0.05975995931303141
+       0.3150668859690571
+     -0.00737106275024517
+     -0.02738944308082004
+       0.3152102038610001
+    -0.003136184704957704
+    -0.007358530258741627
+     -0.05982776564640493
+       0.3088897125511489
+ 4.2e+10     
+       0.3101096792073322
+     -0.05991794105049516
+       0.3157041909696983
+    -0.007398219195451898
+     -0.02747787943935635
+       0.3158477923719425
+    -0.003119100770146737
+    -0.007385738394999274
+     -0.05998579437341105
+       0.3094818660900064
+ 4.21e+10    
+       0.3107019355956535
+     -0.06007607222525581
+       0.3163408374312521
+    -0.007425259398641749
+     -0.02756649556916714
+       0.3164847211613846
+    -0.003101727467069619
+    -0.007412831351852809
+     -0.06014397235772737
+       0.3100730839199072
+ 4.22e+10    
+         0.31129325068164
+     -0.06023435246525369
+       0.3169768244578582
+     -0.00745218176916064
+     -0.02765529168312386
+       0.3171209893352996
+    -0.003084064651655332
+     -0.00743980754226204
+     -0.06030229923681896
+       0.3106633645513704
+ 4.23e+10    
+       0.3118836229695199
+     -0.06039278138261541
+       0.3176121511492375
+    -0.007478984714047376
+     -0.02774426799470867
+       0.3177565959958381
+     -0.00306611219117966
+    -0.007466665376908179
+     -0.06046077463246928
+       0.3112527065123317
+ 4.24e+10    
+       0.3124730509810488
+     -0.06055135857359886
+       0.3182468166006469
+    -0.007505666638110341
+     -0.02783342471803257
+       0.3183915402412744
+    -0.003047869964293147
+    -0.007493403264270143
+     -0.06061939815072372
+       0.3118411083480786
+ 4.25e+10    
+       0.3130615332554537
+     -0.06071008361854154
+       0.3188808199028345
+    -0.007532225944005459
+     -0.02792276206785165
+       0.3190258211659597
+    -0.003029337861050512
+    -0.007520019610701398
+     -0.06077816938183421
+       0.3124285686211857
+ 4.26e+10    
+       0.3136490683493641
+     -0.06086895608180856
+       0.3195141601419977
+    -0.007558661032314271
+     -0.02801228025958452
+       0.3196594378602671
+    -0.003010515782941207
+    -0.007546512820507865
+     -0.06093708790020456
+       0.3130150859114429
+ 4.27e+10    
+       0.3142356548367493
+     -0.06102797551174299
+       0.3201468363997407
+    -0.007584970301623503
+     -0.02810197950932867
+       0.3202923894105482
+    -0.002991403642921249
+    -0.007572881296026231
+     -0.06109615326433902
+       0.3136006588157834
+ 4.28e+10    
+       0.3148212913088468
+     -0.06118714144061863
+       0.3207788477530374
+    -0.007611152148605018
+     -0.02819186003387668
+       0.3209246748990829
+    -0.002972001365446226
+    -0.007599123437703498
+     -0.06125536501679031
+        0.314185285948207
+ 4.29e+10    
+       0.3154059763740893
+     -0.06134645338459176
+       0.3214101932741893
+      -0.0076372049680965
+     -0.02828192205073251
+       0.3215562934040342
+    -0.002952308886505656
+    -0.007625237644176757
+     -0.06141472268411021
+       0.3147689659396992
+ 4.3e+10     
+       0.3159897086580258
+     -0.06150591084365668
+       0.3220408720307896
+    -0.007663127153182986
+     -0.02837216577812689
+       0.3221872439994047
+    -0.002932326153658424
+    -0.007651222312353909
+     -0.06157422577680231
+       0.3153516974381495
+ 4.31e+10    
+       0.3165724868032435
+     -0.06166551330160221
+       0.3226708830856892
+    -0.007688917095279157
+     -0.02846259143503331
+        0.322817525754992
+    -0.002912053126069456
+      -0.0076770758374951
+     -0.06173387378927461
+       0.3159334791082645
+ 4.32e+10    
+       0.3171543094692835
+     -0.06182526022596909
+       0.3233002254969576
+    -0.007714573184212026
+     -0.02855319924118255
+       0.3234471377363461
+    -0.002891489774547615
+    -0.007702796613294814
+     -0.06189366619979488
+       0.3165143096314784
+ 4.33e+10    
+       0.3177351753325542
+     -0.06198515106800932
+       0.3239288983178542
+    -0.007740093808304675
+     -0.02864398941707795
+       0.3240760790047302
+    -0.002870636081584703
+    -0.007728383031964391
+     -0.06205360247044747
+       0.3170941877058612
+ 4.34e+10    
+       0.3183150830862408
+     -0.06214518526264778
+       0.3245569005967934
+    -0.007765477354460282
+     -0.02873496218400982
+       0.3247043486170794
+    -0.002849492041395685
+    -0.007753833484315558
+     -0.06221368204709152
+       0.3176731120460229
+ 4.35e+10    
+       0.3188940314402131
+     -0.06230536222844415
+       0.3251842313773156
+    -0.007790722208247015
+     -0.02882611776406991
+       0.3253319456259638
+    -0.002828057659960003
+    -0.007779146359844214
+      -0.0623739043593204
+       0.3182510813830144
+ 4.36e+10    
+       0.3194720191209284
+     -0.06246568136755706
+       0.3258108896980547
+    -0.007815826753983564
+     -0.02891745638016474
+       0.3259588690795497
+    -0.002806332955064012
+    -0.007804320046815002
+     -0.06253426882042366
+       0.3188280944642266
+ 4.37e+10    
+       0.3200490448713326
+     -0.06262614206571003
+       0.3264368745927128
+    -0.007840789374824911
+     -0.02900897825602986
+       0.3265851180215651
+    -0.002784317956344584
+    -0.007829352932346446
+     -0.06269477482734956
+        0.319404150053286
+ 4.38e+10    
+       0.3206251074507577
+     -0.06278674369215935
+       0.3270621850900335
+    -0.007865608452849157
+     -0.02910068361624253
+       0.3272106914912621
+    -0.002762012705333782
+    -0.007854243402496556
+      -0.0628554217606699
+       0.3199792469299471
+ 4.39e+10    
+       0.3212002056348165
+     -0.06294748559966229
+       0.3276868202137744
+    -0.007890282369144552
+     -0.02919257268623521
+       0.3278355885233885
+    -0.002739417255504578
+    -0.007878989842349114
+     -0.06301620898454703
+       0.3205533838899827
+ 4.4e+10     
+       0.3217743382152952
+     -0.06310836712444817
+       0.3283107789826834
+    -0.007914809503897193
+      -0.0292846456923075
+       0.3284598081481497
+    -0.002716531672317728
+    -0.007903590636100169
+      -0.0631771358467005
+       0.3211265597450686
+ 4.41e+10    
+       0.3223475040000391
+     -0.06326938758619102
+       0.3289340604104749
+    -0.007939188236479164
+      -0.0293769028616389
+       0.3290833493911821
+    -0.002693356033269621
+     -0.00792804416714544
+     -0.06333820167837803
+        0.321698773322671
+ 4.42e+10    
+        0.322919701812842
+     -0.06343054628798311
+       0.3295566635058103
+    -0.007963416945537266
+     -0.02946934442230026
+       0.3297062112735212
+    -0.002669890427941211
+    -0.007952348818167896
+      -0.0634994057943265
+       0.3222700234659257
+ 4.43e+10    
+       0.3234909304933271
+      -0.0635918425163112
+       0.3301785872722752
+    -0.007987494009082177
+     -0.02956197060326561
+       0.3303283928115728
+    -0.002646134958047959
+    -0.007976502971225992
+     -0.06366074749276487
+       0.3228403090335167
+ 4.44e+10    
+       0.3240611888968276
+     -0.06375327554103388
+         0.33079983070836
+    -0.008011417804577998
+      -0.0296547816344231
+       0.3309498930170862
+    -0.002622089737490745
+    -0.008000505007842095
+     -0.06382222605535934
+       0.3234096288995535
+ 4.45e+10    
+       0.3246304758942635
+     -0.06391484461536054
+       0.3314203928074435
+    -0.008035186709032397
+     -0.02974777774658584
+       0.3315707108971282
+    -0.002597754892407901
+    -0.008024353309091558
+     -0.06398384074719971
+       0.3239779819534431
+ 4.46e+10    
+        0.325198790372017
+     -0.06407654897583293
+       0.3320402725577749
+    -0.008058799099086952
+     -0.02984095917150242
+       0.3321908454540582
+    -0.002573130561227971
+    -0.008048046255692195
+     -0.06414559081677793
+       0.3245453670997599
+ 4.47e+10    
+       0.3257661312318032
+     -0.06423838784230718
+       0.3326594689424581
+    -0.008082253351108151
+     -0.02993432614186676
+       0.3328102956855039
+    -0.002548216894723739
+    -0.008071582228093959
+      -0.0643074754959686
+       0.3251117832581171
+ 4.48e+10    
+         0.32633249739054
+      -0.0644003604179387
+       0.3332779809394373
+    -0.008105547841278374
+     -0.03002787889132774
+       0.3334290605843388
+    -0.002523014056066969
+    -0.008094959606569127
+     -0.06446949400001001
+        0.325677229363028
+ 4.49e+10    
+        0.326897887780215
+     -0.06456246588916852
+       0.3338958075214844
+    -0.008128680945687883
+     -0.03012161765449858
+       0.3340471391386604
+     -0.00249752222088409
+    -0.008118176771302764
+      -0.0646316455274888
+       0.3262417043637718
+ 4.5e+10     
+       0.3274623013477465
+     -0.06472470342571122
+        0.334512947656188
+    -0.008151651040426271
+      -0.0302155426669662
+       0.3346645303317732
+    -0.002471741577312903
+    -0.008141232102483595
+     -0.06479392926032512
+       0.3268052072242529
+ 4.51e+10    
+       0.3280257370548492
+     -0.06488707218054507
+       0.3351294003059391
+    -0.008174456501675227
+     -0.03030965416529853
+        0.335281233142165
+    -0.002445672326060047
+    -0.008164123980395083
+     -0.06495634436376017
+       0.3273677369228599
+ 4.52e+10    
+       0.3285881938778893
+     -0.06504957128990348
+        0.335745164427926
+    -0.008197095705800619
+     -0.03040395238705364
+       0.3358972465434927
+    -0.002419314680459475
+    -0.008186850785506895
+     -0.06511888998634562
+       0.3279292924523201
+ 4.53e+10    
+       0.3291496708077422
+     -0.06521219987326869
+        0.336360238974124
+    -0.008219567029445721
+     -0.03049843757078725
+       0.3365125695045654
+    -0.002392668866531589
+    -0.008209410898566536
+     -0.06528156525993428
+        0.328489872819554
+ 4.54e+10    
+       0.3297101668496456
+     -0.06537495703336733
+       0.3369746228912875
+    -0.008241868849624009
+     -0.03059310995605961
+       0.3371272009893279
+    -0.002365735123043387
+    -0.008231802700691265
+     -0.06544436929967387
+       0.3290494770455255
+ 4.55e+10    
+       0.3302696810230503
+     -0.06553784185616762
+       0.3375883151209453
+    -0.008263999543812666
+     -0.03068796978344295
+       0.3377411399568477
+    -0.002338513701569285
+    -0.008254024573460337
+     -0.06560730120400123
+       0.3296081041650907
+ 4.56e+10    
+       0.3308282123614718
+     -0.06570085341087864
+       0.3382013145993968
+    -0.008285957490046181
+     -0.03078301729452753
+       0.3383543853613017
+    -0.002311004866552868
+    -0.008276074899007332
+     -0.06577036005463971
+       0.3301657532268449
+ 4.57e+10    
+       0.3313857599123327
+     -0.06586399074995158
+       0.3388136202577069
+    -0.008307741067009947
+     -0.03087825273192826
+       0.3389669361519657
+    -0.002283208895369271
+    -0.008297952060112681
+     -0.06593354491659781
+        0.330722423292966
+ 4.58e+10    
+       0.3319423227368088
+       -0.066027252909082
+        0.339425231021704
+    -0.008329348654134395
+     -0.03097367633928965
+       0.3395787912732018
+    -0.002255126078388438
+    -0.008319654440296587
+     -0.06609685483816921
+       0.3312781134390572
+ 4.59e+10    
+       0.3324978999096723
+     -0.06619063890721609
+       0.3400361458119802
+    -0.008350778631689091
+     -0.03106928836129183
+       0.3401899496644512
+    -0.002226756719039008
+    -0.008341180423911625
+     -0.06626028885093671
+       0.3318328227539868
+ 4.6e+10     
+       0.3330524905191292
+      -0.0663541477465564
+       0.3406463635438904
+     -0.00837202938087692
+     -0.03116508904365497
+       0.3408004102602259
+    -0.002198101133873001
+    -0.008362528396236179
+     -0.06642384596977596
+       0.3323865503397259
+ 4.61e+10    
+       0.3336060936666571
+     -0.06651777841257107
+       0.3412558831275534
+    -0.008393099283928503
+     -0.03126107863314387
+       0.3414101719901012
+    -0.002169159652631136
+     -0.00838369674356723
+      -0.0665875251928619
+       0.3329392953111822
+ 4.62e+10    
+       0.3341587084668414
+     -0.06668152987400479
+       0.3418647034678564
+    -0.008413986724196888
+     -0.03135725737757196
+       0.3420192337787105
+    -0.002139932618308904
+    -0.008404683853313904
+     -0.06675132550167853
+       0.3334910567960387
+ 4.63e+10    
+       0.3347103340472063
+     -0.06684540108289125
+       0.3424728234644558
+    -0.008434690086251933
+     -0.03145362552580502
+        0.342627594545741
+    -0.002110420387223109
+    -0.008425488114090591
+     -0.06691524586102798
+       0.3340418339345796
+ 4.64e+10    
+       0.3352609695480486
+     -0.06700939097456859
+        0.343080242011785
+    -0.008455207755975167
+     -0.03155018332776438
+       0.3432352532059313
+    -0.002080623329079302
+    -0.008446107915810621
+     -0.06707928521904441
+       0.3345916258795235
+ 4.65e+10    
+       0.3358106141222638
+     -0.06717349846769513
+       0.3436869579990581
+    -0.008475538120654347
+     -0.03164693103442939
+       0.3438422086690669
+    -0.002050541827039606
+    -0.008466541649779509
+     -0.06724344250720789
+         0.33514043179585
+ 4.66e+10    
+        0.336359266935173
+     -0.06733772246426899
+       0.3442929703102786
+     -0.00849567956907844
+     -0.03174386889784035
+        0.344448459839983
+    -0.002020176277791207
+    -0.008486787708788416
+     -0.06740771664036162
+       0.3356882508606253
+ 4.67e+10    
+       0.3369069271643497
+     -0.06750206184964851
+        0.344898277824247
+    -0.008515630491632257
+     -0.03184099717109989
+        0.345054005618562
+    -0.001989527091615404
+    -0.008506844487207883
+     -0.06757210651673046
+       0.3362350822628271
+ 4.68e+10    
+         0.33745359399944
+     -0.06766651549257552
+       0.3455028794145725
+    -0.008535389280391307
+     -0.03193831610837497
+       0.3456588448997374
+    -0.001958594692457229
+    -0.008526710381081149
+     -0.06773661101794194
+       0.3367809252031662
+ 4.69e+10    
+       0.3379992666419853
+     -0.06783108224519974
+         0.34610677394968
+    -0.008554954329216652
+     -0.03203582596489764
+       0.3462629765734946
+    -0.001927379517995513
+     -0.00854638378821756
+     -0.06790122900904898
+       0.3373257788939058
+ 4.7e+10     
+       0.3385439443052402
+     -0.06799576094310635
+       0.3467099602928255
+    -0.008574324033849461
+     -0.03213352699696591
+        0.346866399524876
+    -0.001895882019713561
+    -0.008565863108286199
+     -0.06806595933855525
+       0.3378696425586828
+ 4.71e+10    
+       0.3390876262139894
+     -0.06816055040534442
+       0.3473124373021085
+    -0.008593496792005773
+     -0.03223141946194417
+       0.3474691126339869
+    -0.001864102662970139
+    -0.008585146742909062
+     -0.06823080083844218
+       0.3384125154323221
+ 4.72e+10    
+       0.3396303116043625
+     -0.06832544943445874
+        0.347914203830484
+    -0.008612471003471341
+     -0.03232950361826247
+       0.3480711147760007
+    -0.001832041927071013
+    -0.008604233095754423
+     -0.06839575232419817
+       0.3389543967606526
+ 4.73e+10    
+       0.3401719997236491
+     -0.06849045681652283
+       0.3485152587257825
+     -0.00863124507019576
+     -0.03242777972541688
+       0.3486724048211669
+    -0.001799700305340978
+    -0.008623120572629971
+     -0.06856081259485024
+        0.339495285800321
+ 4.74e+10    
+       0.3407126898301082
+     -0.06865557132117403
+       0.3491156008307211
+    -0.008649817396387103
+     -0.03252624804396734
+       0.3492729816348209
+    -0.001767078305196139
+    -0.008641807581575981
+     -0.06872598043299731
+       0.3400351818186031
+ 4.75e+10    
+       0.3412523811927792
+      -0.0688207917016517
+       0.3497152289829257
+    -0.008668186388606241
+     -0.03262490883553745
+       0.3498728440773936
+    -0.001734176448216608
+    -0.008660292532958131
+     -0.06889125460484674
+       0.3405740840932161
+ 4.76e+10    
+       0.3417910730912889
+     -0.06898611669483629
+       0.3503141420149479
+    -0.008686350455860838
+     -0.03272376236281164
+       0.3504719910044199
+    -0.001700995270219688
+    -0.008678573839560303
+     -0.06905663386025074
+       0.3411119919121227
+ 4.77e+10    
+       0.3423287648156595
+     -0.06915154502129126
+       0.3509123387542853
+    -0.008704308009699501
+     -0.03282280888953366
+       0.3510704212665569
+     -0.00166753532133316
+    -0.008696649916677318
+     -0.06922211693274842
+        0.341648904573345
+ 4.78e+10    
+       0.3428654556661132
+     -0.06931707538530782
+       0.3515098180234039
+    -0.008722057464305434
+     -0.03292204868050365
+       0.3516681337095928
+    -0.001633797166069074
+    -0.008714519182207243
+     -0.06938770253960658
+       0.3421848213847636
+ 4.79e+10    
+       0.3434011449528726
+     -0.06948270647494979
+       0.3521065786397591
+    -0.008739597236590166
+     -0.03302148200157486
+       0.3522651271744625
+    -0.001599781383397669
+    -0.008732180056743815
+     -0.06955338938186495
+       0.3427197416639268
+ 4.8e+10     
+       0.3439358319959666
+     -0.06964843696210327
+        0.352702619415819
+    -0.008756925746286844
+      -0.0331211091196506
+       0.3528614004972659
+    -0.001565488566821664
+     -0.00874963096366815
+     -0.06971917614438287
+       0.3432536647378508
+ 4.81e+10    
+       0.3444695161250267
+     -0.06981426550252635
+       0.3532979391590921
+    -0.008774041416043439
+      -0.0332209303026801
+       0.3534569525092831
+    -0.001530919324450686
+    -0.008766870329240889
+     -0.06988506149588855
+       0.3437865899428232
+ 4.82e+10    
+       0.3450021966790885
+     -0.06998019073590243
+       0.3538925366721487
+    -0.008790942671515692
+     -0.03332094581965424
+       0.3540517820369928
+    -0.001496074279075917
+    -0.008783896582693497
+     -0.07005104408902932
+       0.3443185166241997
+ 4.83e+10    
+       0.3455338730063866
+     -0.07014621128589471
+       0.3544864107526516
+    -0.008807627941459764
+     -0.03342115594060083
+       0.3546458879020932
+    -0.001460954068244938
+     -0.00880070815631962
+     -0.07021712256042681
+       0.3448494441362075
+ 4.84e+10    
+       0.3460645444641517
+     -0.07031232576020409
+       0.3550795601933829
+    -0.008824095657824493
+     -0.03352156093657974
+       0.3552392689215224
+    -0.001425559344336733
+    -0.008817303485566089
+     -0.07038329553073114
+       0.3453793718417396
+ 4.85e+10    
+       0.3465942104184033
+     -0.07047853275062768
+       0.3556719837822727
+    -0.008840344255843702
+     -0.03362216107967707
+        0.355831923907479
+    -0.001389890774636726
+    -0.008833681009123583
+     -0.07054956160467976
+       0.3459082991121518
+ 4.86e+10    
+       0.3471228702437459
+      -0.0706448308331221
+       0.3562636803024311
+    -0.008856372174127679
+     -0.03372295664299953
+       0.3564238516674484
+     -0.00135394904141206
+    -0.008849839169016927
+      -0.0707159193711582
+       0.3464362253270586
+ 4.87e+10    
+       0.3476505233231558
+     -0.07081121856786585
+       0.3568546485321782
+    -0.008872177854754807
+     -0.03382394790066791
+       0.3570150510042241
+    -0.001317734841986744
+    -0.008865776410695338
+     -0.07088236740326176
+       0.3469631498741262
+ 4.88e+10    
+       0.3481771690477752
+     -0.07097769449932656
+       0.3574448872450787
+    -0.008887759743362573
+     -0.03392513512781063
+       0.3576055207159355
+    -0.001281248888817023
+    -0.008881491183121903
+     -0.07104890425836166
+       0.3474890721488669
+ 4.89e+10    
+       0.3487028068166998
+     -0.07114425715632947
+       0.3580343952099739
+     -0.00890311628923833
+     -0.03402651860055651
+       0.3581952595960736
+     -0.00124449190956668
+    -0.008896981938863003
+     -0.07121552847817109
+       0.3480139915544269
+ 4.9e+10     
+       0.3492274360367668
+     -0.07131090505212838
+       0.3586231711910183
+    -0.008918245945409554
+     -0.03412809859602734
+       0.3587842664335189
+    -0.001207464647182259
+    -0.008912247134177331
+     -0.07138223858881584
+        0.348537907501382
+ 4.91e+10    
+       0.3497510561223412
+     -0.07147763668447833
+        0.359211213947715
+    -0.008933147168733882
+     -0.03422987539232995
+        0.359372540012572
+    -0.001170167859968401
+    -0.008927285229104277
+      -0.0715490331009063
+       0.3490608194075231
+ 4.92e+10    
+        0.350273666495101
+      -0.0716444505357117
+       0.3597985222349528
+    -0.008947818419988627
+     -0.03433184926854831
+        0.359960079112983
+    -0.001132602321662915
+    -0.008942094687552238
+     -0.07171591050961126
+       0.3495827266976468
+ 4.93e+10    
+        0.350795266583823
+     -0.07181134507281597
+       0.3603850948030459
+    -0.008962258163959838
+     -0.03443402050473438
+       0.3605468825099827
+    -0.001094768821511919
+    -0.008956673977386295
+     -0.07188286929473488
+       0.3501036288033416
+ 4.94e+10    
+       0.3513158558241635
+     -0.07197831874751386
+       0.3609709303977728
+     -0.00897646486953103
+     -0.03453638938189977
+       0.3611329489743174
+    -0.001056668164344689
+    -0.008971021570515422
+     -0.07204990792079635
+       0.3506235251627757
+ 4.95e+10    
+       0.3518354336584434
+     -0.07214536999634574
+       0.3615560277604165
+     -0.00899043700977142
+     -0.03463895618200565
+       0.3617182772722787
+    -0.001018301170648543
+    -0.008985135942979479
+     -0.07221702483711008
+       0.3511424152204816
+ 4.96e+10    
+       0.3523539995354266
+     -0.07231249724075464
+       0.3621403856278069
+    -0.009004173062023566
+     -0.03474172118795393
+       0.3623028661657463
+   -0.0009796686766433429
+    -0.008999015575035272
+     -0.07238421847787159
+       0.3516602984271412
+ 4.97e+10    
+       0.3528715529101005
+     -0.07247969888717365
+       0.3627240027323656
+    -0.009017671507990736
+     -0.03484468468357637
+       0.3628867144122154
+    -0.000940771534355836
+    -0.009012658951242867
+       -0.072551487262242
+       0.3521771742393706
+ 4.98e+10    
+       0.3533880932434582
+      -0.0726469733271158
+       0.3633068778021469
+    -0.009030930833823688
+     -0.03494784695362459
+       0.3634698207648414
+   -0.0009016106116938725
+    -0.009026064560550544
+     -0.07271882959443773
+       0.3526930421195005
+ 4.99e+10    
+       0.3539036200022719
+     -0.07281431893726532
+       0.3638890095608858
+    -0.009043949530206709
+     -0.03505120828375934
+       0.3640521839724751
+   -0.0008621867925201485
+    -0.009039230896379886
+     -0.07288624386382135
+       0.3532079015353621
+ 5e+10       
+       0.3544181326588736
+     -0.07298173407957294
+       0.3644703967280433
+    -0.009056726092443597
+     -0.03515476896053891
+       0.3646338027797044
+   -0.0008225009767257375
+    -0.009052156456710115
+     -0.07305372844499575
+       0.3537217519600661
+ 5.01e+10    
+       0.3549316306909303
+     -0.07314921710135236
+       0.3650510380188541
+    -0.009069259020542677
+     -0.03525852927140822
+       0.3652146759268939
+   -0.0007825540803033789
+    -0.009064839744161807
+      -0.0732212816978987
+       0.3542345928717828
+ 5.02e+10    
+       0.3554441135812197
+     -0.07331676633537935
+       0.3656309321443754
+    -0.009081546819301435
+     -0.03536248950468663
+       0.3657948021502295
+   -0.0007423470354202078
+    -0.009077279266080132
+     -0.07338890196790357
+       0.3547464237535259
+ 5.03e+10    
+       0.3559555808174055
+     -0.07348438009999426
+       0.3662100778115386
+    -0.009093587998390577
+     -0.03546664994955587
+       0.3663741801817606
+   -0.0007018807904901694
+     -0.00908947353461771
+     -0.07355658758591871
+       0.3552572440929282
+ 5.04e+10    
+       0.3564660318918104
+     -0.07365205669920517
+       0.3667884737231965
+    -0.009105381072437498
+     -0.03557101089604778
+       0.3669528087494455
+   -0.0006611563102460805
+    -0.009101421066816398
+     -0.07372433686849081
+       0.3557670533820204
+ 5.05e+10    
+       0.3569754663011893
+     -0.07381979442279485
+       0.3673661185781797
+    -0.009116924561109168
+     -0.03567557263503107
+       0.3675306865771973
+   -0.0006201745758111145
+    -0.009113120384689149
+     -0.07389214811791209
+       0.3562758511170127
+ 5.06e+10    
+       0.3574838835465028
+     -0.07398759154643009
+        0.367943011071348
+    -0.009128216989194237
+     -0.03578033545819871
+        0.368107812384931
+    -0.000578936584769869
+    -0.009124570015300567
+      -0.0740600196223275
+       0.3567836367980691
+ 5.07e+10    
+       0.3579912831326897
+     -0.07415544633177287
+       0.3685191498936441
+    -0.009139256886684871
+     -0.03588529965805401
+       0.3686841848886127
+   -0.0005374433512388339
+    -0.009135768490847369
+     -0.07422794965584628
+       0.3572904099290849
+ 5.08e+10    
+       0.3584976645684348
+     -0.07432335702659422
+       0.3690945337321511
+    -0.009150042788857535
+      -0.0359904655278971
+       0.3692598028003083
+     -0.00049569590593644
+    -0.009146714348738098
+     -0.07439593647865515
+       0.3577961700174651
+ 5.09e+10    
+       0.3590030273659439
+     -0.07449132186489114
+       0.3696691612701488
+    -0.009160573236353541
+      -0.0360958333618111
+       0.3698346648282352
+   -0.0004536952962523658
+    -0.009157406131671944
+     -0.07456397833713407
+       0.3583009165738986
+ 5.1e+10     
+       0.3595073710407109
+     -0.07465933906700475
+       0.3702430311871695
+    -0.009170846775258529
+     -0.03620140345464724
+       0.3704087696768149
+   -0.0004114425863163094
+    -0.009167842387717114
+      -0.0747320734639756
+       0.3588046491121343
+ 5.11e+10    
+        0.360010695111287
+     -0.07482740683974246
+       0.3708161421590613
+     -0.00918086195718148
+     -0.03630717610201077
+       0.3709821160467242
+   -0.0003689388570661469
+    -0.009178021670388649
+     -0.07490022007830426
+       0.3593073671487563
+ 5.12e+10    
+        0.360512999099052
+     -0.07499552337650137
+       0.3713884928580442
+    -0.009190617339333181
+     -0.03641315160024548
+       0.3715547026349519
+   -0.0003261852063153356
+    -0.009187942538725279
+     -0.07506841638580136
+       0.3598090702029584
+ 5.13e+10    
+       0.3610142825279811
+     -0.07516368685739494
+       0.3719600819527741
+    -0.009200111484603687
+     -0.03651933024641912
+       0.3721265281348544
+   -0.0002831827488196383
+    -0.009197603557365722
+     -0.07523666057883091
+       0.3603097577963199
+ 5.14e+10    
+        0.361514544924412
+      -0.0753318954493816
+       0.3725309081084046
+    -0.009209342961639232
+     -0.03662571233830742
+       0.3726975912362109
+   -0.0002399326163430937
+    -0.009207003296624348
+     -0.07540495083656745
+       0.3608094294525772
+ 5.15e+10    
+        0.362013785816815
+     -0.07550014730639648
+       0.3731009699866504
+    -0.009218310344918492
+     -0.03673229817437841
+       0.3732678906252828
+   -0.0001964359577232078
+    -0.009216140332566056
+     -0.07557328532512787
+       0.3613080846973993
+ 5.16e+10    
+       0.3625120047355578
+     -0.07566844056948527
+       0.3736702662458525
+    -0.009227012214827957
+     -0.03683908805377678
+       0.3738374249848741
+   -0.0001526939389354029
+    -0.009225013247080319
+     -0.07574166219770534
+       0.3618057230581621
+ 5.17e+10    
+       0.3630092012126725
+     -0.07583677336694032
+       0.3742387955410432
+    -0.009235447157736601
+     -0.03694608227630694
+       0.3744061929943899
+   -0.0001087077431565064
+    -0.009233620627954759
+     -0.07591007959470458
+       0.3623023440637186
+ 5.18e+10    
+        0.363505374781624
+      -0.0760051438144403
+       0.3748065565240148
+    -0.009243613766069948
+       -0.037053281142417
+       0.3749741933298991
+   -6.447857082744822e-05
+     -0.00924196106894767
+     -0.07607853564388176
+       0.3627979472441749
+ 5.19e+10    
+       0.3640005249770731
+     -0.07617355001519106
+       0.3753735478433876
+    -0.009251510638382997
+     -0.03716068495318212
+       0.3755414246641977
+   -2.000763971508088e-05
+     -0.00925003316985998
+     -0.07624702846048509
+       0.3632925321306615
+ 5.2e+10     
+       0.3644946513346455
+     -0.07634199006007052
+       0.3759397681446777
+    -0.009259136379432908
+     -0.03726829401028702
+       0.3761078856668732
+    2.470381502706564e-05
+    -0.009257835536606418
+     -0.07641555614739982
+       0.3637860982551073
+ 5.21e+10    
+       0.3649877533906944
+      -0.0765104620277747
+       0.3765052160703697
+     -0.00926648960025038
+     -0.03737610861600897
+       0.3766735750043692
+    6.965454079883859e-05
+    -0.009265366781285856
+     -0.07658411679529382
+       0.3642786451500104
+ 5.22e+10    
+       0.3654798306820673
+     -0.07667896398496653
+       0.3770698902599867
+    -0.009273568918210592
+     -0.03748412907320049
+       0.3772384913400528
+    0.0001148432674946769
+    -0.009272625522250838
+      -0.0767527084827673
+       0.3647701723482116
+ 5.23e+10    
+       0.3659708827458719
+     -0.07684749398642916
+       0.3776337893501646
+    -0.009280372957103091
+     -0.03759235568527138
+       0.3778026333342821
+    0.0001602687074457223
+    -0.009279610384176396
+     -0.07692132927650472
+       0.3652606793826664
+ 5.24e+10    
+       0.3664609091192393
+     -0.07701605007521843
+       0.3781969119747247
+    -0.009286900347201104
+     -0.03770078875617099
+       0.3783659996444745
+    0.0002059295553630664
+    -0.009286319998128009
+     -0.07708997723142864
+       0.3657501657862185
+ 5.25e+10    
+       0.3669499093390902
+     -0.07718463028282101
+       0.3787592567647508
+    -0.009293149725329767
+     -0.03780942859037021
+       0.3789285889251794
+    0.0002518244882821761
+    -0.009292753001628795
+     -0.07725865039085743
+       0.3662386310913703
+ 5.26e+10    
+        0.367437882941899
+     -0.07735323262931347
+       0.3793208223486637
+    -0.009299119734933647
+       -0.037918275492843
+       0.3794903998281469
+    0.0002979521655082271
+    -0.009298908038725689
+     -0.07742734678666433
+       0.3667260748300562
+ 5.27e+10    
+       0.3679248294634591
+     -0.07752185512352452
+       0.3798816073522988
+    -0.009304809026143526
+     -0.03802732976904797
+       0.3800514310024025
+    0.0003443112285628918
+    -0.009304783760055025
+     -0.07759606443943988
+       0.3672124965334152
+ 5.28e+10    
+       0.3684107484386467
+     -0.07769049576319943
+       0.3804416103989869
+    -0.009310216255842062
+     -0.03813659172490989
+       0.3806116810943199
+    0.0003909003011320939
+     -0.00931037882290729
+      -0.0777648013586571
+       0.3676978957315629
+ 5.29e+10    
+       0.3688956394011855
+     -0.07785915253516698
+       0.3810008301096313
+    -0.009315340087728833
+     -0.03824606166680049
+       0.3811711487476969
+    0.0004377179890150947
+    -0.009315691891290605
+     -0.07793355554283815
+       0.3681822719533641
+ 5.3e+10     
+       0.3693795018834115
+     -0.07802782341550966
+       0.3815592651027888
+    -0.009320179192384421
+     -0.03835573990151967
+       0.3817298326038318
+    0.0004847628800748703
+    -0.009320721635993977
+     -0.07810232497972577
+        0.368665624726206
+ 5.31e+10    
+       0.3698623354160391
+     -0.07819650636973699
+       0.3821169139947561
+    -0.009324732247333422
+      -0.0384656267362766
+       0.3822877313016002
+    0.0005320335441897301
+    -0.009325466734649183
+     -0.07827110764645442
+       0.3691479535757698
+ 5.32e+10    
+       0.3703441395279226
+      -0.0783651993529584
+       0.3826737753996466
+    -0.009328997937107088
+     -0.03857572247866968
+       0.3828448434775342
+    0.0005795285332062829
+    -0.009329925871791905
+     -0.07843990150972693
+       0.3696292580258049
+ 5.33e+10    
+       0.3708249137458239
+      -0.0785339003100627
+       0.3832298479294791
+    -0.009332974953304421
+     -0.03868602743666794
+       0.3834011677659035
+    0.0006272463808937533
+    -0.009334097738922201
+     -0.07860870452599182
+       0.3701095375979011
+ 5.34e+10    
+       0.3713046575941768
+     -0.07870260717589787
+        0.383785130194264
+    -0.009336661994652839
+     -0.03879654191859072
+       0.3839567027987947
+    0.0006751856028997427
+    -0.009337981034563833
+     -0.07877751464162458
+       0.3705887918112641
+ 5.35e+10    
+       0.3717833705948504
+     -0.07887131787545273
+       0.3843396208020849
+    -0.009340057767067703
+     -0.03890726623308821
+       0.3845114472061951
+    0.0007233446967073529
+    -0.009341574464322617
+     -0.07894632979311007
+       0.3710670201824854
+ 5.36e+10    
+       0.3722610522669175
+     -0.07904003032404469
+       0.3848933183591936
+    -0.009343160983711027
+     -0.03901820068912171
+       0.3850653996160762
+    0.0007717221415938407
+    -0.009344876740944329
+     -0.07911514790722922
+       0.3715442222253202
+ 5.37e+10    
+       0.3727377021264162
+     -0.07920874242750521
+       0.3854462214700925
+    -0.009345970365049217
+     -0.03912934559594351
+       0.3856185586544791
+    0.0008203163985906674
+    -0.009347886584371089
+     -0.07928396690124766
+        0.372020397450459
+ 5.38e+10    
+       0.3732133196861188
+      -0.0793774520823725
+       0.3859983287376296
+    -0.009348484638909828
+     -0.03924070126307658
+       0.3861709229455988
+    0.0008691259104451905
+    -0.009350602721797351
+     -0.07945278468310615
+       0.3724955453653036
+ 5.39e+10    
+       0.3736879044552964
+     -0.07954615717608346
+       0.3865496387630877
+    -0.009350702540537553
+     -0.03935226800029498
+       0.3867224911118742
+    0.0009181491015838223
+    -0.009353023887724682
+     -0.07962159915161544
+       0.3729696654737419
+ 5.4e+10     
+       0.3741614559394859
+     -0.07971485558717051
+       0.3871001501462761
+    -0.009352622812649038
+     -0.03946404611760286
+       0.3872732617740742
+    0.0009673843780768222
+    -0.009355148824015527
+      -0.0797904081966522
+       0.3734427572759222
+ 5.41e+10    
+       0.3746339736402552
+      -0.0798835451854597
+       0.3876498614856267
+    -0.009354244205486901
+      -0.0395760359252145
+       0.3878232335513885
+     0.001016830127604684
+    -0.009356976279946468
+     -0.07995920969935835
+       0.3739148202680309
+ 5.42e+10    
+       0.3751054570549711
+     -0.08005222383227144
+       0.3881987713782869
+    -0.009355565476872758
+     -0.03968823773353402
+       0.3883724050615204
+     0.001066484719426216
+    -0.009358505012259962
+     -0.08012800153234292
+       0.3743858539420659
+ 5.43e+10    
+       0.3755759056765668
+     -0.08022088938062523
+       0.3887468784202173
+    -0.009356585392259253
+      -0.0398006518531344
+       0.3889207749207749
+     0.001116346504348252
+    -0.009359733785215657
+     -0.08029678155988701
+       0.3748558577856175
+ 5.44e+10    
+       0.3760453189933102
+     -0.08038953967544535
+       0.3892941812062861
+    -0.009357302724781167
+     -0.03991327859473726
+       0.3894683417441571
+     0.001166413814697129
+    -0.009360661370640341
+     -0.08046554763815014
+       0.3753248312816409
+ 5.45e+10    
+       0.3765136964885679
+     -0.08055817255376918
+        0.389840678330369
+    -0.009357716255305551
+     -0.04002611826919169
+       0.3900151041454617
+     0.001216684964291896
+    -0.009361286547977252
+     -0.08063429761537991
+       0.3757927739082362
+ 5.46e+10    
+        0.376981037640581
+     -0.08072678584496115
+       0.3903863683854513
+      -0.0093578247724807
+     -0.04013917118745475
+       0.3905610607373742
+     0.001267158248419228
+     -0.00936160810433416
+     -0.08080302933212621
+       0.3762596851384276
+ 5.47e+10    
+       0.3774473419222266
+     -0.08089537737092384
+       0.3909312499637231
+    -0.009357627072784562
+     -0.04025243766056924
+       0.3911062101315637
+     0.001317831943810333
+    -0.009361624834530714
+     -0.08097174062145426
+       0.3767255644399405
+ 5.48e+10    
+       0.3779126088007927
+     -0.08106394494631768
+       0.3914753216566856
+    -0.009357121960571674
+     -0.04036591799964388
+       0.3916505509387827
+     0.001368704308619527
+    -0.009361335541144699
+     -0.08114042930916313
+       0.3771904112749818
+ 5.49e+10    
+       0.3783768377377462
+     -0.08123248637877856
+       0.3920185820552519
+    -0.009356308248119361
+      -0.0404796125158326
+       0.3921940817689687
+     0.001419773582404647
+     -0.00936073903455701
+     -0.08130909321400687
+       0.3776542251000176
+ 5.5e+10     
+       0.3788400281885022
+     -0.08140099946914045
+       0.3925610297498516
+    -0.009355184755673025
+     -0.04059352152031315
+       0.3927368012313414
+     0.001471037986109658
+    -0.009359834132996592
+     -0.08147773014791666
+       0.3781170053655591
+ 5.51e+10    
+       0.3793021796021982
+     -0.08156948201166057
+       0.3931026633305358
+    -0.009353750311490142
+     -0.04070764532426691
+       0.3932787079345072
+      0.00152249572204881
+    -0.009358619662583067
+     -0.08164633791622654
+       0.3785787515159371
+ 5.52e+10    
+        0.379763291421463
+     -0.08173793179424609
+        0.393643481387084
+    -0.009352003751883522
+     -0.04082198423885752
+        0.393819800486561
+      0.00157414497389302
+     -0.00935709445736959
+     -0.08181491431790257
+       0.3790394629890906
+ 5.53e+10    
+       0.3802233630821912
+     -0.08190634659868452
+       0.3941834825091129
+    -0.009349943921263405
+     -0.04093653857521078
+        0.394360077495192
+     0.001625983906658189
+    -0.009355257359383855
+     -0.08198345714577299
+       0.3794991392163438
+ 5.54e+10    
+       0.3806823940133157
+     -0.08207472420087612
+       0.3947226652861805
+     -0.00934756967217866
+     -0.04105130864439314
+       0.3948995375677887
+     0.001678010666695413
+    -0.009353107218668583
+     -0.08215196418676242
+       0.3799577796221932
+ 5.55e+10    
+       0.3811403836365796
+     -0.08224306237106854
+       0.3952610283079026
+    -0.009344879865356731
+     -0.04116629475739181
+       0.3954381793115444
+     0.001730223381683456
+    -0.009350642893320767
+      -0.0823204332221279
+       0.3804153836240909
+ 5.56e+10    
+       0.3815973313663147
+     -0.08241135887409551
+       0.3957985701640583
+    -0.009341873369743065
+       -0.041281497225093
+        0.395976001333568
+     0.001782620160623122
+    -0.009347863249530236
+     -0.08248886202769772
+       0.3808719506322285
+ 5.57e+10    
+        0.382053236609212
+     -0.08257961146961681
+       0.3963352894447051
+    -0.009338549062538771
+      -0.0413969163582624
+       0.3965130022409915
+     0.001835199093833853
+    -0.009344767161616582
+     -0.08265724837411356
+       0.3813274800493238
+ 5.58e+10    
+       0.3825080987641006
+     -0.08274781791236063
+       0.3968711847402916
+    -0.009334905829237978
+     -0.04151255246752382
+       0.3970491806410801
+     0.001887958252952365
+    -0.009341353512065904
+     -0.08282559002707401
+       0.3817819712704083
+ 5.59e+10    
+       0.3829619172217235
+     -0.08291597595237045
+       0.3974062546417723
+     -0.00933094256366373
+     -0.04162840586333874
+       0.3975845351413452
+     0.001940895690933538
+    -0.009337621191565951
+     -0.08299388474758131
+       0.3822354236826118
+ 5.6e+10     
+       0.3834146913645154
+     -0.08308408333525173
+       0.3979404977407223
+    -0.009326658168003045
+     -0.04174447685598603
+       0.3981190643496569
+     0.001994009442053437
+    -0.009333569099040363
+     -0.08316213029219195
+       0.3826878366649545
+ 5.61e+10    
+       0.3838664205663812
+     -0.08325213780242405
+       0.3984739126294551
+    -0.009322051552840747
+     -0.04186076575554151
+        0.398652766874357
+     0.002047297521914619
+    -0.009329196141682041
+     -0.08333032441326721
+       0.3831392095881322
+ 5.62e+10    
+        0.384317104192474
+     -0.08342013709137341
+       0.3990064979011406
+    -0.009317121637192552
+     -0.04197727287185753
+       0.3991856413243772
+     0.002100757927453549
+    -0.009324501234985369
+      -0.0834984648592291
+         0.38358954181431
+ 5.63e+10    
+       0.3847667415989767
+     -0.08358807893590899
+       0.3995382521499243
+    -0.009311867348536869
+     -0.04209399851454296
+       0.3997176863093522
+     0.002154388636950478
+     -0.00931948330277765
+     -0.08366654937481702
+       0.3840388326969116
+ 5.64e+10    
+       0.3852153321328807
+     -0.08375596106642026
+       0.4000691739710458
+    -0.009306287622845704
+     -0.04221094299294254
+       0.4002489004397398
+     0.002208187610041461
+    -0.009314141277249053
+     -0.08383457570134747
+       0.3844870815804101
+ 5.65e+10    
+       0.3856628751317709
+      -0.0839237812101402
+       0.4005992619609636
+    -0.009300381404614404
+     -0.04232810661611753
+       0.4007792823269384
+     0.002262152787732785
+    -0.009308474098982146
+     -0.08400254157697712
+       0.3849342878001242
+ 5.66e+10    
+       0.3861093699236063
+       -0.084091537091407
+       0.4011285147174745
+    -0.009294147646890573
+     -0.04244548969282542
+       0.4013088305834094
+     0.002316282092417747
+    -0.009302480716979861
+     -0.08417044473696784
+       0.3853804506820091
+ 5.67e+10    
+       0.3865548158265026
+     -0.08425922643193101
+       0.4016569308398388
+    -0.009287585311301543
+     -0.04256309253150029
+       0.4018375438227956
+       0.0023705734278957
+     -0.00929616008869277
+     -0.08433828291395391
+       0.3858255695424531
+ 5.68e+10    
+       0.3869992121485211
+     -0.08442684695106423
+       0.4021845089289059
+    -0.009280693368081509
+     -0.04268091544023291
+       0.4023654206600459
+      0.00242502467939376
+    -0.009289511180045311
+     -0.08450605383821277
+       0.3862696436880739
+ 5.69e+10    
+       0.3874425581874497
+     -0.08459439636607001
+       0.4027112475872398
+    -0.009273470796096703
+     -0.04279895872675173
+       0.4028924597115386
+     0.002479633713590524
+    -0.009282532965460881
+     -0.08467375523793777
+       0.3867126724155155
+ 5.7e+10     
+       0.3878848532305931
+     -0.08476187239239856
+       0.4032371454192449
+    -0.009265916582870385
+     -0.04291722269840337
+       0.4034186595952067
+     0.002534398378642689
+      -0.0092752244278858
+     -0.08484138483951359
+       0.3871546550112451
+ 5.71e+10    
+       0.3883260965545585
+     -0.08492927274396206
+        0.403762201031296
+    -0.009258029724606215
+     -0.04303570766213276
+       0.4039440189306625
+      0.00258931650421385
+    -0.009267584558812726
+     -0.08500894036779369
+       0.3875955907513534
+ 5.72e+10    
+       0.3887662874250456
+     -0.08509659513341473
+       0.4042864130318675
+    -0.009249809226210815
+     -0.04315441392446527
+       0.4044685363393266
+     0.002644385901505798
+     -0.00925961235830239
+     -0.08517641954638197
+        0.388035478901356
+ 5.73e+10    
+       0.3892054250966369
+     -0.08526383727243324
+       0.4048097800316643
+    -0.009241254101315351
+     -0.04327334179148704
+       0.4049922104445564
+     0.002699604363292576
+    -0.009251306835004953
+     -0.08534382009791484
+       0.3884743187159941
+ 5.74e+10    
+       0.3896435088125862
+      -0.0854309968720013
+       0.4053323006437529
+    -0.009232363372295872
+     -0.04339249156882657
+       0.4055150398717748
+     0.002754969663956774
+    -0.009242667006179832
+     -0.08551113974434757
+       0.3889121094390371
+ 5.75e+10    
+       0.3900805378046144
+     -0.08559807164269591
+       0.4058539734836933
+    -0.009223136070292801
+     -0.04351186356163628
+        0.406037023248603
+     0.002810479559528558
+    -0.009233691897714669
+     -0.08567837620724195
+       0.3893488503030863
+ 5.76e+10    
+       0.3905165112927019
+     -0.08576505929497683
+       0.4063747971696766
+    -0.009213571235229276
+     -0.04363145807457421
+       0.4065581592049898
+     0.002866131787727297
+    -0.009224380544143596
+     -0.08584552720805738
+        0.389784540529381
+ 5.77e+10    
+       0.3909514284848803
+     -0.08593195753947706
+       0.4068947703226566
+    -0.009203667915828389
+     -0.04375127541178604
+       0.4070784463733479
+     0.002921924068005682
+    -0.009214731988663894
+     -0.08601259046844378
+       0.3902191793276042
+ 5.78e+10    
+       0.3913852885770319
+     -0.08609876408729784
+       0.4074138915664871
+    -0.009193425169629673
+      -0.0438713158768869
+       0.4075978833886866
+     0.002977854101596528
+    -0.009204745283152184
+     -0.08617956371053756
+       0.3906527658956912
+ 5.79e+10    
+       0.3918180907526844
+     -0.08626547665030446
+       0.4079321595280613
+    -0.009182842063004178
+     -0.04399157977294442
+       0.4081164688887482
+     0.003033919571562284
+    -0.009194419488179117
+     -0.08634644465725969
+       0.3910852994196364
+ 5.8e+10     
+       0.3922498341828098
+     -0.08643209294142529
+       0.4084495728374467
+    -0.009171917671168799
+     -0.04411206740246058
+       0.4086342015141443
+     0.003090118142847056
+    -0.009183753673023569
+     -0.08651323103261674
+        0.391516779073306
+ 5.81e+10    
+       0.3926805180256253
+     -0.08659861067495371
+       0.4089661301280295
+     -0.00916065107819935
+     -0.04423277906735518
+       0.4091510799084943
+     0.003146447462331493
+    -0.009172746915685356
+     -0.08667992056200334
+       0.3919472040182475
+ 5.82e+10    
+       0.3931101414263906
+     -0.08676502756685062
+       0.4094818300366501
+    -0.009149041377042883
+     -0.04435371506894858
+       0.4096671027185657
+      0.00320290515889013
+    -0.009161398302897129
+     -0.08684651097250887
+       0.3923765734035037
+ 5.83e+10    
+       0.3935387035172132
+     -0.08693134133505211
+       0.4099966712037501
+    -0.009137087669528601
+     -0.04447487570794511
+       0.4101822685944108
+     0.003259488843451767
+    -0.009149706930135408
+     -0.08701299999322468
+       0.3928048863654265
+ 5.84e+10    
+       0.3939662034168498
+     -0.08709754969977736
+       0.4105106522735119
+    -0.009124789066378083
+      -0.0445962612844169
+       0.4106965761895126
+     0.003316196109062216
+    -0.009137671901630248
+     -0.08717938535555517
+       0.3932321420274924
+ 5.85e+10    
+        0.394392640230513
+     -0.08726365038383979
+       0.4110237718940049
+    -0.009112144687214371
+     -0.04471787209778767
+       0.4112100241609267
+     0.003373024530950159
+    -0.009125292330374247
+     -0.08734566479353131
+       0.3936583395001196
+ 5.86e+10    
+        0.394818013049675
+     -0.08742964111296105
+       0.4115360287173302
+     -0.00909915366056982
+     -0.04483970844681682
+       0.4117226111694217
+     0.003429971666595447
+    -0.009112567338130401
+     -0.08751183604412438
+       0.3940834778804852
+ 5.87e+10    
+        0.395242320951876
+      -0.0875955196160859
+       0.4120474213997664
+    -0.009085815123893335
+     -0.04496177062958385
+       0.4122343358796283
+     0.003487035055800387
+    -0.009099496055438843
+     -0.08767789684756586
+       0.3945075562523451
+ 5.88e+10    
+       0.3956655630005337
+      -0.0877612836257016
+        0.412557948601917
+    -0.009072128223556289
+     -0.04508405894347346
+       0.4127451969601835
+     0.003544212220763826
+     -0.00908607762162281
+     -0.08784384494766649
+       0.3949305736858583
+ 5.89e+10    
+       0.3960877382447539
+     -0.08792693087815832
+        0.413067608988862
+    -0.009058092114857426
+     -0.04520657368516025
+       0.4132551930838789
+     0.003601500666157848
+    -0.009072311184793503
+     -0.08800967809213936
+       0.3953525292374039
+ 5.9e+10     
+        0.396508845719139
+     -0.08809245911399129
+       0.4135764012303034
+    -0.009043705962026824
+     -0.04532931515059444
+       0.4137643229278081
+     0.003658897879207467
+    -0.009058195901853918
+     -0.08817539403292468
+       0.3957734219494095
+ 5.91e+10    
+       0.3969288844436053
+      -0.0882578660782474
+       0.4140843240007191
+    -0.009028968938228977
+     -0.04545228363498737
+       0.4142725851735173
+      0.00371640132977316
+    -0.009043730938501632
+      -0.0883409905265178
+       0.3961932508501748
+ 5.92e+10    
+       0.3973478534231942
+     -0.08842314952081186
+        0.414591375979513
+    -0.009013880225564597
+     -0.04557547943279726
+       0.4147799785071553
+       0.0037740084704361
+    -0.009028915469230923
+     -0.08850646533429797
+       0.3966120149536986
+ 5.93e+10    
+       0.3977657516478919
+     -0.08858830719673937
+       0.4150975558511696
+    -0.008998439015071627
+     -0.04569890283771634
+       0.4152865016196265
+     0.003831716736586415
+    -0.009013748677333323
+      -0.0886718162228617
+       0.3970297132595081
+ 5.94e+10    
+       0.3981825780924419
+     -0.08875333686658479
+       0.4156028623054075
+    -0.008982644506725021
+     -0.04582255414265715
+       0.4157921532067439
+      0.00388952354651417
+    -0.008998229754897875
+     -0.08883704096435639
+       0.3974463447524879
+ 5.95e+10    
+       0.3985983317161687
+     -0.08891823629673984
+       0.4161072940373347
+    -0.008966495909435898
+     -0.04594643363973909
+         0.41629693196938
+     0.003947426301503341
+     -0.00898235790280999
+     -0.08900213733681668
+       0.3978619084027123
+ 5.96e+10    
+       0.3990130114627967
+     -0.08908300325976794
+        0.416610849747604
+    -0.008949992441049295
+      -0.0460705416202768
+       0.4168008366136279
+     0.004005422385928514
+    -0.008966132330749051
+     -0.08916710312450501
+       0.3982764031652776
+ 5.97e+10    
+       0.3994266162602711
+     -0.08924763553474485
+       0.4171135281425717
+    -0.008933133328341137
+     -0.04619487837476748
+       0.4173038658509536
+     0.004063509167354705
+    -0.008949552257185899
+     -0.08933193611825199
+        0.398689827980138
+ 5.98e+10    
+       0.3998391450205843
+     -0.08941213090759992
+       0.4176153279344561
+     -0.00891591780701418
+     -0.04631944419287896
+       0.4178060183983543
+     0.004121683996639917
+    -0.008932616909378587
+     -0.08949663411579932
+       0.3991021817719402
+ 5.99e+10    
+       0.4002505966395983
+     -0.08957648717145894
+       0.4181162478414959
+    -0.008898345121693097
+     -0.04644423936343833
+       0.4183072929785173
+     0.004179944208040608
+     -0.00891532552336749
+      -0.0896611949221473
+       0.3995134634498632
+ 6e+10       
+       0.4006609699968735
+     -0.08974070212699083
+       0.4186162865881111
+    -0.008880414525918208
+     -0.04656926417442122
+       0.4188076883199809
+     0.004238287119320154
+    -0.008897677343969207
+     -0.08982561634990208
+        0.399923671907455
+ 6.01e+10    
+       0.4010702639554971
+     -0.08990477358275549
+       0.4191154429050666
+    -0.008862125282138689
+     -0.04669451891294067
+       0.4193072031572929
+     0.004296710031860176
+    -0.008879671624770066
+     -0.08998989621962543
+       0.4003328060224769
+ 6.02e+10    
+       0.4014784773619129
+      -0.0900686993555542
+       0.4196137155296312
+    -0.008843476661704496
+     -0.04682000386523722
+        0.419805836231175
+     0.004355210230774825
+    -0.008861307628117942
+     -0.09015403236018858
+       0.4007408646567437
+ 6.03e+10    
+       0.4018856090457525
+     -0.09023247727078193
+       0.4201111032057461
+    -0.008824467944857417
+     -0.04694571931666892
+        0.420303586288684
+     0.004413784985027893
+    -0.008842584625113677
+     -0.09031802260912607
+       0.4011478466559693
+ 6.04e+10    
+       0.4022916578196686
+     -0.09039610516278197
+       0.4206076046841844
+    -0.008805098420721131
+     -0.04707166555170198
+       0.4208004520833776
+     0.004472431547553042
+     -0.00882350189560119
+     -0.09048186481299318
+       0.4015537508496123
+ 6.05e+10    
+       0.4026966224791727
+     -0.09055958087520313
+       0.4211032187227226
+    -0.008785367387290497
+     -0.04719784285390163
+       0.4212964323754775
+     0.004531147155376921
+    -0.008804058728157118
+     -0.09064555682772439
+       0.4019585760507241
+ 6.06e+10    
+       0.4031005018024684
+     -0.09072290226135798
+       0.4215979440863025
+    -0.008765274151419495
+     -0.04732425150592385
+       0.4217915259320395
+     0.004589929029744907
+    -0.008784254420078789
+      -0.0908090965189958
+       0.4023623210557983
+ 6.07e+10    
+       0.4035032945502919
+     -0.09088606718458471
+       0.4220917795472026
+    -0.008744818028808485
+     -0.04745089178950704
+       0.4222857315271154
+     0.004648774376250335
+    -0.008764088277372004
+     -0.09097248176258695
+       0.4027649846446202
+ 6.08e+10    
+       0.4039049994657522
+     -0.09104907351860936
+       0.4225847238852057
+    -0.008723998343990614
+     -0.04757776398546427
+        0.422779047941926
+     0.004707680384966191
+    -0.008743559614737512
+      -0.0911357104447473
+       0.4031665655801228
+ 6.09e+10    
+       0.4043056152741717
+     -0.09121191914791164
+       0.4230767758877684
+    -0.008702814430316936
+      -0.0477048683736765
+       0.4232714739650295
+     0.004766644230580018
+    -0.008722667755556447
+     -0.09129878046256404
+       0.4035670626082386
+ 6.1e+10     
+       0.4047051406829326
+     -0.09137460196809238
+       0.4235679343501944
+    -0.008681265629940912
+     -0.04783220523308547
+        0.423763008392491
+      0.00482566307253163
+    -0.008701412031875314
+     -0.09146168972433101
+       0.4039664744577576
+ 6.11e+10    
+       0.4051035743813184
+     -0.09153711988624198
+       0.4240581980758036
+    -0.008659351293801739
+      -0.0479597748416876
+       0.4242536500280553
+     0.004884734055153758
+    -0.008679791784389254
+      -0.0916244361499205
+        0.404364799840183
+ 6.12e+10    
+       0.4055009150403647
+     -0.09169947082131229
+       0.4245475658761065
+     -0.00863707078160705
+     -0.04808757747652787
+       0.4247433976833184
+     0.004943854307815833
+    -0.008657806362425633
+     -0.09178701767115756
+       0.4047620374495949
+ 6.13e+10    
+       0.4058971613127061
+     -0.09186165270449019
+       0.4250360365709794
+    -0.008614423461814133
+     -0.04821561341369513
+       0.4252322501779016
+     0.005003020945070243
+     -0.00863545512392525
+     -0.09194943223219509
+       0.4051581859625088
+ 6.14e+10    
+        0.406292311832428
+     -0.09202366347957257
+       0.4255236089888379
+    -0.008591408711611017
+     -0.04834388292831683
+       0.4257202063396285
+     0.005062231066802132
+    -0.008612737435423892
+     -0.09211167778989204
+       0.4055532440377391
+ 6.15e+10    
+       0.4066863652149184
+     -0.09218550110334313
+       0.4260102819668128
+    -0.008568025916895889
+     -0.04847238629455482
+       0.4262072650046968
+     0.005121481758381564
+    -0.008589652672032183
+     -0.09227375231419302
+       0.4059472103162664
+ 6.16e+10    
+       0.4070793200567239
+     -0.09234716354595297
+       0.4264960543509291
+    -0.008544274472256025
+     -0.04860112378560148
+       0.4266934250178578
+     0.005180770090818895
+    -0.008566200217415151
+     -0.09243565378850974
+       0.4063400834211029
+ 6.17e+10    
+       0.4074711749354029
+     -0.09250864879129984
+       0.4269809249962811
+    -0.008520153780945823
+     -0.04873009567367656
+       0.4271786852325937
+     0.005240093120923028
+    -0.008542379463770108
+      -0.0925973802101053
+       0.4067318619571616
+ 6.18e+10    
+       0.4078619284093871
+     -0.09266995483741342
+       0.4274648927672143
+    -0.008495663254863516
+     -0.04885930223002451
+        0.427663044511296
+      0.00529944789146246
+    -0.008518189811804664
+     -0.09275892959047891
+       0.4071225445111262
+ 6.19e+10    
+       0.4082515790178394
+     -0.09283107969683813
+       0.4279479565375029
+    -0.008470802314527645
+     -0.04898874372491156
+       0.4281465017254452
+     0.005358831431329315
+    -0.008493630670713032
+     -0.09292029995575361
+       0.4075121296513248
+ 6.2e+10     
+       0.4086401252805156
+     -0.09299202139702147
+       0.4284301151905328
+    -0.008445570389051972
+     -0.04911842042762511
+       0.4286290557557921
+     0.005418240755706249
+    -0.008468701458151772
+     -0.09308148934706598
+       0.4079006159276047
+ 6.21e+10    
+       0.4090275656976288
+     -0.09315277798070154
+       0.4289113676194815
+    -0.008419966916120059
+     -0.04924833260647157
+        0.429110705492539
+     0.005477672866236144
+    -0.008443401600214716
+     -0.09324249582095696
+       0.4082880018712063
+ 6.22e+10    
+        0.409413898749716
+     -0.09331334750629854
+        0.429391712727502
+    -0.008393991341958632
+      -0.0493784805287761
+       0.4295914498355236
+     0.005537124751194764
+    -0.008417730531406962
+     -0.09340331744976495
+       0.4086742859946436
+ 6.23e+10    
+       0.4097991228975018
+     -0.09347372804830664
+       0.4298711494279079
+    -0.008367643121309991
+     -0.04950886446088295
+       0.4300712876944013
+     0.005596593385666279
+     -0.00839168769461798
+     -0.09356395232202054
+       0.4090594667915827
+ 6.24e+10    
+       0.4101832365817721
+     -0.09363391769768736
+       0.4303496766443542
+    -0.008340921717403953
+     -0.04963948466815502
+         0.43055021798883
+     0.005656075731721396
+     -0.00836527254109388
+     -0.09372439854284288
+        0.409443542736724
+ 6.25e+10    
+       0.4105662382232425
+     -0.09379391456226638
+       0.4308272933110268
+     -0.00831382660192862
+     -0.04977034141497574
+       0.4310282396486571
+     0.005715568738598699
+    -0.008338484530408911
+     -0.09388465423433869
+       0.4098265122856859
+ 6.26e+10    
+       0.4109481262224322
+     -0.09395371676713053
+       0.4313039983728268
+    -0.008286357255000204
+     -0.04990143496475014
+       0.4315053516141046
+     0.005775069342888432
+    -0.008311323130435973
+     -0.09404471753600196
+       0.4102083738748912
+ 6.27e+10    
+       0.4113288989595406
+     -0.09411332245502715
+       0.4317797907855588
+    -0.008258513165132392
+     -0.05003276557990747
+       0.4319815528359578
+     0.005834574468719292
+    -0.008283787817316417
+     -0.09420458660511588
+       0.4105891259214532
+ 6.28e+10    
+       0.4117085547943204
+     -0.09427272978676499
+       0.4322546695161185
+     -0.00823029382920438
+     -0.05016433352190377
+       0.4324568422757525
+     0.005894081027947933
+    -0.008255878075428911
+     -0.09436425961715585
+       0.4109687668230663
+ 6.29e+10    
+       0.4120870920659613
+     -0.09443193694161688
+       0.4327286335426833
+     -0.00820169875242838
+     -0.05029613905122515
+       0.4329312189059654
+      0.00595358592035123
+    -0.008227593397357602
+      -0.0945237347661958
+       0.4113472949578968
+ 6.3e+10     
+       0.4124645090929682
+     -0.09459094211772398
+       0.4332016818548998
+    -0.008172727448316238
+      -0.0504281824273915
+        0.433404681710202
+     0.006013086033821358
+    -0.008198933283859336
+     -0.09468301026531357
+       0.4117247086844769
+ 6.31e+10    
+       0.4128408041730437
+     -0.09474974353250125
+       0.4336738134540778
+    -0.008143379438645003
+     -0.05056046390896221
+       0.4338772296833934
+     0.006072578244563357
+    -0.008169897243830026
+     -0.09484208434700089
+       0.4121010063415985
+ 6.32e+10    
+        0.413215975582974
+     -0.09490833942304533
+       0.4341450273533798
+    -0.008113654253422118
+     -0.05069298375353978
+        0.434348861831982
+     0.006132059417295874
+    -0.008140484794270346
+      -0.0950009552635724
+       0.4124761862482118
+ 6.33e+10    
+        0.413590021578516
+     -0.09506672804654387
+       0.4346153225780152
+    -0.008083551430849125
+      -0.0508257422177768
+       0.4348195771741169
+     0.006191526405454012
+    -0.008110695460250568
+     -0.09515962128757738
+       0.4128502467033238
+ 6.34e+10    
+       0.4139629403942854
+     -0.09522490768068469
+       0.4350846981654324
+    -0.008053070517285266
+     -0.05095873955738167
+         0.43528937473985
+     0.006250976051395388
+    -0.008080528774874567
+      -0.0953180807122137
+       0.4132231859858999
+ 6.35e+10    
+        0.414334730243647
+     -0.09538287662406937
+       0.4355531531655137
+    -0.008022211067209661
+     -0.05109197602712589
+       0.4357582535713261
+     0.006310405186608399
+    -0.008049984279242965
+     -0.09547633185174138
+       0.4135950023547659
+ 6.36e+10    
+       0.4147053893186095
+     -0.09554063319662638
+       0.4360206866407726
+    -0.007990972643183126
+     -0.05122545188085197
+       0.4362262127229833
+      0.00636981063192342
+    -0.008019061522415586
+     -0.09563437304189998
+       0.4139656940485137
+ 6.37e+10    
+       0.4150749157897173
+     -0.09569817574002544
+       0.4364872976665451
+    -0.007959354815808856
+     -0.05135916737148102
+       0.4366932512617456
+      0.00642918919772647
+    -0.007987760061373146
+     -0.09579220264032522
+       0.4143352592854077
+ 6.38e+10    
+       0.4154433078059488
+     -0.09585550261809436
+       0.4369529853311911
+    -0.007927357163692502
+     -0.05149312275102242
+       0.4371593682672216
+     0.006488537684175406
+    -0.007956079460977941
+      -0.0959498190269689
+       0.4147036962632953
+ 6.39e+10    
+       0.4158105634946168
+     -0.09601261221723764
+       0.4374177487362899
+    -0.007894979273401388
+      -0.0516273182705831
+       0.4376245628319039
+     0.006547852881418827
+    -0.007924019293934076
+     -0.09610722060451921
+       0.4150710031595159
+ 6.4e+10     
+       0.4161766809612659
+     -0.09616950294685427
+       0.4378815869968384
+    -0.007862220739422972
+     -0.05176175418037775
+       0.4380888340613651
+     0.006607131569817393
+    -0.007891579140746594
+     -0.09626440579882216
+       0.4154371781308136
+ 6.41e+10    
+        0.416541658289578
+     -0.09632617323975971
+       0.4383444992414505
+    -0.007829081164122405
+     -0.05189643072973955
+       0.4385521810744596
+     0.006666370520167556
+    -0.007858758589680164
+     -0.09642137305930594
+       0.4158022193132555
+ 6.42e+10    
+       0.4169054935412757
+      -0.0964826215526072
+       0.4388064846125598
+    -0.007795560157699427
+     -0.05203134816713254
+       0.4390146030035239
+     0.006725566493928092
+     -0.00782555723671664
+     -0.09657812085940415
+       0.4161661248221427
+ 6.43e+10    
+       0.4172681847560299
+     -0.09663884636631112
+       0.4392675422666147
+    -0.007761657338144609
+     -0.05216650674016261
+       0.4394760989945769
+     0.006784716243448674
+    -0.007791974685512185
+     -0.09673464769698324
+       0.4165288927519341
+ 6.44e+10    
+       0.4176297299513685
+     -0.09679484618647122
+       0.4397276713742852
+    -0.007727372331194331
+     -0.05230190669559127
+       0.4399366682075224
+      0.00684381651220111
+    -0.007758010547353441
+     -0.09689095209476881
+       0.4168905211761666
+ 6.45e+10    
+       0.4179901271225871
+     -0.09695061954379863
+       0.4401868711206602
+    -0.007692704770285793
+     -0.05243754827934893
+       0.4403963098163522
+     0.006902864035012933
+    -0.007723664441113055
+     -0.09704703260077391
+       0.4172510081473751
+ 6.46e+10    
+       0.4183493742426612
+     -0.09710616499454351
+       0.4406451407054573
+    -0.007657654296510307
+     -0.05257343173654967
+       0.4408550230093502
+     0.006961855538303405
+    -0.007688935993204314
+     -0.09720288778872999
+       0.4176103516970193
+ 6.47e+10    
+       0.4187074692621631
+     -0.09726148112092214
+         0.44110247934322
+    -0.007622220558566668
+     -0.05270955731150508
+       0.4413128069892951
+     0.007020787740321531
+    -0.007653824837535302
+     -0.09735851625851616
+       0.4179685498354105
+ 6.48e+10    
+       0.4190644101091778
+     -0.09741656653154662
+       0.4415588862635235
+     -0.00758640321271339
+     -0.05284592524774125
+       0.4417696609736669
+     0.007079657351386905
+    -0.007618330615461868
+     -0.09751391663659292
+       0.4183256005516407
+ 6.49e+10    
+       0.4194201946892214
+     -0.09757141986185611
+       0.4420143607111825
+    -0.007550201922720099
+     -0.05298253578801392
+       0.4422255841948508
+     0.007138461074132332
+    -0.007582452975740559
+     -0.09766908757643339
+       0.4186815018135109
+ 6.5e+10     
+       0.4197748208851628
+     -0.09772603977454723
+       0.4424689019464543
+    -0.007513616359818387
+     -0.05311938917432641
+       0.4426805759003469
+     0.007197195603748836
+    -0.007546191574479959
+      -0.0978240277589599
+       0.4190362515674675
+ 6.51e+10    
+       0.4201282865571486
+     -0.09788042496000807
+       0.4429225092452466
+    -0.007476646202652007
+     -0.05325648564794697
+       0.4431346353529743
+     0.007255857628233144
+    -0.007509546075092088
+      -0.0979787358929778
+       0.4193898477385345
+ 6.52e+10    
+       0.4204805895425237
+     -0.09803457413675021
+       0.4433751818993231
+    -0.007439291137225932
+     -0.05339382544942729
+       0.4435877618310803
+     0.007314443828636823
+      -0.0074725161482426
+      -0.0981332107156126
+       0.4197422882302519
+ 6.53e+10    
+       0.4208317276557638
+      -0.0981884860518453
+       0.4438269192165131
+    -0.007401550856855107
+     -0.05353140881862164
+       0.4440399546287481
+     0.007372950879317966
+    -0.007435101471800435
+     -0.09828745099274674
+        0.420093570924612
+ 6.54e+10    
+       0.4211816986884022
+     -0.09834215948135994
+       0.4442777205209195
+    -0.007363425062112354
+     -0.05366923599470717
+       0.4444912130560077
+     0.007431375448194728
+    -0.007397301730786733
+     -0.09844145551945901
+       0.4204436936820033
+ 6.55e+10    
+       0.4215305004089598
+      -0.0984955932307916
+        0.444727585153125
+    -0.007324913460775453
+      -0.0538073072162038
+       0.4449415364390434
+     0.007489714197001038
+    -0.007359116617323051
+     -0.09859522312046362
+       0.4207926543411507
+ 6.56e+10    
+       0.4218781305628816
+     -0.09864878613550787
+       0.4451765124704066
+    -0.007286015767773512
+     -0.05394562272099621
+       0.4453909241204068
+     0.007547963781544325
+    -0.007320545830578883
+     -0.09874875265055025
+       0.4211404507190625
+ 6.57e+10    
+       0.4222245868724696
+     -0.09880173706118366
+       0.4456245018469415
+    -0.007246731705132702
+     -0.05408418274635587
+       0.4458393754592255
+     0.007606120851965057
+    -0.007281589076718446
+     -0.09890204299502536
+       0.4214870806109746
+ 6.58e+10    
+       0.4225698670368204
+     -0.09895444490424113
+        0.446071552674021
+    -0.007207061001921503
+     -0.05422298752896369
+       0.4462868898314158
+     0.007664182052998491
+    -0.007242246068846823
+     -0.09905509307015464
+       0.4218325417903014
+ 6.59e+10    
+       0.4229139687317668
+     -0.09910690859228964
+       0.4465176643602592
+    -0.007167003394194693
+     -0.05436203730493342
+       0.4467334666298964
+     0.007722144024238103
+    -0.007202516526955379
+     -0.09920790182360598
+       0.4221768320085853
+ 6.6e+10     
+       0.4232568896098177
+     -0.09925912708456727
+       0.4469628363318065
+    -0.007126558624937119
+     -0.05450133230983646
+       0.4471791052647985
+     0.007780003400400868
+    -0.007162400177866447
+     -0.09936046823489247
+       0.4225199489954501
+ 6.61e+10    
+       0.4235986273001015
+      -0.0994110993723821
+       0.4474070680325622
+    -0.007085726444006625
+     -0.05464087277872672
+       0.4476238051636819
+     0.007837756811594669
+    -0.007121896755177414
+     -0.09951279131581819
+       0.4228618904585552
+ 6.62e+10    
+       0.4239391794083118
+     -0.09956282447955465
+       0.4478503589243887
+    -0.007044506608076219
+     -0.05478065894616628
+       0.4480675657717463
+     0.007895400883587023
+    -0.007081005999204217
+     -0.09966487011092195
+       0.4232026540835526
+ 6.63e+10    
+       0.4242785435166565
+     -0.09971430146286141
+       0.4482927084873205
+    -0.007002898880575814
+     -0.05492069104625217
+       0.4485103865520497
+     0.007952932238075902
+    -0.007039727656923817
+     -0.09981670369792459
+       0.4235422375340444
+ 6.64e+10    
+       0.4246167171838054
+     -0.09986552941247914
+       0.4487341162197845
+    -0.006960903031632645
+      -0.0550609693126438
+       0.4489522669857188
+     0.008010347492962026
+    -0.006998061481916402
+     -0.09996829118817513
+       0.4238806384515462
+ 6.65e+10    
+       0.4249536979448434
+      -0.1000165074524282
+       0.4491745816388087
+     -0.00691851883801205
+      -0.0552014939785907
+       0.4493932065721692
+     0.008067643262623023
+    -0.006956007234306673
+      -0.1001196317270975
+        0.424217854455446
+ 6.66e+10    
+       0.4252894833112245
+      -0.1001672347410188
+       0.4496141042802422
+    -0.006875746083056513
+     -0.05534226527696186
+       0.4498332048293174
+     0.008124816158188962
+    -0.006913564680704552
+      -0.1002707244946395
+       0.4245538831429718
+ 6.67e+10    
+       0.4256240707707249
+      -0.1003177104712964
+       0.4500526836989672
+    -0.006832584556624752
+     -0.05548328344027495
+       0.4502722612938008
+      0.00818186278781952
+    -0.006870733594145289
+      -0.1004215687057202
+       0.4248887220891561
+ 6.68e+10    
+       0.4259574577874046
+      -0.1004679338714878
+       0.4504903194691173
+    -0.006789034055029763
+     -0.05562454870072732
+       0.4507103755211928
+     0.008238779756982848
+    -0.006827513754028783
+      -0.1005721636106797
+       0.4252223688468059
+ 6.69e+10    
+       0.4262896418015641
+      -0.1006179042054479
+       0.4509270111842925
+    -0.006745094380976447
+     -0.05576606129022638
+       0.4511475470862196
+     0.008295563668735581
+    -0.006783904946058262
+      -0.1007225084957281
+       0.4255548209464714
+ 6.7e+10     
+       0.4266206202297067
+      -0.1007676207731069
+       0.4513627584577755
+    -0.006700765343498363
+     -0.05590782144042257
+       0.4515837755829824
+     0.008352211124004534
+    -0.006739906962178402
+      -0.1008726026833962
+       0.4258860758964201
+ 6.71e+10    
+       0.4269503904645057
+      -0.1009170829109191
+       0.4517975609227527
+    -0.006656046757894038
+     -0.05604982938274142
+       0.4520190606251708
+     0.008408718721869624
+    -0.006695519600512853
+      -0.1010224455329852
+       0.4262161311826094
+ 6.72e+10    
+       0.4272789498747641
+      -0.1010662899923086
+       0.4522314182325264
+    -0.006610938445662406
+     -0.05619208534841721
+       0.4524534018462832
+     0.008465083059848263
+    -0.006650742665300892
+      -0.1011720364410171
+       0.4265449842686638
+ 6.73e+10    
+       0.4276062958053874
+      -0.1012152414281204
+        0.452664330060738
+     -0.00656544023443777
+     -0.05633458956852784
+       0.4528867988998482
+     0.008521300734180875
+    -0.006605575966833624
+      -0.1013213748416879
+       0.4268726325958537
+ 6.74e+10    
+       0.4279324255773517
+      -0.1013639366670672
+       0.4530962961015814
+     -0.00651955195792418
+     -0.05647734227402908
+       0.4533192514596419
+      0.00857736834011774
+    -0.006560019321389537
+      -0.1014704602073168
+       0.4271990735830736
+ 6.75e+10    
+       0.4282573364876741
+      -0.1015123751961797
+       0.4535273160700263
+    -0.006473273455828715
+     -0.05662034369579128
+       0.4537507592199074
+     0.008633282472206891
+    -0.006514072551169313
+      -0.1016192920487988
+       0.4275243046268241
+ 6.76e+10    
+       0.4285810258093887
+      -0.1016605565412551
+       0.4539573897020354
+    -0.006426604573794853
+     -0.05676359406463609
+       0.4541813218955787
+      0.00868903972458347
+    -0.006467735484230076
+       -0.101767869916058
+       0.4278483231011987
+ 6.77e+10    
+       0.4289034907915206
+      -0.1018084802673077
+       0.4543865167547835
+    -0.006379545163334495
+     -0.05690709361137338
+       0.4546109392224967
+     0.008744636691259822
+    -0.006421007954419128
+      -0.1019161933984979
+       0.4281711263578657
+ 6.78e+10    
+        0.429224728659065
+      -0.1019561459790178
+       0.4548146970068776
+    -0.006332095081759947
+     -0.05705084256684033
+       0.4550396109576343
+     0.008800069966416624
+    -0.006373889801306768
+      -0.1020642621254552
+       0.4284927117260586
+ 6.79e+10    
+       0.4295447366129633
+      -0.1021035533211816
+       0.4552419302585767
+     -0.00628425419211473
+     -0.05719484116193992
+       0.4554673368793135
+     0.008855336144695306
+    -0.006326380870118792
+       -0.102212075766652
+       0.4288130765125629
+ 6.8e+10     
+       0.4298635118300906
+      -0.1022507019791627
+       0.4556682163320134
+    -0.006236022363104354
+     -0.05733908962768153
+       0.4558941167874325
+     0.008910431821491272
+    -0.006278481011668219
+      -0.1023596340326496
+       0.4291322180017111
+ 6.81e+10    
+       0.4301810514632319
+      -0.1023975916793397
+       0.4560935550714112
+    -0.006187399469025899
+     -0.05748358819522117
+       0.4563199505036827
+     0.008965353593247738
+    -0.006230190082286409
+      -0.1025069366752993
+       0.4294501334553721
+ 6.82e+10    
+       0.4304973526410737
+      -0.1025442221895595
+        0.456517946343311
+    -0.006138385389697258
+     -0.05762833709590367
+       0.4567448378717731
+     0.009020098057750689
+    -0.006181507943753594
+      -0.1026539834881973
+       0.4297668201129488
+ 6.83e+10    
+        0.430812412468187
+      -0.1026905933195849
+       0.4569413900367859
+    -0.006088980010385901
+     -0.05777333656130443
+       0.4571687787576518
+     0.009074661814424612
+    -0.006132434463228801
+      -0.1028007743071367
+       0.4300822751913732
+ 6.84e+10    
+       0.4311262280250197
+      -0.1028367049215464
+       0.4573638860636666
+    -0.006039183221736758
+     -0.05791858682327302
+       0.4575917730497297
+     0.009129041464628739
+    -0.006082969513179145
+      -0.1029473090105601
+       0.4303964958851063
+ 6.85e+10    
+       0.4314387963678836
+      -0.1029825568903913
+       0.4577854343587606
+    -0.005988994919699554
+     -0.05806408811397719
+       0.4580138206591021
+     0.009183233611954262
+    -0.006033112971308578
+      -0.1030935875200136
+       0.4307094793661388
+ 6.86e+10    
+       0.4317501145289515
+      -0.1031281491643354
+       0.4582060348800762
+    -0.005938415005455605
+     -0.05820984066594793
+       0.4584349215197737
+     0.009237234862521849
+    -0.005982864720485885
+      -0.1032396098005985
+       0.4310212227839924
+ 6.87e+10    
+       0.4320601795162496
+      -0.1032734817253107
+       0.4586256876090414
+    -0.005887443385344105
+     -0.05835584471212452
+        0.458855075588878
+     0.009291041825280013
+    -0.005932224648672336
+      -0.1033853758614243
+       0.4313317232657241
+ 6.88e+10    
+       0.4323689883136537
+      -0.1034185545994168
+       0.4590443925507278
+    -0.005836079970787525
+     -0.05850210048590185
+       0.4592742828469054
+     0.009344651112303573
+    -0.005881192648848307
+      -0.1035308857560612
+       0.4316409779159319
+ 6.89e+10    
+       0.4326765378808894
+      -0.1035633678573704
+       0.4594621497340731
+    -0.005784324678216612
+     -0.05864860822117736
+       0.4596925432979239
+      0.00939805933909324
+    -0.005829768618939891
+      -0.1036761395829926
+       0.4319489838167646
+ 6.9e+10     
+        0.432982825153531
+      -0.1037079216149533
+       0.4598789592120996
+    -0.005732177428994905
+      -0.0587953681523988
+       0.4601098569698016
+     0.009451263124874897
+    -0.005777952461744457
+      -0.1038211374860659
+       0.4322557380279266
+ 6.91e+10    
+       0.4332878470430048
+      -0.1038522160334633
+       0.4602948210621423
+    -0.005679638149342178
+     -0.05894238051461435
+       0.4605262239144337
+     0.009504259092899592
+     -0.00572574408485577
+      -0.1039658796549458
+       0.4325612375866946
+ 6.92e+10    
+       0.4335916004365921
+      -0.1039962513201621
+       0.4607097353860668
+    -0.005626706770257959
+     -0.05908964554352134
+       0.4609416442079641
+     0.009557043870744008
+    -0.005673143400588471
+      -0.1041103663255647
+       0.4328654795079251
+ 6.93e+10    
+       0.4338940821974335
+      -0.1041400277287225
+       0.4611237023104924
+    -0.005573383227443982
+      -0.0592371634755173
+       0.4613561179510092
+     0.009609614090610482
+    -0.005620150325902077
+      -0.1042545977805739
+       0.4331684607840728
+ 6.94e+10    
+       0.4341952891645405
+      -0.1042835455596786
+       0.4615367219870153
+    -0.005519667461226084
+     -0.05938493454775191
+       0.4617696452688839
+     0.009661966389628126
+    -0.005566764782324379
+      -0.1043985743497947
+       0.4334701783852064
+ 6.95e+10    
+       0.4344952181528002
+      -0.1044268051608719
+       0.4619487945924324
+     -0.00546555941647576
+     -0.05953295899817848
+       0.4621822263118222
+     0.009714097410153187
+     -0.00551298669587404
+      -0.1045422964106673
+       0.4337706292590235
+ 6.96e+10    
+         0.43479386595299
+      -0.1045698069278986
+       0.4623599203289606
+    -0.005411059042530961
+     -0.05968123706560789
+       0.4625938612552054
+     0.009766003800070165
+     -0.00545881599698299
+      -0.1046857643887029
+       0.4340698103308743
+ 6.97e+10    
+       0.4350912293317874
+      -0.1047125513045569
+        0.462770099424461
+    -0.005356166293116317
+     -0.05982976898976206
+       0.4630045502997817
+     0.009817682213092503
+    -0.005404252620417788
+      -0.1048289787579298
+       0.4343677185037799
+ 6.98e+10    
+       0.4353873050317857
+      -0.1048550387832915
+       0.4631793321326616
+    -0.005300881126262789
+     -0.05997855501132893
+       0.4634142936718921
+     0.009869129309063408
+    -0.005349296505200947
+      -0.1049719400413445
+        0.434664350658456
+ 6.99e+10    
+       0.4356820897715125
+      -0.1049972699056416
+       0.4635876187333802
+    -0.005245203504226736
+     -0.06012759537201869
+        0.463823091623697
+     0.009920341754256681
+    -0.005293947594531066
+      -0.1051146488113592
+       0.4349597036533392
+ 7e+10       
+        0.435975580245442
+      -0.1051392452626825
+       0.4639949595327433
+    -0.005189133393408644
+     -0.06027689031461914
+       0.4642309444333952
+     0.009971316221677054
+    -0.005238205835702979
+      -0.1052571056902485
+       0.4352537743246102
* NOTE: Solution at 1e+08 Hz used as DC point.

.model c_m4lines_HFSS_W_1 sp N=4 SPACING=nonuniform VALTYPE=real
+ INTERPOLATION=spline
+ INFINITY =
+    7.938621322074103e-11
+   -2.234686778922564e-11
+    8.350721157248263e-11
+   -1.872746540418529e-12
+   -1.142445181304755e-11
+    8.352938776572516e-11
+   -2.203335273976321e-13
+   -1.872043010176729e-12
+   -2.235002713338225e-11
+     7.92698254841625e-11
+ DATA = 700
+ 0           
+    8.640174920590117e-11
+    -2.14416090728894e-11
+    8.793408763567512e-11
+   -8.389673395611541e-13
+   -1.021175218891604e-11
+    8.796128153242538e-11
+   -3.023047060529615e-13
+   -8.359493564182524e-13
+   -2.144637104119777e-11
+    8.625786243188311e-11
+ 2e+08       
+    8.579356517807833e-11
+   -2.133018481287351e-11
+    8.732273804978702e-11
+   -8.409745571171349e-13
+   -1.015945392081564e-11
+    8.734928774723289e-11
+   -3.017209077407336e-13
+   -8.379727382415652e-13
+   -2.133396863163589e-11
+    8.565048805585838e-11
+ 3e+08       
+    8.543439129147498e-11
+   -2.125919358636875e-11
+    8.696147697909173e-11
+   -8.388714817469942e-13
+   -1.013212095931011e-11
+    8.698809761386621e-11
+   -3.016053761501185e-13
+   -8.358583481642005e-13
+   -2.126333912016844e-11
+    8.529262847560166e-11
+ 4e+08       
+     8.51973785006239e-11
+   -2.121611624896911e-11
+    8.672397360039697e-11
+   -8.370576263106825e-13
+    -1.01144905578764e-11
+    8.675056048629885e-11
+   -3.015461469017349e-13
+   -8.340441696890575e-13
+   -2.122041112324275e-11
+    8.505609369460387e-11
+ 5e+08       
+    8.501308142501136e-11
+   -2.118240268346723e-11
+    8.653926817497166e-11
+   -8.358747223385644e-13
+   -1.009992154090721e-11
+    8.656576400727495e-11
+   -3.012893316516853e-13
+   -8.328633203687275e-13
+   -2.118669760698499e-11
+    8.487204370126886e-11
+ 6e+08       
+    8.485906137203432e-11
+    -2.11533346653181e-11
+    8.638463937856391e-11
+   -8.349758688101932e-13
+   -1.008711758231931e-11
+    8.641104847680747e-11
+   -3.008173216221576e-13
+   -8.319664423778381e-13
+   -2.115758882075701e-11
+     8.47182727872951e-11
+ 7e+08       
+    8.472695307073616e-11
+   -2.112780632516672e-11
+    8.625179551406494e-11
+   -8.341174077938374e-13
+   -1.007578659555687e-11
+    8.627813731849719e-11
+   -3.001762091430381e-13
+   -8.311096585892238e-13
+   -2.113201709725078e-11
+     8.45864327515991e-11
+ 8e+08       
+    8.461229945786495e-11
+   -2.110531332881669e-11
+    8.613639890603737e-11
+   -8.331937424130681e-13
+   -1.006572106061007e-11
+    8.616268716773436e-11
+   -2.994151589074017e-13
+   -8.301876066807383e-13
+   -2.110948556650975e-11
+    8.447203040662894e-11
+ 9e+08       
+    8.451184222347195e-11
+   -2.108535962900842e-11
+    8.603526482545168e-11
+   -8.321766378163135e-13
+    -1.00566835807289e-11
+    8.606150428414358e-11
+    -2.98570621181589e-13
+   -8.291723195167683e-13
+   -2.108949872180673e-11
+    8.437178184932172e-11
+ 1e+09       
+    8.442288424772558e-11
+   -2.106742960264604e-11
+    8.594571214091148e-11
+   -8.310706423844269e-13
+    -1.00484331775308e-11
+    8.597190206687965e-11
+   -2.976659995362326e-13
+   -8.280685677340599e-13
+   -2.107154255125035e-11
+    8.428298725200001e-11
+ 1.1e+09     
+    8.437460507791684e-11
+   -2.106624074547515e-11
+    8.589805476139957e-11
+   -8.239465012216544e-13
+   -1.004552064913586e-11
+    8.592413259584436e-11
+   -2.964899427887409e-13
+   -8.209940977364336e-13
+   -2.107014523867967e-11
+    8.423447568500969e-11
+ 1.2e+09     
+     8.43245663974042e-11
+   -2.106233839222982e-11
+    8.584835482871661e-11
+   -8.176495839037098e-13
+   -1.004129128696384e-11
+    8.587432691337147e-11
+   -2.950683251965018e-13
+   -8.147242930860823e-13
+   -2.106605289143358e-11
+    8.418423233417252e-11
+ 1.3e+09     
+    8.427348347863223e-11
+   -2.105619764460884e-11
+    8.579737854348914e-11
+   -8.120816160966631e-13
+   -1.003609607263911e-11
+    8.582325255344668e-11
+   -2.934383948906261e-13
+   -8.091670836177758e-13
+   -2.105974252581142e-11
+    8.413297630310995e-11
+ 1.4e+09     
+    8.422198447874124e-11
+   -2.104826086692808e-11
+    8.574579286412157e-11
+   -8.071507419404161e-13
+   -1.003020671643005e-11
+     8.57715772640569e-11
+   -2.916359239640621e-13
+   -8.042356180334973e-13
+   -2.105165715359212e-11
+    8.408133775151999e-11
+ 1.5e+09     
+    8.417060450730928e-11
+   -2.103892206532189e-11
+    8.569416348395644e-11
+   -8.027736976958999e-13
+   -1.002383528259889e-11
+     8.57198671152423e-11
+   -2.896942242071174e-13
+   -7.998505001503724e-13
+   -2.104219055273919e-11
+    8.402985227937574e-11
+ 1.6e+09     
+    8.411978678206185e-11
+   -2.102852170767522e-11
+    8.564295849298016e-11
+   -7.988765243830525e-13
+   -1.001714788028125e-11
+    8.566859026324317e-11
+   -2.876435674601692e-13
+    -7.95940665847512e-13
+   -2.103168238190677e-11
+    8.397896239793878e-11
+ 1.7e+09     
+    8.406988822017556e-11
+   -2.101734750701204e-11
+    8.559255557568778e-11
+   -7.953943938286889e-13
+   -1.001027455692468e-11
+     8.56181242275682e-11
+   -2.855109252620918e-13
+   -7.924433978815882e-13
+   -2.102041917795803e-11
+    8.392902341443424e-11
+ 1.8e+09     
+    8.402118754988145e-11
+   -2.100563833763528e-11
+    8.554325115714106e-11
+   -7.922709571671941e-13
+   -1.000331669784981e-11
+    8.556876509874973e-11
+   -2.833199379111761e-13
+    -7.89303850394293e-13
+   -2.100863842489831e-11
+    8.388031180405749e-11
+ 1.9e+09     
+       8.397389460195e-11
+   -2.099358956582531e-11
+    8.549527036746823e-11
+   -7.894574809001196e-13
+   -9.996352726713894e-12
+    8.552073755158072e-11
+    -2.81091036365744e-13
+   -7.864743338712114e-13
+   -2.099653399236813e-11
+    8.383303472394389e-11
+ 2e+09       
+    8.392815987371647e-11
+   -2.098135879148791e-11
+    8.544877705245908e-11
+   -7.869119293487982e-13
+   -9.989442599220102e-12
+    8.547420489465154e-11
+   -2.788416580462351e-13
+    -7.83913516778218e-13
+   -2.098426195255009e-11
+    8.378733976081267e-11
+ 2.1e+09     
+    8.388408377819229e-11
+   -2.096907144194183e-11
+    8.540388332881279e-11
+   -7.845980810007209e-13
+   -9.982631403961308e-12
+    8.542927865685387e-11
+   -2.765865138451134e-13
+   -7.815856340359866e-13
+   -2.097194622573455e-11
+    8.374332432653029e-11
+ 2.2e+09     
+    8.384172522303675e-11
+   -2.095682592970669e-11
+    8.536065838308113e-11
+   -7.824847214995741e-13
+   -9.975952278494238e-12
+    8.538602741130715e-11
+   -2.743378767379694e-13
+   -7.794597495733617e-13
+   -2.095968377287441e-11
+     8.37010443497313e-11
+ 2.3e+09     
+    8.380110932925539e-11
+   -2.094469824741965e-11
+    8.531913635788977e-11
+   -7.805449295475684e-13
+   -9.969428785070778e-12
+    8.534448468130195e-11
+   -2.721058722469524e-13
+   -7.775090938887741e-13
+   -2.094754921288971e-11
+     8.36605220776313e-11
+ 2.4e+09     
+     8.37622342136142e-11
+   -2.093274596658718e-11
+    8.527932326991699e-11
+   -7.787554572719812e-13
+    -9.96307685112063e-12
+    8.530465587353196e-11
+    -2.69898758150362e-13
+    -7.75710482305071e-13
+   -2.093559883478369e-11
+    8.362175291662427e-11
+ 2.5e+09     
+     8.37250768346537e-11
+   -2.092101165898519e-11
+    8.524120297159354e-11
+    -7.77096199101624e-13
+   -9.956906354343927e-12
+    8.526652425124387e-11
+   -2.677231858773431e-13
+   -7.740438113589374e-13
+   -2.092387402584967e-11
+    8.358471131607552e-11
+ 2.6e+09     
+    8.368959794989149e-11
+   -2.090952578645482e-11
+     8.52047422109606e-11
+   -7.755497399184461e-13
+   -9.950922415282258e-12
+    8.523005600234436e-11
+   -2.655844395192381e-13
+   -7.724916267588425e-13
+   -2.091240416355471e-11
+    8.354935574709566e-11
+ 2.7e+09     
+    8.365574625922425e-11
+   -2.089830911669424e-11
+    8.516989486837121e-11
+   -7.741009723267556e-13
+   -9.945126448164106e-12
+    8.519520448168605e-11
+    -2.63486650759463e-13
+   -7.710387547948227e-13
+   -2.090120903008251e-11
+    8.351563285501788e-11
+ 2.8e+09     
+    8.362346182275519e-11
+   -2.088737472565504e-11
+    8.513660546009465e-11
+   -7.727367731910079e-13
+   -9.939517011781159e-12
+     8.51619137180878e-11
+   -2.614329895931576e-13
+    -7.69671988883333e-13
+   -2.089030081118862e-11
+    8.348348087697058e-11
+ 2.9e+09     
+    8.359267884491582e-11
+   -2.087672964517384e-11
+    8.510481200153078e-11
+   -7.714457304773174e-13
+   -9.934090495075022e-12
+    8.513012127922784e-11
+   -2.594258317109687e-13
+   -7.683798234194198e-13
+   -2.087968573878684e-11
+    8.345283241904081e-11
+ 3e+09       
+    8.356332791425514e-11
+   -2.086637620987677e-11
+     8.50744483197437e-11
+   -7.702179125270195e-13
+    -9.92884166638844e-12
+    8.509976058450765e-11
+   -2.574669040275244e-13
+   -7.671522279005185e-13
+   -2.086936543189445e-11
+    8.342361668451188e-11
+ 3.1e+09     
+    8.353533778210108e-11
+   -2.085631315162771e-11
+    8.504544589867172e-11
+   -7.690446729987935e-13
+   -9.923764110602195e-12
+    8.507076274956859e-11
+   -2.555574101657824e-13
+   -7.659804551695532e-13
+   -2.085933798464651e-11
+      8.3395761238047e-11
+ 3.2e+09     
+    8.350863675521079e-11
+   -2.084653648371604e-11
+    8.501773533224297e-11
+   -7.679184857435841e-13
+   -9.918850574420401e-12
+    8.504305803796828e-11
+   -2.536981378506696e-13
+   -7.648568784863931e-13
+    -2.08495988438939e-11
+    8.336919338220913e-11
+ 3.3e+09     
+    8.348315376867641e-11
+   -2.083704021108556e-11
+    8.499124745182819e-11
+   -7.668328047854111e-13
+   -9.914093236740164e-12
+    8.501657698667354e-11
+   -2.518895501817527e-13
+   -7.637748529231612e-13
+   -2.084014151291486e-11
+    8.334384121353976e-11
+ 3.4e+09     
+    8.345881919651734e-11
+   -2.082781689745869e-11
+    8.496591418570073e-11
+   -7.657819453618638e-13
+   -9.909483918246677e-12
+    8.499125126322584e-11
+   -2.501318626896018e-13
+   -7.627285972702954e-13
+   -2.083095811225276e-11
+    8.331963441632407e-11
+ 3.5e+09     
+    8.343556544902443e-11
+   -2.081885811533263e-11
+    8.494166919988745e-11
+   -7.647609826364102e-13
+   -9.905014242034174e-12
+    8.496701430410684e-11
+   -2.484251079656327e-13
+   -7.617130932333311e-13
+   -2.082203982376043e-11
+    8.329650484359301e-11
+ 3.6e+09     
+    8.341332739827877e-11
+   -2.081015480054896e-11
+    8.491844836222584e-11
+   -7.637656652429803e-13
+   -9.900675755104275e-12
+     8.49438017762299e-11
+   -2.467691895129345e-13
+   -7.607239992017769e-13
+   -2.081337723961679e-11
+     8.32743869271183e-11
+ 3.7e+09     
+    8.339204266647787e-11
+   -2.080169752945212e-11
+    8.489619006469673e-11
+   -7.627923412763014e-13
+   -9.896460018983533e-12
+    8.492155189671331e-11
+   -2.451639263111069e-13
+   -7.597575762896345e-13
+   -2.080496063436553e-11
+      8.3253217951232e-11
+ 3.8e+09     
+    8.337165180576088e-11
+   -2.079347673351197e-11
+    8.487483543321042e-11
+   -7.618378947130726e-13
+   -9.892358676382076e-12
+     8.49002056401747e-11
+   -2.436090894320529e-13
+   -7.588106246944749e-13
+   -2.079678017486359e-11
+    8.323293821928147e-11
+ 3.9e+09     
+    8.335209839313658e-11
+   -2.078548286363725e-11
+    8.485432844894897e-11
+   -7.608996905526249e-13
+   -9.888363499745811e-12
+    8.487970685769248e-11
+   -2.421044318926161e-13
+   -7.578804287071768e-13
+    -2.07888260803635e-11
+    8.321349113636718e-11
+ 4e+09       
+    8.333332905977977e-11
+    -2.07777065141868e-11
+    8.483461600105146e-11
+   -7.599755272126889e-13
+   -9.884466426696411e-12
+    8.486000232725074e-11
+   -2.406497127882133e-13
+   -7.569647089387849e-13
+   -2.078108874272305e-11
+    8.319482322762901e-11
+ 4.1e+09     
+    8.331529347032924e-11
+    -2.07701385148415e-11
+    8.481564788679407e-11
+     -7.5906359491642e-13
+   -9.880659586670524e-12
+     8.48410417518371e-11
+   -2.392447166213628e-13
+   -7.560615805219996e-13
+   -2.077355881488424e-11
+    8.317688410767872e-11
+ 4.2e+09     
+    8.329794426478199e-11
+   -2.076276999696981e-11
+    8.479737677237883e-11
+   -7.581624389698094e-13
+   -9.876935322531008e-12
+    8.482277771831569e-11
+   -2.378892686213871e-13
+    -7.55169516201203e-13
+   -2.076622727422989e-11
+    8.315962641371717e-11
+ 4.3e+09     
+    8.328123697306673e-11
+   -2.075559243986129e-11
+    8.477975812492582e-11
+   -7.572709269620781e-13
+   -9.873286210493813e-12
+    8.480516562767506e-11
+   -2.365832467462516e-13
+   -7.542873133536138e-13
+   -2.075908546616508e-11
+    8.314300571235097e-11
+ 4.4e+09     
+    8.326512991031394e-11
+   -2.074859770116746e-11
+    8.476275012418314e-11
+   -7.563882190330851e-13
+   -9.869705081362319e-12
+    8.478816360515985e-11
+   -2.353265909642827e-13
+    -7.53414064092236e-13
+   -2.075212513223451e-11
+    8.312698038804697e-11
+ 4.5e+09     
+    8.324958405915143e-11
+   -2.074177803504395e-11
+    8.474631356075768e-11
+   -7.555137404484584e-13
+    -9.86618504575115e-12
+    8.477173239708613e-11
+   -2.341193103307798e-13
+   -7.525491276955131e-13
+   -2.074533842624111e-11
+    8.311151151947351e-11
+ 4.6e+09     
+    8.323456294397341e-11
+   -2.073512610079575e-11
+    8.473041172626343e-11
+   -7.546471558120446e-13
+   -9.862719525675323e-12
+    8.475583525972882e-11
+   -2.329614883011739e-13
+    -7.51692104695937e-13
+   -2.073871792114108e-11
+    8.309656274859854e-11
+ 4.7e+09     
+    8.322003250102418e-11
+   -2.072863496426713e-11
+    8.471501029962669e-11
+   -7.537883443344915e-13
+   -9.859302294537604e-12
+    8.474043784450956e-11
+   -2.318532866564696e-13
+   -7.508428120477884e-13
+   -2.073225660892985e-11
+    8.308210014630609e-11
+ 4.8e+09     
+     8.32059609472368e-11
+   -2.072229809376132e-11
+    8.470007723282714e-11
+   -7.529373756728991e-13
+   -9.855927527122391e-12
+    8.472550808275479e-11
+   -2.307949483566619e-13
+   -7.500012588896035e-13
+   -2.072594789527999e-11
+    8.306809207739955e-11
+ 4.9e+09     
+     8.31923186500486e-11
+   -2.071610935190722e-11
+    8.468558263854508e-11
+   -7.520944859681707e-13
+   -9.852589860653958e-12
+    8.471101607248576e-11
+   -2.297867995813312e-13
+   -7.491676225281557e-13
+   -2.071978559032449e-11
+    8.305450906714383e-11
+ 5e+09       
+    8.317907799984759e-11
+   -2.071006298459431e-11
+    8.467149868150085e-11
+   -7.512600538401991e-13
+   -9.849284467257982e-12
+    8.469693396900967e-11
+   -2.288292511624622e-13
+    -7.48342224403974e-13
+   -2.071376389668501e-11
+    8.304132367093616e-11
+ 5.1e+09     
+    8.316621328624557e-11
+   -2.070415360785845e-11
+    8.465779947465871e-11
+   -7.504345762623582e-13
+   -9.846007137244163e-12
+    8.468323588048167e-11
+   -2.279227995607326e-13
+   -7.475255059592271e-13
+   -2.070787739560884e-11
+     8.30285103482446e-11
+ 5.2e+09     
+    8.315370057902299e-11
+   -2.069837619341264e-11
+    8.464446098092966e-11
+   -7.496186444285036e-13
+   -9.842754371488154e-12
+    8.466989776905474e-11
+   -2.270680274821684e-13
+   -7.467180045210113e-13
+   -2.070212103188863e-11
+    8.301604534160405e-11
+ 5.3e+09     
+    8.314151761431461e-11
+   -2.069272605336643e-11
+    8.463146092050412e-11
+     -7.4881291994669e-13
+   -9.839523479845461e-12
+    8.465689735774398e-11
+   -2.262656041769715e-13
+   -7.459203295333745e-13
+   -2.069649009809338e-11
+    8.300390656119107e-11
+ 5.4e+09     
+    8.312964368638912e-11
+   -2.068719882455853e-11
+    8.461877868348323e-11
+   -7.480181119364553e-13
+   -9.836312681026916e-12
+    8.464421404266127e-11
+   -2.255162854068487e-13
+   -7.451331397145541e-13
+    -2.06909802185182e-11
+    8.299207347528808e-11
+ 5.5e+09     
+    8.311805954521732e-11
+   -2.068179045283539e-11
+    8.460639524705884e-11
+   -7.472349558550189e-13
+   -9.833121197811067e-12
+    8.463182880986402e-11
+   -2.248209130136789e-13
+   -7.443571219641143e-13
+   -2.068558733317268e-11
+    8.298052700679099e-11
+ 5.6e+09     
+     8.31067472999018e-11
+   -2.067649717753492e-11
+    8.459429309612675e-11
+    -7.46464195109326e-13
+   -9.829949340016967e-12
+    8.461972415569466e-11
+   -2.241804139738643e-13
+   -7.435929730763689e-13
+   -2.068030768205328e-11
+     8.29692494358001e-11
+ 5.7e+09     
+    8.309569032794694e-11
+   -2.067131551637735e-11
+    8.458245614594078e-11
+   -7.457065666919324e-13
+   -9.826798566527944e-12
+    8.460788400920794e-11
+   -2.235957987841259e-13
+   -7.428413854976882e-13
+   -2.067513778988974e-11
+    8.295822430824051e-11
+ 5.8e+09     
+    8.308487319028226e-11
+   -2.066624225091893e-11
+    8.457086966524679e-11
+   -7.449627921724789e-13
+   -9.823671517092105e-12
+    8.459629365512347e-11
+   -2.230681590014779e-13
+   -7.421030384588567e-13
+   -2.067007445151071e-11
+      8.2947436350399e-11
+ 5.9e+09     
+    8.307428155189982e-11
+   -2.066127441268534e-11
+    8.455952019832548e-11
+   -7.442335753433323e-13
+    -9.82057200488514e-12
+    8.458493965572112e-11
+   -2.225986637585083e-13
+   -7.413785957808529e-13
+   -2.066511471793455e-11
+     8.29368713892125e-11
+ 6e+09       
+     8.30639021079221e-11
+   -2.065640927006667e-11
+    8.454839548453854e-11
+   -7.435196076255713e-13
+   -9.817504962122929e-12
+    8.457380977027119e-11
+    -2.22188555099615e-13
+   -7.406687114598608e-13
+   -2.066025588325886e-11
+    8.292651627810421e-11
+ 6.1e+09     
+    8.305372251488596e-11
+   -2.065164431602547e-11
+    8.453748437433438e-11
+   -7.428215819730112e-13
+   -9.814476333465621e-12
+    8.456289287094941e-11
+    -2.21839142037398e-13
+   -7.399740437690363e-13
+   -2.065549547239035e-11
+    8.291635882813305e-11
+ 6.2e+09     
+    8.304373132699277e-11
+   -2.064697725663567e-11
+    8.452677674121946e-11
+   -7.421402154738556e-13
+   -9.811492915520345e-12
+    8.455217885473729e-11
+   -2.215517933090998e-13
+     -7.3929527807655e-13
+   -2.065083122962645e-11
+    8.290638774419067e-11
+ 6.3e+09     
+    8.303391793705023e-11
+   -2.064240600044267e-11
+    8.451626338988916e-11
+   -7.414762801799254e-13
+   -9.808562145179838e-12
+     8.45416585514996e-11
+   -2.213279289154051e-13
+   -7.386331579098831e-13
+   -2.064626110807001e-11
+    8.289659256595644e-11
+ 6.4e+09     
+    8.302427252180642e-11
+   -2.063792864860372e-11
+    8.450593596147945e-11
+    -7.40830640959647e-13
+    -9.80569184438404e-12
+    8.453132362919377e-11
+   -2.211690106367023e-13
+   -7.379885230625792e-13
+   -2.064178325983118e-11
+    8.288696361329831e-11
+ 6.5e+09     
+     8.30147859913543e-11
+   -2.063354348574402e-11
+    8.449578683763708e-11
+   -7.402042984660215e-13
+   -9.802889933551992e-12
+    8.452116649790751e-11
+   -2.210765318307917e-13
+   -7.373623528349138e-13
+   -2.063739602694423e-11
+    8.287749193578777e-11
+ 6.6e+09     
+    8.300544994227763e-11
+   -2.062924897144222e-11
+    8.448580904570703e-11
+   -7.395984347377455e-13
+   -9.800164129726576e-12
+    8.451118021501961e-11
+   -2.210520069043559e-13
+   -7.367558119266803e-13
+   -2.063309793290767e-11
+     8.28681692659867e-11
+ 6.7e+09     
+    8.299625661420202e-11
+   -2.062504373224702e-11
+    8.447599616771298e-11
+   -7.390144586036288e-13
+   -9.797521647787353e-12
+    8.450135839415725e-11
+   -2.210969609038778e-13
+   -7.361702961524465e-13
+   -2.062888767474411e-11
+     8.28589879761659e-11
+ 6.8e+09     
+    8.298719884942497e-11
+   -2.062092655412128e-11
+    8.446634225587342e-11
+   -7.384540480031781e-13
+   -9.794968923488711e-12
+     8.44916951206888e-11
+   -2.212129196794569e-13
+   -7.356074750921374e-13
+   -2.062476411547046e-11
+    8.284994103811851e-11
+ 6.9e+09     
+    8.297827005532058e-11
+   -2.061689637521573e-11
+    8.445684175714736e-11
+   -7.379191865893014e-13
+   -9.792511375438406e-12
+     8.44821848762456e-11
+   -2.214014010342915e-13
+   -7.350693290427601e-13
+   -2.062072627687553e-11
+    8.284102198575772e-11
+ 7e+09       
+    8.296946416923711e-11
+   -2.061295227888608e-11
+    8.444748944876119e-11
+   -7.374121925123044e-13
+   -9.790153219642842e-12
+    8.447282247422039e-11
+   -2.216639071879018e-13
+    -7.34558178170165e-13
+   -2.061677333251369e-11
+    8.283222488021256e-11
+ 7.1e+09     
+    8.296077562564993e-11
+   -2.060909348688716e-11
+    8.443828038591558e-11
+   -7.369357380218036e-13
+   -9.787897345410014e-12
+    8.446360300743907e-11
+   -2.220019187647677e-13
+   -7.340767024969229e-13
+   -2.061290460084301e-11
+    8.282354427717781e-11
+ 7.2e+09     
+    8.295219932536518e-11
+   -2.060531935269908e-11
+     8.44292098620121e-11
+   -7.364928593587344e-13
+   -9.785745255913043e-12
+    8.445452180834529e-11
+   -2.224168903883057e-13
+   -7.336279521978192e-13
+   -2.060911953845782e-11
+    8.281497519630876e-11
+ 7.3e+09     
+    8.294373060661025e-11
+   -2.060162935496313e-11
+    8.442027338090125e-11
+   -7.360869572294559e-13
+   -9.783697071329157e-12
+    8.444557442119444e-11
+   -2.229102478310335e-13
+   -7.332153484938229e-13
+   -2.060541773338808e-11
+    8.280651309249373e-11
+ 7.4e+09     
+    8.293536521788246e-11
+   -2.059802309102512e-11
+    8.441146663993183e-11
+   -7.357217888564608e-13
+   -9.781751587843696e-12
+    8.443675658503777e-11
+   -2.234833865614156e-13
+   -7.328426761380034e-13
+   -2.060179889845813e-11
+    8.279815382887154e-11
+ 7.5e+09     
+    8.292709929245543e-11
+    -2.05945002705987e-11
+    8.440278552205728e-11
+   -7.354014531153158e-13
+   -9.779906382415696e-12
+    8.442806422574638e-11
+   -2.241376714470123e-13
+     -7.3251406900141e-13
+   -2.059826286471163e-11
+    8.278989365148872e-11
+ 7.6e+09     
+      8.2918929324459e-11
+   -2.059106070957123e-11
+    8.439422609495685e-11
+    -7.35130370560537e-13
+   -9.778157951261381e-12
+    8.441949345503677e-11
+   -2.248744373278353e-13
+   -7.322339905600582e-13
+   -2.059480957492088e-11
+    8.278172916551188e-11
+ 7.7e+09     
+    8.291085214646771e-11
+   -2.058770432397944e-11
+    8.438578461506094e-11
+   -7.349132602193656e-13
+   -9.776501869499357e-12
+    8.441104057437749e-11
+   -2.256949901621265e-13
+   -7.320072111600453e-13
+   -2.059143907720128e-11
+    8.277365731292453e-11
+ 7.8e+09     
+    8.290286490853215e-11
+   -2.058443112418047e-11
+    8.437745753448779e-11
+   -7.347551149228759e-13
+   -9.774932960106893e-12
+    8.440270208179008e-11
+   -2.266006084645112e-13
+   -7.318387838281038e-13
+   -2.058815151875275e-11
+     8.27656753516427e-11
+ 7.9e+09     
+     8.28949650585932e-11
+   -2.058124120924139e-11
+    8.436924150916315e-11
+   -7.346611766999939e-13
+   -9.773445461927443e-12
+    8.439447467980651e-11
+   -2.275925447951805e-13
+   -7.317340201509525e-13
+   -2.058494713974442e-11
+    8.275778083598452e-11
+ 8e+09       
+    8.288715032421435e-11
+   -2.057813476156186e-11
+    8.436113340673153e-11
+    -7.34636913436694e-13
+   -9.772033188582923e-12
+    8.438635528319736e-11
+   -2.286720271101535e-13
+   -7.316984674228855e-13
+   -2.058182626735428e-11
+    8.274997159842957e-11
+ 8.1e+09     
+    8.287941869556513e-11
+   -2.057511204173946e-11
+    8.435313031324226e-11
+   -7.346879976511787e-13
+   -9.770689672441251e-12
+    8.437834102544563e-11
+   -2.298402598382809e-13
+   -7.317378879098036e-13
+   -2.057878930996625e-11
+     8.27422457325949e-11
+ 8.2e+09     
+    8.287176840958236e-11
+   -2.057217338367856e-11
+    8.434522953794941e-11
+   -7.348202878983681e-13
+    -9.76940828999901e-12
+    8.437042926330778e-11
+   -2.310984246042283e-13
+   -7.318582407395794e-13
+   -2.057583675152278e-11
+    8.273460157735844e-11
+ 8.3e+09     
+    8.286419793523731e-11
+   -2.056931918993821e-11
+    8.433742861587283e-11
+   -7.350398130200691e-13
+   -9.768182366977123e-12
+    8.436261757910686e-11
+   -2.324476805637957e-13
+   -7.320656666317065e-13
+   -2.057296914602248e-11
+    8.272703770204975e-11
+ 8.4e+09     
+    8.285670595982946e-11
+   -2.056654992730983e-11
+    8.432972530802703e-11
+   -7.353527592175308e-13
+   -9.767005262992649e-12
+    8.435490378066194e-11
+   -2.338891643560127e-13
+    -7.32366475438946e-13
+   -2.057018711214971e-11
+    8.271955289263225e-11
+ 8.5e+09     
+    8.284929137623391e-11
+   -2.056386612261182e-11
+     8.43221175994086e-11
+   -7.357654597442553e-13
+   -9.765870436831231e-12
+    8.434728589894471e-11
+   -2.354239897050487e-13
+   -7.327671362945123e-13
+   -2.056749132801895e-11
+    8.271214613879844e-11
+ 8.6e+09     
+    8.284195327102339e-11
+   -2.056126835868613e-11
+    8.431460369496183e-11
+    -7.36284386896502e-13
+   -9.764771494123485e-12
+     8.43397621836812e-11
+   -2.370532467243063e-13
+   -7.332742700373401e-13
+   -2.056488252601509e-11
+    8.270481662190137e-11
+ 8.7e+09     
+     8.28346909133954e-11
+   -2.055875727058249e-11
+    8.430718201381925e-11
+   -7.369161459083857e-13
+    -9.76370221967594e-12
+    8.433233109719281e-11
+    -2.38778000986679e-13
+   -7.338946435170757e-13
+   -2.056236148771102e-11
+    8.269756370364895e-11
+ 8.8e+09     
+    8.282750374483507e-11
+   -2.055633354191476e-11
+    8.429985118214368e-11
+   -7.376674703284475e-13
+   -9.762656596889196e-12
+    8.432499130680574e-11
+   -2.405992924300376e-13
+   -7.346351653497506e-13
+   -2.055992903884414e-11
+    8.269038691549028e-11
+ 8.9e+09     
+    8.282039136944703e-11
+   -2.055399790137632e-11
+    8.429261002490222e-11
+    -7.38545218453771e-13
+   -9.761628816681852e-12
+    8.431774167615475e-11
+   -2.425181341677006e-13
+   -7.355028826937526e-13
+   -2.055758604433496e-11
+     8.26832859486279e-11
+ 9e+09       
+    8.281335354489834e-11
+   -2.055175111940255e-11
+    8.428545755688054e-11
+   -7.395563704173848e-13
+   -9.760613278190592e-12
+    8.431058125569073e-11
+   -2.445355112710266e-13
+   -7.365049786349072e-13
+   -2.055533340333302e-11
+     8.26762606445954e-11
+ 9.1e+09     
+    8.280639017391434e-11
+   -2.054959400497015e-11
+    8.427839297321514e-11
+   -7.407080255562522e-13
+   -9.759604583288945e-12
+    8.430350927266945e-11
+   -2.466523795867825e-13
+   -7.376487698001375e-13
+   -2.055317204427797e-11
+    8.266931098634165e-11
+ 9.2e+09     
+    8.279950129627701e-11
+   -2.054752740252615e-11
+    8.427141563967941e-11
+   -7.420073997245918e-13
+   -9.758597526697741e-12
+    8.429652512085552e-11
+   -2.488696646465763e-13
+   -7.389417038562997e-13
+   -2.055110291996563e-11
+    8.266243708977065e-11
+ 9.3e+09     
+    8.279268708127859e-11
+   -2.054555218904038e-11
+    8.426452508291827e-11
+   -7.434618222561149e-13
+   -9.757587083183213e-12
+    8.428962835013844e-11
+   -2.511882607201816e-13
+   -7.403913565884849e-13
+   -2.054912700261259e-11
+    8.265563919568804e-11
+ 9.4e+09     
+      8.2785947820586e-11
+   -2.054366927117849e-11
+    8.425772098078905e-11
+    -7.45078732315494e-13
+   -9.756568393071056e-12
+    8.428281865621544e-11
+   -2.536090300591445e-13
+   -7.420054282886404e-13
+   -2.054724527891407e-11
+    8.264891766211066e-11
+ 9.5e+09     
+    8.277928392147759e-11
+   -2.054187958259365e-11
+    8.425100315292453e-11
+    -7.46865674413014e-13
+    -9.75553674706053e-12
+    8.427609587046008e-11
+   -2.561328023725619e-13
+   -7.437917392176244e-13
+   -2.054545874509388e-11
+    8.264227295689748e-11
+ 9.6e+09     
+    8.277269590041285e-11
+    -2.05401840813371e-11
+    8.424437155160711e-11
+   -7.488302928846911e-13
+   -9.754487571108763e-12
+    8.426945995006505e-11
+   -2.587603745728125e-13
+   -7.457582239318163e-13
+   -2.054376840194702e-11
+    8.263570565066554e-11
+ 9.7e+09     
+    8.276618437690431e-11
+   -2.053858374739031e-11
+    8.423782625301308e-11
+   -7.509803251640719e-13
+    -9.75341641197253e-12
+    8.426291096851782e-11
+   -2.614925108259813e-13
+   -7.479129242882627e-13
+    -2.05421752498778e-11
+    8.262921640995647e-11
+ 9.8e+09     
+    8.275975006765587e-11
+   -2.053707958032144e-11
+    8.423136744886365e-11
+   -7.533235936908259e-13
+   -9.752318923844321e-12
+    8.425644910644894e-11
+   -2.643299429391396e-13
+   -7.502639809603384e-13
+   -2.054068028393952e-11
+     8.26228059906204e-11
+ 9.9e+09     
+    8.275339378094116e-11
+   -2.053567259707204e-11
+    8.422499543850235e-11
+   -7.558679963156253e-13
+   -9.751190856396836e-12
+    8.425007464287346e-11
+   -2.672733711150228e-13
+   -7.528196233095554e-13
+   -2.053928448888313e-11
+    8.261647523138868e-11
+ 1e+10       
+    8.274711641119144e-11
+   -2.053436382987935e-11
+    8.421871062140328e-11
+   -7.586214950716547e-13
+   -9.750028044454334e-12
+    8.424378794683085e-11
+    -2.70323465103354e-13
+   -7.555881574687884e-13
+   -2.053798883422521e-11
+    8.261022504760704e-11
+ 1.01e+10    
+    8.274046670555712e-11
+   -2.053421894857917e-11
+    8.421057255650754e-11
+   -7.603598366570135e-13
+   -9.751573808028176e-12
+    8.423599112079564e-11
+   -2.732389437670171e-13
+   -7.573093908460148e-13
+   -2.053791467638209e-11
+    8.260361709451382e-11
+ 1.02e+10    
+    8.273386489301764e-11
+   -2.053407790984924e-11
+    8.420260598918166e-11
+   -7.621405680592108e-13
+   -9.753049521172555e-12
+    8.422834169872604e-11
+    -2.76185478942822e-13
+   -7.590736801128107e-13
+   -2.053783927675941e-11
+    8.259705557416601e-11
+ 1.03e+10    
+    8.272731123821393e-11
+   -2.053394032965235e-11
+     8.41948065268367e-11
+   -7.639627068445014e-13
+   -9.754458091283077e-12
+    8.422083658805324e-11
+   -2.791628557786777e-13
+   -7.608800039610581e-13
+    -2.05377625172344e-11
+    8.259054080471093e-11
+ 1.04e+10    
+    8.272080597481111e-11
+   -2.053380586625661e-11
+    8.418716991778352e-11
+   -7.658252959419342e-13
+   -9.755802315657977e-12
+    8.421347277036487e-11
+   -2.821708423231979e-13
+   -7.627273684668009e-13
+   -2.053768430866087e-11
+    8.258407307115293e-11
+ 1.05e+10    
+    8.271434930634816e-11
+   -2.053367421799218e-11
+    8.417969204620122e-11
+   -7.677274027937633e-13
+   -9.757084886169103e-12
+    8.420624729983936e-11
+   -2.852091902170224e-13
+   -7.646148061378244e-13
+   -2.053760458930631e-11
+     8.25776526263104e-11
+ 1.06e+10    
+     8.27079414070866e-11
+   -2.053354512109613e-11
+     8.41723689272898e-11
+   -7.696681185412689e-13
+   -9.758308393720954e-12
+    8.419915730167814e-11
+   -2.882776353709749e-13
+   -7.665413750023033e-13
+   -2.053752332334139e-11
+     8.25712796917677e-11
+ 1.07e+10    
+    8.270158242285659e-11
+   -2.053341834764374e-11
+    8.416519670260063e-11
+   -7.716465572453645e-13
+   -9.759475332506849e-12
+    8.419219997054006e-11
+   -2.913758986307197e-13
+   -7.685061577371551e-13
+   -2.053744049938164e-11
+    8.256495445881721e-11
+ 1.08e+10    
+    8.269527247189942e-11
+   -2.053329370356318e-11
+    8.415817163553649e-11
+   -7.736618551397248e-13
+   -9.760588104071106e-12
+    8.418537256897932e-11
+   -2.945036864280211e-13
+   -7.705082608338388e-13
+   -2.053735612907986e-11
+    8.255867708939331e-11
+ 1.09e+10    
+    8.268901164570542e-11
+   -2.053317102673185e-11
+    8.415129010701719e-11
+   -7.757131699155359e-13
+    -9.76164902118615e-12
+    8.417867242589324e-11
+   -2.976606914184358e-13
+   -7.725468138001284e-13
+    -2.05372702457701e-11
+    8.255244771699526e-11
+ 1.1e+10     
+    8.268280000984503e-11
+   -2.053305018515123e-11
+    8.414454861130301e-11
+    -7.77799680035848e-13
+   -9.762660311552609e-12
+     8.41720969349792e-11
+   -3.008465931054761e-13
+   -7.746209683962462e-13
+   -2.053718290316117e-11
+    8.254626644760014e-11
+ 1.11e+10    
+    8.267663760479262e-11
+   -2.053293107519796e-11
+    8.413794375197114e-11
+   -7.799205840789284e-13
+   -9.763624121330453e-12
+    8.416564355320572e-11
+   -3.040610584511368e-13
+   -7.767298979036179e-13
+   -2.053709417407927e-11
+     8.25401333605623e-11
+ 1.12e+10    
+    8.267052444674239e-11
+   -2.053281361994934e-11
+    8.413147223803909e-11
+   -7.820751001087023e-13
+   -9.764542518509273e-12
+    8.415930979929874e-11
+    -3.07303742472859e-13
+    -7.78872796424743e-13
+   -2.053700414925936e-11
+    8.253404850950191e-11
+ 1.13e+10    
+    8.266446052841456e-11
+   -2.053269776758046e-11
+    8.412513088023132e-11
+   -7.842624650710928e-13
+   -9.765417496124801e-12
+    8.415309325224564e-11
+   -3.105742888269529e-13
+   -7.810488782127668e-13
+   -2.053691293618374e-11
+    8.252801192317908e-11
+ 1.14e+10    
+    8.265844581985179e-11
+   -2.053258348983041e-11
+    8.411891658738095e-11
+   -7.864819342154261e-13
+   -9.766250975328903e-12
+    8.414699154981826e-11
+   -3.138723303784533e-13
+   -7.832573770292235e-13
+   -2.053682065796702e-11
+    8.252202360635413e-11
+ 1.15e+10    
+    8.265248026920431e-11
+   -2.053247078053586e-11
+     8.41128263629652e-11
+   -7.887327805393946e-13
+   -9.767044808319998e-12
+    8.414100238711646e-11
+   -3.171974897574532e-13
+   -7.854975455288519e-13
+   -2.053672745228657e-11
+    8.251608354063417e-11
+ 1.16e+10    
+     8.26465638035042e-11
+   -2.053235965422952e-11
+    8.410685730176722e-11
+   -7.910142942563536e-13
+   -9.767800781140419e-12
+    8.413512351513425e-11
+   -3.205493799021162e-13
+   -7.877686546697875e-13
+   -2.053663347035739e-11
+    8.251019168530445e-11
+ 1.17e+10    
+    8.264069632942684e-11
+   -2.053225014480128e-11
+    8.410100658666137e-11
+   -7.933257822843026e-13
+    -9.76852061634698e-12
+    8.412935273934892e-11
+   -3.239276045882505e-13
+   -7.900699931482342e-13
+   -2.053653887595015e-11
+    8.250434797814389e-11
+ 1.18e+10    
+     8.26348777340403e-11
+   -2.053214230421973e-11
+    8.409527148551593e-11
+   -7.956665677552388e-13
+   -9.769205975560732e-12
+    8.412368791833401e-11
+   -3.273317589456234e-13
+   -7.924008668563772e-13
+   -2.053644384445139e-11
+    8.249855233622599e-11
+ 1.19e+10    
+    8.262910788554097e-11
+   -2.053203620131222e-11
+    8.408964934821117e-11
+   -7.980359895439492e-13
+   -9.769858461901728e-12
+    8.411812696239853e-11
+   -3.307614299611372e-13
+   -7.947605983623195e-13
+   -2.053634856196498e-11
+     8.24928046567031e-11
+ 1.2e+10     
+     8.26233866339764e-11
+   -2.053193192060145e-11
+    8.408413760376653e-11
+   -8.004334018151924e-13
+   -9.770479622314327e-12
+    8.411266783225013e-11
+   -3.342161969689798e-13
+    -7.97148526410812e-13
+   -2.053625322445308e-11
+    8.248710481757496e-11
+ 1.21e+10    
+    8.261771381195385e-11
+   -2.053182956119605e-11
+    8.407873375757431e-11
+   -8.028581735886347e-13
+   -9.771070949788001e-12
+    8.410730853768614e-11
+   -3.376956321277596e-13
+    -7.99564005444367e-13
+   -2.053615803691624e-11
+    8.248145267844061e-11
+ 1.22e+10    
+    8.261208923533435e-11
+   -2.053172923573377e-11
+    8.407343538873548e-11
+   -8.053096883207753e-13
+   -9.771633885478882e-12
+    8.410204713631065e-11
+   -3.411993008848365e-13
+   -8.020064051430319e-13
+    -2.05360632126108e-11
+    8.247584808123375e-11
+ 1.23e+10    
+    8.260651270391292e-11
+   -2.053163106937491e-11
+    8.406824014749391e-11
+   -8.077873435021923e-13
+   -9.772169820736858e-12
+    8.409688173227848e-11
+   -3.447267624281106e-13
+   -8.044751099822337e-13
+   -2.053596897230294e-11
+    8.247029085094205e-11
+ 1.24e+10    
+    8.260098400208371e-11
+   -2.053153519884443e-11
+    8.406314575276546e-11
+   -8.102905502708543e-13
+   -9.772680099042416e-12
+    8.409181047506706e-11
+   -3.482775701250444e-13
+   -8.069695188080263e-13
+   -2.053587554355801e-11
+     8.24647807963089e-11
+ 1.25e+10    
+    8.259550289949063e-11
+   -2.053144177152071e-11
+    8.405814998975942e-11
+   -8.128187330390544e-13
+   -9.773166017857845e-12
+    8.408683155827484e-11
+   -3.518512719495244e-13
+   -8.094890444286005e-13
+   -2.053578316006379e-11
+    8.245931771051923e-11
+ 1.26e+10    
+      8.2590069151663e-11
+   -2.053135094456919e-11
+    8.405325070768659e-11
+   -8.153713291349354e-13
+   -9.773628830396802e-12
+    8.408194321844784e-11
+    -3.55447410896303e-13
+   -8.120331132212978e-13
+   -2.053569206098705e-11
+    8.245390137186798e-11
+ 1.27e+10    
+     8.25846825006357e-11
+   -2.053126288411911e-11
+    8.404844581755357e-11
+   -8.179477884563322e-13
+   -9.774069747316196e-12
+    8.407714373393385e-11
+   -3.590655253835331e-13
+   -8.146011647544806e-13
+   -2.053560249036201e-11
+    8.244853154441215e-11
+ 1.28e+10    
+    8.257934267555514e-11
+   -2.053117776448202e-11
+    8.404373329003831e-11
+   -8.205475731377487e-13
+   -9.774489938333938e-12
+    8.407243142376307e-11
+   -3.627051496432652e-13
+   -8.171926514235992e-13
+   -2.053551469650938e-11
+    8.244320797860654e-11
+ 1.29e+10    
+    8.257404939326972e-11
+   -2.053109576740958e-11
+    8.403911115344404e-11
+   -8.231701572288939e-13
+   -9.774890533776317e-12
+    8.406780464655677e-11
+   -3.663658141003235e-13
+   -8.198070381003937e-13
+   -2.053542893148524e-11
+     8.24379304119217e-11
+ 1.3e+10     
+    8.256880235890445e-11
+   -2.053101708139006e-11
+    8.403457749172973e-11
+   -8.258150263845089e-13
+   -9.775272626058246e-12
+    8.406326179946249e-11
+   -3.700470457395491e-13
+   -8.224438017952016e-13
+    -2.05353454505587e-11
+    8.243269856944738e-11
+ 1.31e+10    
+    8.256360126642265e-11
+    -2.05309419009814e-11
+    8.403013044261326e-11
+   -8.284816775652701e-13
+    -9.77563727109963e-12
+    8.405880131711673e-11
+   -3.737483684616824e-13
+    -8.25102431331232e-13
+   -2.053526451171693e-11
+    8.242751216447702e-11
+ 1.32e+10    
+    8.255844579917028e-11
+   -2.053087042617924e-11
+    8.402576819574452e-11
+   -8.311696187486925e-13
+   -9.775985489680754e-12
+    8.405442167063283e-11
+    -3.77469303428083e-13
+   -8.277824270304228e-13
+   -2.053518637519689e-11
+    8.242237089907898e-11
+ 1.33e+10    
+     8.25533356304068e-11
+   -2.053080286181874e-11
+     8.40214889909466e-11
+   -8.338783686498946e-13
+   -9.776318268739735e-12
+    8.405012136661621e-11
+   -3.812093693943976e-13
+   -8.304833004105161e-13
+   -2.053511130304247e-11
+    8.241727446464899e-11
+ 1.34e+10    
+    8.254827042382148e-11
+   -2.053073941700916e-11
+    8.401729111652248e-11
+   -8.366074564518203e-13
+    -9.77663656261489e-12
+    8.404589894620497e-11
+   -3.849680830334492e-13
+   -8.332045738922826e-13
+    -2.05350395586864e-11
+     8.24122225424486e-11
+ 1.35e+10    
+    8.254324983403419e-11
+   -2.053068030459845e-11
+    8.401317290762333e-11
+   -8.393564215443048e-13
+   -9.776941294234185e-12
+    8.404175298413566e-11
+   -3.887449592474384e-13
+   -8.359457805171795e-13
+   -2.053497140655555e-11
+    8.240721480412728e-11
+ 1.36e+10    
+     8.25382735070822e-11
+   -2.053062574066835e-11
+    8.400913274467784e-11
+   -8.421248132714692e-13
+   -9.777233356254867e-12
+    8.403768208783431e-11
+   -3.925395114697847e-13
+   -8.387064636742333e-13
+   -2.053490711169904e-11
+    8.240225091222888e-11
+ 1.37e+10    
+    8.253334108089293e-11
+   -2.053057594405726e-11
+    8.400516905187964e-11
+   -8.449121906875497e-13
+   -9.777513612154917e-12
+    8.403368489653187e-11
+   -3.963512519566426e-13
+   -8.414861768362626e-13
+   -2.053484693943796e-11
+    8.239733052068343e-11
+ 1.38e+10    
+     8.25284521857422e-11
+   -2.053053113591064e-11
+    8.400128029573011e-11
+   -8.477181223201785e-13
+   -9.777782897279424e-12
+    8.402976008040371e-11
+   -4.001796920684193e-13
+   -8.442844833045388e-13
+   -2.053479115503596e-11
+    8.239245327528306e-11
+ 1.39e+10    
+    8.252360644469866e-11
+    -2.05304915392569e-11
+    8.399746498363569e-11
+   -8.505421859411667e-13
+   -9.778042019843118e-12
+    8.402590633973318e-11
+   -4.040243425414128e-13
+   -8.471009559620703e-13
+   -2.053474002338999e-11
+    8.238761881414445e-11
+ 1.4e+10     
+    8.251880347405469e-11
+   -2.053045737860833e-11
+    8.399372166255563e-11
+   -8.533839683443662e-13
+   -9.778291761891736e-12
+    8.402212240409747e-11
+   -4.078847137497976e-13
+   -8.499351770344671e-13
+   -2.053469380873977e-11
+    8.238282676815498e-11
+ 1.41e+10    
+    8.251404288374341e-11
+   -2.053042887958577e-11
+    8.399004891770069e-11
+   -8.562430651302003e-13
+   -9.778532880223896e-12
+      8.4018407031577e-11
+   -4.117603159581585e-13
+   -8.527867378585226e-13
+   -2.053465277439614e-11
+     8.23780767614069e-11
+ 1.42e+10    
+    8.250932427774259e-11
+    -2.05304062685655e-11
+    8.398644537127926e-11
+   -8.591190804966824e-13
+   -9.778766107275231e-12
+     8.40147590079865e-11
+   -4.156506595647199e-13
+   -8.556552386580539e-13
+   -2.053461718248628e-11
+    8.237336841161506e-11
+ 1.43e+10    
+    8.250464725446637e-11
+   -2.053038977234829e-11
+    8.398290968128901e-11
+   -8.620116270366223e-13
+   -9.778992151966702e-12
+    8.401117714612782e-11
+   -4.195552553355678e-13
+   -8.585402883264798e-13
+   -2.053458729371637e-11
+    8.236870133052328e-11
+ 1.44e+10    
+    8.250001140714234e-11
+   -2.053037961784837e-11
+    8.397944054035324e-11
+   -8.649203255406237e-13
+   -9.779211700518564e-12
+     8.40076602850636e-11
+   -4.234736146299253e-13
+   -8.614415042162021e-13
+   -2.053456336714949e-11
+     8.23640751242951e-11
+ 1.45e+10    
+     8.24954163241775e-11
+   -2.053037603180247e-11
+    8.397603667459999e-11
+   -8.678448048059089e-13
+   -9.779425417231759e-12
+    8.400420728941297e-11
+   -4.274052496167915e-13
+   -8.643585119341303e-13
+   -2.053454565999964e-11
+    8.235948939389336e-11
+ 1.46e+10    
+     8.24908615895117e-11
+   -2.053037924049752e-11
+    8.397269684258132e-11
+   -8.707847014503113e-13
+   -9.779633945237953e-12
+    8.400081704866506e-11
+   -4.313496734831125e-13
+   -8.672909451431942e-13
+   -2.053453442743952e-11
+      8.2354943735445e-11
+ 1.47e+10    
+     8.24863467829585e-11
+   -2.053038946951606e-11
+     8.39694198342326e-11
+    -8.73739659731622e-13
+   -9.779837907219887e-12
+     8.39974884765146e-11
+   -4.353064006335813e-13
+   -8.702384453699616e-13
+   -2.053452992242294e-11
+    8.235043774059502e-11
+ 1.48e+10    
+    8.248187148053452e-11
+   -2.053040694349853e-11
+    8.396620446986917e-11
+   -8.767093313719501e-13
+   -9.780037906103239e-12
+    8.399422051021467e-11
+   -4.392749468824243e-13
+   -8.732006618173035e-13
+   -2.053453239551997e-11
+    8.234597099684703e-11
+ 1.49e+10    
+    8.247743525477745e-11
+   -2.053043188592225e-11
+    8.396304959922033e-11
+   -8.796933753864452e-13
+   -9.780234525721451e-12
+    8.399101210994951e-11
+   -4.432548296372699e-13
+   -8.761772511827442e-13
+   -2.053454209476503e-11
+     8.23415430878919e-11
+ 1.5e+10     
+    8.247303767505243e-11
+   -2.053046451889508e-11
+    8.395995410049647e-11
+    -8.82691457917251e-13
+   -9.780428331454303e-12
+    8.398786225822476e-11
+   -4.472455680751929e-13
+   -8.791678774817592e-13
+    -2.05345592655169e-11
+    8.233715359392481e-11
+ 1.51e+10    
+    8.246867830784739e-11
+   -2.053050506296429e-11
+    8.395691687949185e-11
+   -8.857032520712001e-13
+   -9.780619870842098e-12
+    8.398476995927581e-11
+   -4.512466833113638e-13
+   -8.821722118758904e-13
+   -2.053458415033019e-11
+    8.233280209195129e-11
+ 1.52e+10    
+    8.246435671705786e-11
+   -2.053055373693905e-11
+    8.395393686871887e-11
+   -8.887284377620442e-13
+   -9.780809674175878e-12
+    8.398173423849284e-11
+   -4.552576985602814e-13
+   -8.851899325056357e-13
+   -2.053461698883779e-11
+    8.232848815608099e-11
+ 1.53e+10    
+    8.246007246426112e-11
+    -2.05306107577262e-11
+    8.395101302657247e-11
+   -8.917667015568017e-13
+   -9.780998255064995e-12
+    8.397875414186269e-11
+    -4.59278139289807e-13
+   -8.882207243278346e-13
+   -2.053465801764337e-11
+    8.232421135781163e-11
+ 1.54e+10    
+    8.245582510898008e-11
+   -2.053067634017866e-11
+    8.394814433652637e-11
+   -8.948177365256848e-13
+   -9.781186110983319e-12
+    8.397582873542754e-11
+   -4.633075333683448e-13
+    -8.91264278957149e-13
+   -2.053470747022428e-11
+     8.23199712663018e-11
+ 1.55e+10    
+    8.245161420893734e-11
+   -2.053075069695582e-11
+    8.394532980635668e-11
+   -8.978812420961128e-13
+   -9.781373723794437e-12
+    8.397295710475912e-11
+   -4.673454112050387e-13
+   -8.943202945120642e-13
+   -2.053476557684317e-11
+    8.231576744863324e-11
+ 1.56e+10    
+    8.244743932029882e-11
+   -2.053083403839497e-11
+    8.394256846739376e-11
+   -9.009569239100483e-13
+    -9.78156156025722e-12
+    8.397013835444733e-11
+    -4.71391305883516e-13
+   -8.973884754645839e-13
+   -2.053483256446883e-11
+    8.231159947006393e-11
+ 1.57e+10    
+    8.244329999790923e-11
+   -2.053092657239386e-11
+    8.393985937379991e-11
+   -9.040444936850694e-13
+   -9.781750072512399e-12
+    8.396737160760557e-11
+   -4.754447532890786e-13
+   -9.004685324937488e-13
+   -2.053490865670545e-11
+    8.230746689427007e-11
+ 1.58e+10    
+    8.243919579551691e-11
+   -2.053102850430317e-11
+    8.393720160187409e-11
+   -9.071436690785195e-13
+   -9.781939698551107e-12
+    8.396465600538863e-11
+   -4.795052922296472e-13
+   -9.035601823431579e-13
+   -2.053499407372944e-11
+    8.230336928357955e-11
+ 1.59e+10    
+    8.243512626599061e-11
+   -2.053114003682869e-11
+    8.393459424937928e-11
+   -9.102541735550815e-13
+   -9.782130862665919e-12
+    8.396199070652617e-11
+   -4.835724645506283e-13
+   -9.066631476816463e-13
+   -2.053508903223431e-11
+    8.229930619919591e-11
+ 1.6e+10     
+    8.243109096152695e-11
+   -2.053126136994274e-11
+    8.393203643489525e-11
+   -9.133757362574492e-13
+   -9.782323975885526e-12
+    8.395937488686907e-11
+   -4.876458152437759e-13
+   -9.097771569676914e-13
+   -2.053519374538235e-11
+    8.229527720141307e-11
+ 1.61e+10    
+    8.242708943384999e-11
+   -2.053139270080414e-11
+    8.392952729719342e-11
+   -9.165080918798373e-13
+   -9.782519436393313e-12
+    8.395680773894896e-11
+   -4.917248925503637e-13
+   -9.129019443169735e-13
+   -2.053530842276311e-11
+    8.229128184982153e-11
+ 1.62e+10    
+    8.242312123440193e-11
+   -2.053153422368634e-11
+    8.392706599463268e-11
+   -9.196509805446363e-13
+   -9.782717629930738e-12
+    8.395428847155086e-11
+    -4.95809248058702e-13
+    -9.16037249373154e-13
+   -2.053543327035814e-11
+    8.228731970350627e-11
+ 1.63e+10    
+    8.241918591452621e-11
+   -2.053168612991345e-11
+    8.392465170457784e-11
+   -9.228041476816483e-13
+     -9.7829189301863e-12
+    8.395181630929827e-11
+   -4.998984367961929e-13
+   -9.191828171818111e-13
+     -2.0535568490512e-11
+    8.228339032123543e-11
+ 1.64e+10    
+    8.241528302564284e-11
+   -2.053184860780342e-11
+     8.39222836228373e-11
+   -9.259673439102859e-13
+   -9.783123699170386e-12
+    8.394939049225017e-11
+   -5.039920173161388e-13
+   -9.223383980671941e-13
+   -2.053571428190868e-11
+    8.227949326164249e-11
+ 1.65e+10    
+    8.241141211941576e-11
+   -2.053202184261811e-11
+    8.391996096312034e-11
+   -9.291403249241266e-13
+   -9.783332287576731e-12
+    8.394701027550976e-11
+   -5.080895517793901e-13
+   -9.255037475119946e-13
+   -2.053587083955337e-11
+    8.227562808339952e-11
+ 1.66e+10    
+    8.240757274791325e-11
+   -2.053220601652003e-11
+    8.391768295651307e-11
+   -9.323228513782186e-13
+   -9.783545035131098e-12
+    8.394467492884464e-11
+    -5.12190606031014e-13
+   -9.286786260398424e-13
+   -2.053603835475952e-11
+    8.227179434538358e-11
+ 1.67e+10    
+    8.240376446376129e-11
+   -2.053240130853508e-11
+    8.391544885097263e-11
+    -9.35514688778793e-13
+   -9.783762270927632e-12
+    8.394238373631805e-11
+   -5.162947496721097e-13
+    -9.31862799100509e-13
+   -2.053621701514015e-11
+    8.226799160683505e-11
+ 1.68e+10    
+    8.239998682029008e-11
+   -2.053260789452118e-11
+    8.391325791083865e-11
+   -9.387156073753331e-13
+    -9.78398431375345e-12
+    8.394013599593042e-11
+   -5.204015561269916e-13
+   -9.350560369576642e-13
+   -2.053640700460406e-11
+    8.226421942751003e-11
+ 1.69e+10    
+    8.239623937167319e-11
+   -2.053282594714226e-11
+    8.391110941636101e-11
+   -9.419253820550161e-13
+    -9.78421147240179e-12
+    8.393793101927169e-11
+   -5.245106027057593e-13
+   -9.382581145792398e-13
+   -2.053660850335591e-11
+    8.226047736782467e-11
+ 1.7e+10     
+    8.239252167306111e-11
+   -2.053305563584735e-11
+    8.390900266324411e-11
+   -9.451437922393102e-13
+   -9.784444045974518e-12
+    8.393576813118351e-11
+   -5.286214706625419e-13
+   -9.414688115301379e-13
+   -2.053682168790036e-11
+    8.225676498899406e-11
+ 1.71e+10    
+    8.238883328070846e-11
+   -2.053329712685475e-11
+    8.390693696220649e-11
+   -9.483706217829121e-13
+   -9.784682324173954e-12
+    8.393364666943094e-11
+   -5.327337452494141e-13
+   -9.446879118674188e-13
+    -2.05370467310497e-11
+    8.225308185316377e-11
+ 1.72e+10    
+    8.238517375209434e-11
+   -2.053355058314027e-11
+    8.390491163855446e-11
+   -9.516056588747385e-13
+   -9.784926587584864e-12
+    8.393156598438402e-11
+   -5.368470157662035e-13
+   -9.479152040376832e-13
+   -2.053728380193503e-11
+    8.224942752353522e-11
+ 1.73e+10    
+    8.238154264603783e-11
+   -2.053381616443021e-11
+    8.390292603177158e-11
+   -9.548486959408361e-13
+    -9.78517710794682e-12
+    8.392952543870759e-11
+   -5.409608756063522e-13
+    -9.51150480776809e-13
+   -2.053753306602063e-11
+    8.224580156448645e-11
+ 1.74e+10    
+    8.237793952280734e-11
+   -2.053409402719789e-11
+    8.390097949512059e-11
+   -9.580995295495883e-13
+   -9.785434148417268e-12
+    8.392752440706129e-11
+   -5.450749222988391e-13
+   -9.543935390117258e-13
+    -2.05377946851212e-11
+    8.224220354168476e-11
+ 1.75e+10    
+    8.237436394422421e-11
+   -2.053438432466421e-11
+    8.389907139525871e-11
+   -9.613579603186899e-13
+   -9.785697963825785e-12
+    8.392556227580656e-11
+    -5.49188757546416e-13
+   -9.576441797643636e-13
+   -2.053806881742191e-11
+    8.223863302219558e-11
+ 1.76e+10    
+    8.237081547376176e-11
+   -2.053468720680159e-11
+    8.389720111186642e-11
+    -9.64623792823945e-13
+   -9.785968800919844e-12
+    8.392363844272339e-11
+   -5.533019872602334e-13
+   -9.609022080577137e-13
+   -2.053835561750112e-11
+     8.22350895745856e-11
+ 1.77e+10    
+    8.236729367663897e-11
+   -2.053500282034113e-11
+    8.389536803728772e-11
+   -9.678968355102281e-13
+   -9.786246898602279e-12
+    8.392175231673393e-11
+     -5.5741422159094e-13
+   -9.641674328237407e-13
+   -2.053865523635525e-11
+    8.223157276901966e-11
+ 1.78e+10    
+    8.236379811990801e-11
+   -2.053533130878275e-11
+    8.389357157618254e-11
+   -9.711769006038694e-13
+    -9.78653248816104e-12
+    8.391990331763451e-11
+   -5.615250749564651e-13
+   -9.674396668133383e-13
+   -2.053896782142619e-11
+    8.222808217735382e-11
+ 1.79e+10    
+     8.23603283725394e-11
+   -2.053567281240848e-11
+    8.389181114519072e-11
+    -9.74463804027147e-13
+    -9.78682579349134e-12
+    8.391809087583534e-11
+   -5.656341660664972e-13
+   -9.707187265081651e-13
+   -2.053929351663054e-11
+    8.222461737322323e-11
+ 1.8e+10     
+    8.235688400550039e-11
+   -2.053602746829793e-11
+    8.389008617260627e-11
+   -9.777573653142338e-13
+    -9.78712703131036e-12
+    8.391631443210659e-11
+   -5.697411179438599e-13
+   -9.740044320342943e-13
+   -2.053963246239047e-11
+      8.2221177932124e-11
+ 1.81e+10    
+    8.235346459182969e-11
+   -2.053639541034645e-11
+    8.388839609806274e-11
+   -9.810574075290316e-13
+   -9.787436411365186e-12
+    8.391457343733284e-11
+    -5.73845557942842e-13
+   -9.772966070776497e-13
+   -2.053998479566712e-11
+    8.221776343149322e-11
+ 1.82e+10    
+    8.235006970670859e-11
+   -2.053677676928566e-11
+     8.38867403722286e-11
+   -9.843637571844536e-13
+   -9.787754136633973e-12
+    8.391286735227364e-11
+   -5.779471177646301e-13
+   -9.805950788012025e-13
+   -2.054035064999455e-11
+    8.221437345078149e-11
+ 1.83e+10    
+    8.234669892752663e-11
+   -2.053717167270593e-11
+    8.388511845651239e-11
+   -9.876762441634626e-13
+   -9.788080403520449e-12
+    8.391119564732996e-11
+   -5.820454334698964e-13
+   -9.838996777639278e-13
+   -2.054073015551597e-11
+    8.221100757152359e-11
+ 1.84e+10    
+    8.234335183394431e-11
+   -2.053758024508063e-11
+    8.388352982277732e-11
+   -9.909947016415552e-13
+   -9.788415402042444e-12
+    8.390955780231929e-11
+   -5.861401454887164e-13
+   -9.872102378412713e-13
+   -2.054112343902086e-11
+    8.220766537740372e-11
+ 1.85e+10    
+    8.234002800795162e-11
+   -2.053800260779266e-11
+    8.388197395306466e-11
+   -9.943189660108903e-13
+   -9.788759316014172e-12
+    8.390795330625433e-11
+   -5.902308986278382e-13
+   -9.905265961475136e-13
+   -2.054153062398337e-11
+    8.220434645431786e-11
+ 1.86e+10    
+    8.233672703392254e-11
+     -2.0538438879162e-11
+    8.388045033932641e-11
+   -9.976488768058704e-13
+   -9.789112323222936e-12
+    8.390638165712968e-11
+   -5.943173420754741e-13
+   -9.938485929593386e-13
+   -2.054195183060187e-11
+    8.220105039043084e-11
+ 1.87e+10    
+    8.233344849866662e-11
+   -2.053888917447538e-11
+    8.387895848316561e-11
+   -1.000984276630021e-12
+   -9.789474595600119e-12
+    8.390484236171327e-11
+   -5.983991294037014e-13
+   -9.971760716413153e-13
+   -2.054238717583935e-11
+    8.219777677623164e-11
+ 1.88e+10    
+    8.233019199147671e-11
+   -2.053935360601681e-11
+      8.3877497895586e-11
+   -1.004325011084605e-12
+   -9.789846299386931e-12
+    8.390333493534444e-11
+   -6.024759185684592e-13
+   -1.000508878572696e-12
+   -2.054283677346484e-11
+    8.219452520458342e-11
+ 1.89e+10    
+    8.232695710417378e-11
+   -2.053983228309975e-11
+    8.387606809674802e-11
+   -1.007670928698412e-12
+   -9.790227595294846e-12
+    8.390185890173619e-11
+    -6.06547371907423e-13
+   -1.003846863075742e-12
+   -2.054330073409541e-11
+    8.219129527077164e-11
+ 1.9e+10     
+    8.232374343114744e-11
+   -2.054032531210009e-11
+    8.387466861573356e-11
+   -1.011021880858968e-12
+   -9.790618638661188e-12
+    8.390041379278392e-11
+   -6.106131561356699e-13
+   -1.007189877345465e-12
+   -2.054377916523903e-11
+    8.218808657254766e-11
+ 1.91e+10    
+    8.232055056939532e-11
+   -2.054083279649051e-11
+    8.387329899031732e-11
+   -1.014377721745143e-12
+   -9.791019579599884e-12
+    8.389899914837904e-11
+   -6.146729423393374e-13
+   -1.010537776380846e-12
+    -2.05442721713378e-11
+    8.218489871017014e-11
+ 1.92e+10    
+    8.231737811855742e-11
+   -2.054135483687537e-11
+    8.387195876674533e-11
+   -1.017738308261018e-12
+   -9.791430563147467e-12
+     8.38976145162271e-11
+   -6.187264059672531e-13
+   -1.013890417917426e-12
+   -2.054477985381197e-11
+    8.218173128644311e-11
+ 1.93e+10    
+    8.231422568094956e-11
+   -2.054189153102684e-11
+    8.387064749952085e-11
+   -1.021103499971067e-12
+   -9.791851729404853e-12
+    8.389625945167114e-11
+   -6.227732268207733e-13
+   -1.017247662361192e-12
+   -2.054530231110394e-11
+    8.217858390675078e-11
+ 1.94e+10    
+    8.231109286159246e-11
+   -2.054244297392134e-11
+    8.386936475119526e-11
+   -1.024473159036595e-12
+   -9.792283213674543e-12
+    8.389493351751983e-11
+   -6.268130890417402e-13
+   -1.020609372723826e-12
+   -2.054583963872316e-11
+    8.217545617909031e-11
+ 1.95e+10    
+    8.230797926823927e-11
+   -2.054300925777702e-11
+      8.3868110092167e-11
+   -1.027847150153385e-12
+     -9.7927251465939e-12
+    8.389363628388014e-11
+    -6.30845681098748e-13
+   -1.023975414559298e-12
+   -2.054639192929088e-11
+    8.217234771410142e-11
+ 1.96e+10    
+    8.230488451140045e-11
+    -2.05435904720916e-11
+    8.386688310048584e-11
+   -1.031225340490666e-12
+   -9.793177654264266e-12
+    8.389236732799422e-11
+   -6.348706957717394e-13
+   -1.027345655901684e-12
+   -2.054695927258532e-11
+    8.216925812509338e-11
+ 1.97e+10    
+    8.230180820436601e-11
+   -2.054418670368064e-11
+    8.386568336166267e-11
+   -1.034607599631129e-12
+   -9.793640858376261e-12
+    8.389112623408026e-11
+   -6.388878301350481e-13
+   -1.030719967204241e-12
+   -2.054754175558675e-11
+    8.216618702806969e-11
+ 1.98e+10    
+    8.229874996322505e-11
+   -2.054479803671635e-11
+     8.38645104684852e-11
+    -1.03799379951219e-12
+   -9.794114876331346e-12
+    8.388991259317861e-11
+    -6.42896785538938e-13
+    -1.03409822127966e-12
+   -2.054813946252307e-11
+    8.216313404175064e-11
+ 1.99e+10    
+    8.229570940688438e-11
+   -2.054542455276669e-11
+    8.386336402083937e-11
+   -1.041383814368464e-12
+   -9.794599821359784e-12
+    8.388872600300077e-11
+   -6.468972675896559e-13
+   -1.037480293241642e-12
+   -2.054875247491517e-11
+    8.216009878759327e-11
+ 2e+10       
+    8.229268615708352e-11
+   -2.054606633083478e-11
+    8.386224362553612e-11
+   -1.044777520675186e-12
+   -9.795095802635156e-12
+    8.388756606778283e-11
+    -6.50888986128202e-13
+   -1.040866060447497e-12
+   -2.054938087162212e-11
+      8.2157080889809e-11
+ 2.01e+10    
+    8.228967983840891e-11
+   -2.054672344739858e-11
+    8.386114889614256e-11
+   -1.048174797092946e-12
+   -9.795602925385369e-12
+     8.38864323981425e-11
+   -6.548716552077138e-13
+   -1.044255402442032e-12
+   -2.055002472888667e-11
+    8.215407997537977e-11
+ 2.02e+10    
+    8.228669007830517e-11
+   -2.054739597645047e-11
+    8.386007945281863e-11
+   -1.051575524413347e-12
+    -9.79612129100062e-12
+    8.388532461094002e-11
+   -6.588449930696676e-13
+   -1.047648200902434e-12
+    -2.05506841203804e-11
+    8.215109567407156e-11
+ 2.03e+10    
+    8.228371650708546e-11
+   -2.054808398953732e-11
+    8.385903492215821e-11
+   -1.054979585505828e-12
+   -9.796650997138034e-12
+    8.388424232914263e-11
+   -6.628087221188935e-13
+   -1.051044339584354e-12
+   -2.055135911724885e-11
+    8.214812761844671e-11
+ 2.04e+10    
+    8.228075875793904e-11
+   -2.054878755580038e-11
+     8.38580149370357e-11
+   -1.058386865265471e-12
+   -9.797192137823422e-12
+    8.388318518169187e-11
+   -6.667625688974377e-13
+   -1.054443704269134e-12
+   -2.055204978815617e-11
+    8.214517544387322e-11
+ 2.05e+10    
+    8.227781646693792e-11
+   -2.054950674201507e-11
+    8.385701913645507e-11
+   -1.061797250561909e-12
+   -9.797744803549957e-12
+    8.388215280337538e-11
+   -6.707062640574147e-13
+   -1.057846182711876e-12
+   -2.055275619933015e-11
+    8.214223878853395e-11
+ 2.06e+10    
+    8.227488927304172e-11
+   -2.055024161263112e-11
+    8.385604716540556e-11
+    -1.06521063018914e-12
+   -9.798309081374137e-12
+    8.388114483470086e-11
+   -6.746395423328502e-13
+   -1.061251664590812e-12
+   -2.055347841460629e-11
+    8.213931729343265e-11
+ 2.07e+10    
+    8.227197681810106e-11
+   -2.055099222981235e-11
+    8.385509867471955e-11
+   -1.068626894816407e-12
+    -9.79888505500896e-12
+    8.388016092177395e-11
+   -6.785621425105472e-13
+   -1.064660041457559e-12
+   -2.055421649547213e-11
+    8.213641060239916e-11
+ 2.08e+10    
+    8.226907874685857e-11
+   -2.055175865347628e-11
+    8.385417332093597e-11
+   -1.072045936940113e-12
+   -9.799472804914431e-12
+    8.387920071617872e-11
+   -6.824738074000648e-13
+   -1.068071206688411e-12
+   -2.055497050111105e-11
+     8.21335183620932e-11
+ 2.09e+10    
+    8.226619470694962e-11
+   -2.055254094133376e-11
+    8.385327076616619e-11
+   -1.075467650836493e-12
+   -9.800072408385509e-12
+    8.387826387486129e-11
+   -6.863742838029012e-13
+   -1.071485055436618e-12
+   -2.055574048844553e-11
+    8.213064022200569e-11
+ 2.1e+10     
+    8.226332434890167e-11
+   -2.055333914892844e-11
+    8.385239067796468e-11
+   -1.078891932515456e-12
+   -9.800683939637571e-12
+    8.387735006001604e-11
+    -6.90263322480829e-13
+   -1.074901484585682e-12
+   -2.055652651218046e-11
+    8.212777583446042e-11
+ 2.11e+10    
+    8.226046732613158e-11
+   -2.055415332967598e-11
+     8.38515327292031e-11
+   -1.082318679675207e-12
+   -9.801307469889548e-12
+    8.387645893897566e-11
+   -6.941406781235099e-13
+   -1.078320392703506e-12
+   -2.055732862484585e-11
+    8.212492485461257e-11
+ 2.12e+10    
+    8.225762329494163e-11
+   -2.055498353490277e-11
+    8.385069659794724e-11
+   -1.085747791657801e-12
+   -9.801943067444622e-12
+    8.387559018410256e-11
+   -6.980061093154143e-13
+   -1.081741679997609e-12
+   -2.055814687683894e-11
+    8.212208694044692e-11
+ 2.13e+10    
+    8.225479191451574e-11
+    -2.05558298138848e-11
+    8.384988196733803e-11
+   -1.089179169405699e-12
+   -9.802590797768731e-12
+    8.387474347268367e-11
+   -7.018593785020809e-13
+   -1.085165248271137e-12
+   -2.055898131646634e-11
+    8.211926175277519e-11
+ 2.14e+10    
+    8.225197284691248e-11
+   -2.055669221388594e-11
+    8.384908852547553e-11
+   -1.092612715418964e-12
+   -9.803250723566877e-12
+    8.387391848682767e-11
+   -7.057002519557786e-13
+   -1.088591000879903e-12
+   -2.055983198998516e-11
+    8.211644895523105e-11
+ 2.15e+10    
+    8.224916575705946e-11
+   -2.055757078019611e-11
+    8.384831596530674e-11
+   -1.096048333713603e-12
+   -9.803922904857454e-12
+    8.387311491336519e-11
+   -7.095284997405959e-13
+   -1.092018842690153e-12
+   -2.056069894164428e-11
+    8.211364821426515e-11
+ 2.16e+10    
+    8.224637031274452e-11
+   -2.055846555616891e-11
+    8.384756398451474e-11
+   -1.099485929780599e-12
+   -9.804607399044249e-12
+    8.387233244374996e-11
+   -7.133438956769981e-13
+   -1.095448680037406e-12
+   -2.056158221372451e-11
+    8.211085919913859e-11
+ 2.17e+10    
+    8.224358618460693e-11
+   -2.055937658325889e-11
+    8.384683228541294e-11
+   -1.102925410545718e-12
+   -9.805304260986776e-12
+    8.387157077396463e-11
+    -7.17146217305922e-13
+   -1.098880420685944e-12
+   -2.056248184657892e-11
+    8.210808158191554e-11
+ 2.18e+10    
+    8.224081304612825e-11
+   -2.056030390105882e-11
+     8.38461205748408e-11
+   -1.106366684330328e-12
+   -9.806013543068479e-12
+     8.38708296044264e-11
+   -7.209352458523963e-13
+   -1.102313973789333e-12
+   -2.056339787867203e-11
+    8.210531503745472e-11
+ 2.19e+10    
+    8.223805057362123e-11
+   -2.056124754733604e-11
+    8.384542856406246e-11
+   -1.109809660812866e-12
+   -9.806735295263225e-12
+    8.387010863989695e-11
+   -7.247107661887756e-13
+    -1.10574924985158e-12
+   -2.056433034661907e-11
+    8.210255924340032e-11
+ 2.2e+10     
+    8.223529844621831e-11
+   -2.056220755806883e-11
+    8.384475596866923e-11
+   -1.113254250991125e-12
+   -9.807469565199904e-12
+      8.3869407589393e-11
+   -7.284725667975906e-13
+   -1.109186160689292e-12
+   -2.056527928522416e-11
+    8.209981388017188e-11
+ 2.21e+10    
+     8.22325563458595e-11
+   -2.056318396748189e-11
+     8.38441025084826e-11
+    -1.11670036714541e-12
+   -9.808216398225288e-12
+    8.386872616610007e-11
+   -7.322204397340394e-13
+   -1.112624619394474e-12
+   -2.056624472751848e-11
+    8.209707863095307e-11
+ 2.22e+10    
+    8.222982395727998e-11
+   -2.056417680808218e-11
+     8.38434679074619e-11
+   -1.120147922802313e-12
+    -9.80897583746527e-12
+    8.386806408728748e-11
+   -7.359541805882226e-13
+   -1.116064540298226e-12
+   -2.056722670479751e-11
+    8.209435318168052e-11
+ 2.23e+10    
+    8.222710096799564e-11
+   -2.056518611069335e-11
+    8.384285189361294e-11
+    -1.12359683269939e-12
+   -9.809747923884479e-12
+    8.386742107422626e-11
+   -7.396735884470574e-13
+   -1.119505838935106e-12
+   -2.056822524665807e-11
+    8.209163722103129e-11
+ 2.24e+10    
+    8.222438706828967e-11
+   -2.056621190449056e-11
+    8.384225419889986e-11
+   -1.127047012750476e-12
+   -9.810532696344088e-12
+    8.386679685210744e-11
+   -7.433784658559476e-13
+   -1.122948432008367e-12
+   -2.056924038103434e-11
+    8.208893044040952e-11
+ 2.25e+10    
+    8.222168195119681e-11
+   -2.056725421703412e-11
+    8.384167455915869e-11
+   -1.130498380011731e-12
+   -9.811330191658436e-12
+    8.386619114996412e-11
+    -7.47068618780299e-13
+   -1.126392237355812e-12
+    -2.05702721342338e-11
+    8.208623253393303e-11
+ 2.26e+10    
+    8.221898531248884e-11
+   -2.056831307430335e-11
+    8.384111271401368e-11
+   -1.133950852648539e-12
+    -9.81214044464989e-12
+    8.386560370059416e-11
+    -7.50743856566762e-13
+   -1.129837173916482e-12
+   -2.057132053097253e-11
+     8.20835431984192e-11
+ 2.27e+10    
+    8.221629685065798e-11
+    -2.05693885007295e-11
+    8.384056840679516e-11
+   -1.137404349902838e-12
+   -9.812963488202325e-12
+    8.386503424048497e-11
+   -7.544039919043927e-13
+   -1.133283161698005e-12
+   -2.057238559440956e-11
+    8.208086213336929e-11
+ 2.28e+10    
+    8.221361626690056e-11
+   -2.057048051922829e-11
+    8.384004138446039e-11
+   -1.140858792061466e-12
+   -9.813799353313289e-12
+     8.38644825097395e-11
+   -7.580488407856456e-13
+   -1.136730121744643e-12
+   -2.057346734618118e-11
+    8.207818904095428e-11
+ 2.29e+10    
+    8.221094326510019e-11
+   -2.057158915123205e-11
+    8.383953139751528e-11
+   -1.144314100424897e-12
+   -9.814648069144645e-12
+    8.386394825200547e-11
+   -7.616782224672658e-13
+   -1.140177976106107e-12
+   -2.057456580643442e-11
+    8.207552362599786e-11
+ 2.3e+10     
+     8.22082775518102e-11
+   -2.057271441672134e-11
+    8.383903819993915e-11
+   -1.147770197276895e-12
+   -9.815509663072078e-12
+    8.386343121440416e-11
+   -7.652919594311085e-13
+   -1.143626647806925e-12
+   -2.057568099385995e-11
+     8.20728655959609e-11
+ 2.31e+10    
+     8.22056188362362e-11
+   -2.057385633425604e-11
+    8.383856154911079e-11
+   -1.151227005854588e-12
+   -9.816384160733146e-12
+    8.386293114746244e-11
+   -7.688898773449069e-13
+   -1.147076060816614e-12
+   -2.057681292572451e-11
+     8.20702146609241e-11
+ 2.32e+10    
+    8.220296683021735e-11
+   -2.057501492100598e-11
+    8.383810120573641e-11
+   -1.154684450319376e-12
+   -9.817271586074199e-12
+     8.38624478050455e-11
+    -7.72471805022981e-13
+   -1.150526140020373e-12
+    -2.05779616179027e-11
+    8.206757053357079e-11
+ 2.33e+10    
+    8.220032124820815e-11
+   -2.057619019278107e-11
+    8.383765693377977e-11
+   -1.158142455728381e-12
+   -9.818171961396097e-12
+    8.386198094429166e-11
+   -7.760375743869748e-13
+   -1.153976811190555e-12
+   -2.057912708490845e-11
+    8.206493292917008e-11
+ 2.34e+10    
+    8.219768180725967e-11
+     -2.0577382164061e-11
+    8.383722850039373e-11
+   -1.161600948006523e-12
+   -9.819085307398646e-12
+    8.386153032554773e-11
+   -7.795870204265629e-13
+   -1.157428000958675e-12
+   -2.058030933992544e-11
+    8.206230156555781e-11
+ 2.35e+10    
+    8.219504822700021e-11
+   -2.057859084802422e-11
+    8.383681567585327e-11
+    -1.16505985391927e-12
+   -9.820011643223956e-12
+    8.386109571230678e-11
+   -7.831199811602097e-13
+   -1.160879636788087e-12
+   -2.058150839483744e-11
+     8.20596761631193e-11
+ 2.36e+10    
+    8.219242022961575e-11
+   -2.057981625657676e-11
+    8.383641823349084e-11
+    -1.16851910104587e-12
+   -9.820950986498812e-12
+    8.386067687114728e-11
+   -7.866362975959817e-13
+   -1.164331646947218e-12
+   -2.058272426025801e-11
+    8.205705644477012e-11
+ 2.37e+10    
+    8.218979753983037e-11
+   -2.058105840038009e-11
+    8.383603594963247e-11
+   -1.171978617753337e-12
+   -9.821903353375709e-12
+    8.386027357167264e-11
+   -7.901358136924017e-13
+   -1.167783960483516e-12
+   -2.058395694555934e-11
+    8.205444213593763e-11
+ 2.38e+10    
+    8.218717988488647e-11
+   -2.058231728887923e-11
+    8.383566860353649e-11
+   -1.175438333170869e-12
+   -9.822868758573137e-12
+    8.385988558645293e-11
+   -7.936183763194221e-13
+    -1.17123650719782e-12
+   -2.058520645890091e-11
+    8.205183296454166e-11
+ 2.39e+10    
+     8.21845669945243e-11
+   -2.058359293032943e-11
+    8.383531597733253e-11
+   -1.178898177164925e-12
+   -9.823847215414592e-12
+     8.38595126909678e-11
+   -7.970838352194705e-13
+   -1.174689217619508e-12
+   -2.058647280725748e-11
+    8.204922866097521e-11
+ 2.4e+10     
+    8.218195860096182e-11
+   -2.058488533182311e-11
+    8.383497785596282e-11
+   -1.182358080314846e-12
+   -9.824838735866819e-12
+    8.385915466355042e-11
+   -8.005320429686388e-13
+   -1.178142022981986e-12
+   -2.058775599644641e-11
+    8.204662895808506e-11
+ 2.41e+10    
+    8.217935443887418e-11
+   -2.058619449931595e-11
+    8.383465402712482e-11
+   -1.185817973888992e-12
+   -9.825843330576965e-12
+    8.385881128533276e-11
+   -8.039628549379776e-13
+   -1.181594855198968e-12
+   -2.058905603115467e-11
+     8.20440335911519e-11
+ 2.42e+10    
+    8.217675424537273e-11
+   -2.058752043765257e-11
+      8.3834344281215e-11
+   -1.189277789821488e-12
+   -9.826861008908802e-12
+    8.385848234019184e-11
+   -8.073761292549768e-13
+   -1.185047646841122e-12
+   -2.059037291496513e-11
+    8.204144229787043e-11
+ 2.43e+10    
+     8.21741577599848e-11
+    -2.05888631505917e-11
+    8.383404841127374e-11
+   -1.192737460689415e-12
+   -9.827891778978146e-12
+    8.385816761469774e-11
+   -8.107717267651744e-13
+    -1.18850033111336e-12
+   -2.059170665038247e-11
+    8.203885481832929e-11
+ 2.44e+10    
+    8.217156472463221e-11
+   -2.059022264083098e-11
+    8.383376621293238e-11
+   -1.196196919690625e-12
+   -9.828935647687335e-12
+    8.385786689806225e-11
+   -8.141495109939717e-13
+    -1.19195284183259e-12
+   -2.059305723885843e-11
+    8.203627089499076e-11
+ 2.45e+10    
+    8.216897488361055e-11
+   -2.059159891003117e-11
+    8.383349748436072e-11
+    -1.19965610062201e-12
+   -9.829992620758807e-12
+    8.385757998208865e-11
+   -8.175093481085959e-13
+   -1.195405113406081e-12
+   -2.059442468081668e-11
+    8.203369027267077e-11
+ 2.46e+10    
+    8.216638798356786e-11
+   -2.059299195883981e-11
+      8.3833242026216e-11
+   -1.203114937858224e-12
+   -9.831062702767969e-12
+    8.385730666112254e-11
+   -8.208511068803384e-13
+   -1.198857080810194e-12
+   -2.059580897567714e-11
+    8.203111269851813e-11
+ 2.47e+10    
+    8.216380377348375e-11
+   -2.059440178691473e-11
+     8.38329996415933e-11
+   -1.206573366331043e-12
+   -9.832145897175113e-12
+    8.385704673200435e-11
+   -8.241746586469227e-13
+   -1.202308679569771e-12
+   -2.059721012187974e-11
+    8.202853792199423e-11
+ 2.48e+10    
+    8.216122200464772e-11
+   -2.059582839294663e-11
+     8.38327701359767e-11
+   -1.210031321509101e-12
+   -9.833242206356698e-12
+    8.385679999402176e-11
+   -8.274798772751465e-13
+   -1.205759845737914e-12
+   -2.059862811690759e-11
+    8.202596569485215e-11
+ 2.49e+10    
+    8.215864243063831e-11
+   -2.059727177468167e-11
+    8.383255331719217e-11
+   -1.213488739378092e-12
+   -9.834351631635803e-12
+    8.385656624886444e-11
+   -8.307666391237609e-13
+   -1.209210515876232e-12
+   -2.060006295731015e-11
+    8.202339577111642e-11
+ 2.5e+10     
+    8.215606480730143e-11
+   -2.059873192894321e-11
+    8.383234899536045e-11
+   -1.216945556421566e-12
+   -9.835474173311699e-12
+    8.385634530057832e-11
+    -8.34034823006569e-13
+    -1.21266062703569e-12
+   -2.060151463872504e-11
+    8.202082790706202e-11
+ 2.51e+10    
+    8.215348889272919e-11
+   -2.060020885165343e-11
+    8.383215698285286e-11
+   -1.220401709602015e-12
+   -9.836609830689042e-12
+    8.385613695552221e-11
+   -8.372843101558047e-13
+   -1.216110116737765e-12
+   -2.060298315590038e-11
+     8.20182618611937e-11
+ 2.52e+10    
+    8.215091444723865e-11
+   -2.060170253785428e-11
+    8.383197709424619e-11
+   -1.223857136342581e-12
+   -9.837758602105968e-12
+    8.385594102232444e-11
+   -8.405149841857587e-13
+   -1.219558922956164e-12
+   -2.060446850271581e-11
+    8.201569739422536e-11
+ 2.53e+10    
+    8.214834123335021e-11
+   -2.060321298172791e-11
+    8.383180914627952e-11
+    -1.22731177450908e-12
+   -9.838920484961844e-12
+    8.385575731184078e-11
+   -8.437267310566871e-13
+   -1.223006984098951e-12
+   -2.060597067220361e-11
+    8.201313426905915e-11
+ 2.54e+10    
+    8.214576901576644e-11
+   -2.060474017661704e-11
+    8.383165295781252e-11
+    -1.23076556239249e-12
+   -9.840095475744128e-12
+    8.385558563711292e-11
+   -8.469194390390069e-13
+   -1.226454238991104e-12
+   -2.060748965656893e-11
+     8.20105722507647e-11
+ 2.55e+10    
+    8.214319756135091e-11
+   -2.060628411504458e-11
+    8.383150834978364e-11
+    -1.23421843869199e-12
+   -9.841283570054627e-12
+    8.385542581332851e-11
+   -8.500929986777478e-13
+   -1.229900626857548e-12
+   -2.060902544721001e-11
+    8.200801110655863e-11
+ 2.56e+10    
+    8.214062663910668e-11
+   -2.060784478873284e-11
+    8.383137514516993e-11
+   -1.237670342498222e-12
+   -9.842484762635295e-12
+    8.385527765778126e-11
+   -8.532473027573392e-13
+   -1.233346087306567e-12
+   -2.061057803473753e-11
+    8.200545060578334e-11
+ 2.57e+10    
+    8.213805602015525e-11
+   -2.060942218862245e-11
+    8.383125316894762e-11
+   -1.241121213277094e-12
+   -9.843699047393091e-12
+    8.385514098983197e-11
+   -8.563822462666878e-13
+   -1.236790560313661e-12
+   -2.061214740899378e-11
+    8.200289051988679e-11
+ 2.58e+10    
+    8.213548547771528e-11
+   -2.061101630489077e-11
+    8.383114224805368e-11
+    -1.24457099085399e-12
+   -9.844926417424633e-12
+    8.385501563087144e-11
+   -8.594977263645418e-13
+   -1.240233986205766e-12
+   -2.061373355907138e-11
+    8.200033062240154e-11
+ 2.59e+10    
+    8.213291478708181e-11
+   -2.061262712697011e-11
+    8.383104221134813e-11
+   -1.248019615398284e-12
+   -9.846166865039978e-12
+    8.385490140428247e-11
+   -8.625936423452051e-13
+   -1.243676305645949e-12
+   -2.061533647333141e-11
+    8.199777068892444e-11
+ 2.6e+10     
+    8.213034372560468e-11
+   -2.061425464356499e-11
+    8.383095288957679e-11
+    -1.25146702740838e-12
+   -9.847420381785866e-12
+    8.385479813540364e-11
+   -8.656698956045377e-13
+   -1.247117459618441e-12
+   -2.061695613942122e-11
+    8.199521049709561e-11
+ 2.61e+10    
+    8.212777207266813e-11
+   -2.061589884266974e-11
+    8.383087411533592e-11
+   -1.254913167697022e-12
+   -9.848686958468648e-12
+     8.38547056514943e-11
+   -8.687263896063106e-13
+   -1.250557389414025e-12
+   -2.061859254429201e-11
+     8.19926498265786e-11
+ 2.62e+10    
+    8.212519960966962e-11
+   -2.061755971158523e-11
+    8.383080572303683e-11
+   -1.258357977377037e-12
+   -9.849966585176386e-12
+    8.385462378169893e-11
+   -8.717630298488573e-13
+   -1.253996036615926e-12
+   -2.062024567421563e-11
+    8.199008845903931e-11
+ 2.63e+10    
+    8.212262611999913e-11
+   -2.061923723693516e-11
+    8.383074754887087e-11
+   -1.261801397847434e-12
+    -9.85125925130059e-12
+    8.385455235701324e-11
+   -8.747797238321004e-13
+   -1.257433343085946e-12
+   -2.062191551480117e-11
+    8.198752617812621e-11
+ 2.64e+10    
+    8.212005138901855e-11
+   -2.062093140468243e-11
+    8.383069943077672e-11
+   -1.265243370779844e-12
+   -9.852564945557456e-12
+    8.385449121025104e-11
+   -8.777763810248924e-13
+   -1.260869250950986e-12
+   -2.062360205101128e-11
+    8.198496276944981e-11
+ 2.65e+10    
+    8.211747520404096e-11
+   -2.062264220014463e-11
+    8.383066120840685e-11
+   -1.268683838105379e-12
+   -9.853883656008501e-12
+    8.385444017601075e-11
+    -8.80752912832683e-13
+   -1.264303702590009e-12
+   -2.062530526717793e-11
+    8.198239802056255e-11
+ 2.66e+10    
+    8.211489735431064e-11
+   -2.062436960800951e-11
+    8.383063272309539e-11
+   -1.272122742001765e-12
+   -9.855215370080859e-12
+    8.385439909064409e-11
+   -8.837092325655778e-13
+   -1.267736640621233e-12
+   -2.062702514701781e-11
+    8.197983172093902e-11
+ 2.67e+10    
+    8.211231763098192e-11
+   -2.062611361234989e-11
+    8.383061381782666e-11
+   -1.275560024880861e-12
+   -9.856560074587007e-12
+    8.385436779222397e-11
+   -8.866452554067055e-13
+    -1.27116800788975e-12
+   -2.062876167364737e-11
+    8.197726366195546e-11
+ 2.68e+10    
+    8.210973582709979e-11
+   -2.062787419663822e-11
+     8.38306043372049e-11
+   -1.278995629376508e-12
+   -9.857917755744046e-12
+    8.385434612051403e-11
+   -8.895608983809364e-13
+   -1.274597747455506e-12
+   -2.063051482959758e-11
+    8.197469363687049e-11
+ 2.69e+10    
+    8.210715173757924e-11
+     -2.0629651343761e-11
+    8.383060412742306e-11
+   -1.282429498332703e-12
+   -9.859288399192547e-12
+    8.385433391693832e-11
+   -8.924560803240047e-13
+   -1.278025802581476e-12
+   -2.063228459682811e-11
+     8.19721214408051e-11
+ 2.7e+10     
+     8.21045651591855e-11
+   -2.063144503603259e-11
+    8.383061303623432e-11
+   -1.285861574792095e-12
+   -9.860671990015024e-12
+     8.38543310245516e-11
+    -8.95330721851921e-13
+   -1.281452116722319e-12
+   -2.063407095674145e-11
+    8.196954687072322e-11
+ 2.71e+10    
+    8.210197589051441e-11
+   -2.063325525520886e-11
+    8.383063091292273e-11
+   -1.289291801984799e-12
+   -9.862068512753851e-12
+    8.385433728801076e-11
+   -8.981847453307911e-13
+   -1.284876633513257e-12
+   -2.063587389019646e-11
+    8.196696972541198e-11
+ 2.72e+10    
+    8.209938373197243e-11
+   -2.063508198250046e-11
+    8.383065760827525e-11
+   -1.292720123317534e-12
+   -9.863477951428904e-12
+    8.385435255354591e-11
+   -9.010180748469699e-13
+   -1.288299296759313e-12
+   -2.063769337752165e-11
+    8.196438980546281e-11
+ 2.73e+10    
+     8.20967884857571e-11
+    -2.06369251985856e-11
+    8.383069297455381e-11
+   -1.296146482363035e-12
+   -9.864900289554725e-12
+    8.385437666893289e-11
+   -9.038306361775972e-13
+   -1.291720050424794e-12
+   -2.063952939852806e-11
+    8.196180691325167e-11
+ 2.74e+10    
+    8.209418995583793e-11
+   -2.063878488362295e-11
+    8.383073686546882e-11
+   -1.299570822849812e-12
+   -9.866335510157321e-12
+    8.385440948346601e-11
+   -9.066223567614689e-13
+   -1.295138838623152e-12
+   -2.064138193252204e-11
+    8.195922085292063e-11
+ 2.75e+10    
+    8.209158794793695e-11
+   -2.064066101726358e-11
+    8.383078913615198e-11
+   -1.302993088652154e-12
+   -9.867783595790479e-12
+    8.385445084793075e-11
+   -9.093931656703152e-13
+   -1.298555605607087e-12
+   -2.064325095831723e-11
+    8.195663143035823e-11
+ 2.76e+10    
+    8.208898226950947e-11
+   -2.064255357866321e-11
+    8.383084964313143e-11
+   -1.306413223780441e-12
+   -9.869244528551972e-12
+    8.385450061457856e-11
+   -9.121429935803954e-13
+    -1.30197029575897e-12
+   -2.064513645424687e-11
+    8.195403845318132e-11
+ 2.77e+10    
+    8.208637272972547e-11
+   -2.064446254649373e-11
+    8.383091824430541e-11
+   -1.309831172371744e-12
+   -9.870718290099084e-12
+    8.385455863710041e-11
+   -9.148717727444983e-13
+   -1.305382853581467e-12
+   -2.064703839817526e-11
+    8.195144173071601e-11
+ 2.78e+10    
+    8.208375913945056e-11
+   -2.064638789895473e-11
+    8.383099479891782e-11
+   -1.313246878680726e-12
+   -9.872204861663946e-12
+    8.385462477060175e-11
+   -9.175794369642791e-13
+   -1.308793223688592e-12
+   -2.064895676750911e-11
+     8.19488410739795e-11
+ 2.79e+10    
+    8.208114131122748e-11
+   -2.064832961378451e-11
+    8.383107916753459e-11
+   -1.316660287070706e-12
+   -9.873704224068605e-12
+    8.385469887157802e-11
+   -9.202659215629968e-13
+   -1.312201350796883e-12
+    -2.06508915392086e-11
+     8.19462362956613e-11
+ 2.8e+10     
+    8.207851905925753e-11
+   -2.065028766827068e-11
+    8.383117121201873e-11
+   -1.320071342005181e-12
+   -9.875216357739495e-12
+    8.385478079789058e-11
+   -9.229311633585802e-13
+   -1.315607179716902e-12
+   -2.065284268979825e-11
+     8.19436272101054e-11
+ 2.81e+10    
+    8.207589219938223e-11
+   -2.065226203926109e-11
+    8.383127079550825e-11
+   -1.323479988039381e-12
+   -9.876741242721913e-12
+    8.385487040874272e-11
+   -9.255751006370902e-13
+   -1.319010655345029e-12
+   -2.065481019537721e-11
+     8.19410136332922e-11
+ 2.82e+10    
+    8.207326054906552e-11
+   -2.065425270317373e-11
+    8.383137778239244e-11
+   -1.326886169812282e-12
+   -9.878278858693829e-12
+    8.385496756465657e-11
+    -9.28197673126534e-13
+   -1.322411722655453e-12
+    -2.06567940316296e-11
+    8.193839538282055e-11
+ 2.83e+10    
+    8.207062392737543e-11
+   -2.065625963600687e-11
+    8.383149203829054e-11
+   -1.330289832038743e-12
+   -9.879829184979735e-12
+    8.385507212745043e-11
+   -9.307988219710582e-13
+   -1.325810326692449e-12
+   -2.065879417383427e-11
+    8.193577227788994e-11
+ 2.84e+10    
+    8.206798215496639e-11
+    -2.06582828133487e-11
+    8.383161343002899e-11
+   -1.333690919501908e-12
+    -9.88139220056383e-12
+    8.385518396021597e-11
+   -9.333784897054979e-13
+   -1.329206412562878e-12
+   -2.066081059687449e-11
+    8.193314413928315e-11
+ 2.85e+10    
+    8.206533505406139e-11
+   -2.066032221038669e-11
+    8.383174182562059e-11
+   -1.337089377045916e-12
+   -9.882967884103212e-12
+     8.38553029272972e-11
+    -9.35936620230273e-13
+   -1.332599925428974e-12
+   -2.066284327524742e-11
+    8.193051078934856e-11
+ 2.86e+10    
+    8.206268244843494e-11
+   -2.066237780191696e-11
+    8.383187709424361e-11
+   -1.340485149568765e-12
+   -9.884556213940624e-12
+    8.385542889426824e-11
+   -9.384731587866987e-13
+   -1.335990810501277e-12
+   -2.066489218307315e-11
+    8.192787205198345e-11
+ 2.87e+10    
+    8.206002416339561e-11
+   -2.066444956235309e-11
+    8.383201910622093e-11
+    -1.34387818201546e-12
+    -9.88615716811688e-12
+    8.385556172791273e-11
+   -9.409880519326111e-13
+   -1.339379013031892e-12
+   -2.066695729410344e-11
+    8.192522775261626e-11
+ 2.88e+10    
+    8.205736002576865e-11
+   -2.066653746573485e-11
+    8.383216773300032e-11
+   -1.347268419371361e-12
+   -9.887770724383128e-12
+    8.385570129620291e-11
+   -9.434812475183748e-13
+   -1.342764478307939e-12
+   -2.066903858173049e-11
+    8.192257771819018e-11
+ 2.89e+10    
+    8.205468986387956e-11
+   -2.066864148573661e-11
+     8.38323228471348e-11
+   -1.350655806655733e-12
+   -9.889396860212837e-12
+    8.385584746827974e-11
+   -9.459526946632607e-13
+   -1.346147151645168e-12
+   -2.067113601899527e-11
+    8.191992177714632e-11
+ 2.9e+10     
+    8.205201350753659e-11
+    -2.06707615956756e-11
+    8.383248432226329e-11
+   -1.354040288915598e-12
+   -9.891035552813378e-12
+    8.385600011443259e-11
+   -9.484023437321557e-13
+   -1.349526978381909e-12
+   -2.067324957859548e-11
+     8.19172597594068e-11
+ 2.91e+10    
+    8.204933078801499e-11
+    -2.06728977685199e-11
+    8.383265203309143e-11
+   -1.357421811219694e-12
+   -9.892686779137456e-12
+    8.385615910608013e-11
+   -9.508301463126653e-13
+   -1.352903903873121e-12
+   -2.067537923289371e-11
+    8.191459149635912e-11
+ 2.92e+10    
+    8.204664153803969e-11
+   -2.067504997689601e-11
+    8.383282585537369e-11
+   -1.360800318652724e-12
+   -9.894350515894348e-12
+    8.385632431575151e-11
+   -9.532360551925326e-13
+   -1.356277873484704e-12
+   -2.067752495392487e-11
+    8.191191682083885e-11
+ 2.93e+10    
+    8.204394559176989e-11
+   -2.067721819309671e-11
+    8.383300566589502e-11
+   -1.364175756309743e-12
+   -9.896026739560761e-12
+     8.38564956170671e-11
+   -9.556200243374666e-13
+   -1.359648832588018e-12
+    -2.06796867134037e-11
+    8.190923556711461e-11
+ 2.94e+10    
+    8.204124278478246e-11
+   -2.067940238908812e-11
+    8.383319134245307e-11
+   -1.367548069290817e-12
+   -9.897715426391473e-12
+    8.385667288472027e-11
+   -9.579820088692588e-13
+    -1.36301672655458e-12
+   -2.068186448273196e-11
+    8.190654757087144e-11
+ 2.95e+10    
+    8.203853295405635e-11
+   -2.068160253651686e-11
+     8.38333827638409e-11
+   -1.370917202695838e-12
+   -9.899416552429866e-12
+    8.385685599445996e-11
+   -9.603219650443157e-13
+   -1.366381500750955e-12
+   -2.068405823300551e-11
+    8.190385266919538e-11
+ 2.96e+10    
+    8.203581593795629e-11
+   -2.068381860671704e-11
+    8.383357980983015e-11
+   -1.374283101619457e-12
+   -9.901130093518105e-12
+    8.385704482307225e-11
+   -9.626398502324825e-13
+   -1.369743100533889e-12
+   -2.068626793502099e-11
+     8.19011507005582e-11
+ 2.97e+10    
+    8.203309157621825e-11
+   -2.068605057071683e-11
+    8.383378236115406e-11
+   -1.377645711146404e-12
+   -9.902856025307042e-12
+    8.385723924836365e-11
+   -9.649356228962673e-13
+   -1.373101471245537e-12
+   -2.068849355928241e-11
+    8.189844150480127e-11
+ 2.98e+10    
+    8.203035970993283e-11
+   -2.068829839924495e-11
+    8.383399029949133e-11
+   -1.381004976346805e-12
+   -9.904594323266113e-12
+    8.385743914914406e-11
+   -9.672092425703599e-13
+   -1.376456558208963e-12
+   -2.069073507600765e-11
+    8.189572492312093e-11
+ 2.99e+10    
+    8.202762018153124e-11
+   -2.069056206273706e-11
+    8.383420350744991e-11
+   -1.384360842271704e-12
+   -9.906344962692748e-12
+    8.385764440520952e-11
+   -9.694606698415557e-13
+   -1.379808306723781e-12
+   -2.069299245513443e-11
+    8.189300079805341e-11
+ 3e+10       
+    8.202487283476924e-11
+   -2.069284153134178e-11
+    8.383442186855192e-11
+   -1.387713253948905e-12
+   -9.908107918721887e-12
+    8.385785489732687e-11
+   -9.716898663289328e-13
+   -1.383156662061952e-12
+   -2.069526566632652e-11
+    8.189026897345962e-11
+ 3.01e+10    
+    8.202211751471312e-11
+   -2.069513677492671e-11
+    8.383464526721759e-11
+   -1.391062156378793e-12
+   -9.909883166334898e-12
+    8.385807050721691e-11
+   -9.738967946644664e-13
+   -1.386501569463823e-12
+   -2.069755467897939e-11
+    8.188752929451081e-11
+ 3.02e+10    
+    8.201935406772459e-11
+   -2.069744776308402e-11
+    8.383487358875065e-11
+   -1.394407494530454e-12
+   -9.911670680368727e-12
+    8.385829111753925e-11
+   -9.760814184739255e-13
+   -1.389842974134213e-12
+   -2.069985946222588e-11
+    8.188478160767372e-11
+ 3.03e+10    
+    8.201658234144627e-11
+   -2.069977446513612e-11
+    8.383510671932337e-11
+   -1.397749213337941e-12
+   -9.913470435524468e-12
+    8.385851661187655e-11
+   -9.782437023580811e-13
+   -1.393180821238829e-12
+   -2.070217998494165e-11
+    8.188202576069651e-11
+ 3.04e+10    
+    8.201380218478726e-11
+   -2.070211685014096e-11
+     8.38353445459621e-11
+   -1.401087257696629e-12
+   -9.915282406376012e-12
+    8.385874687471957e-11
+   -9.803836118743109e-13
+   -1.396515055900664e-12
+   -2.070451621575041e-11
+    8.187926160259421e-11
+ 3.05e+10    
+    8.201101344790954e-11
+   -2.070447488689733e-11
+    8.383558695653331e-11
+    -1.40442157245986e-12
+   -9.917106567378381e-12
+    8.385898179145257e-11
+   -9.825011135184822e-13
+   -1.399845623196714e-12
+   -2.070686812302903e-11
+    8.187648898363484e-11
+ 3.06e+10    
+    8.200821598221341e-11
+   -2.070684854394986e-11
+    8.383583383972968e-11
+   -1.407752102435595e-12
+   -9.918942892875867e-12
+    8.385922124833794e-11
+   -9.845961747071903e-13
+   -1.403172468154732e-12
+   -2.070923567491238e-11
+    8.187370775532564e-11
+ 3.07e+10    
+    8.200540964032345e-11
+   -2.070923778959382e-11
+    8.383608508505628e-11
+   -1.411078792383316e-12
+   -9.920791357110043e-12
+    8.385946513250292e-11
+   -9.866687637602866e-13
+   -1.406495535750224e-12
+   -2.071161883929824e-11
+    8.187091777039929e-11
+ 3.08e+10    
+    8.200259427607588e-11
+   -2.071164259187998e-11
+    8.383634058281723e-11
+   -1.414401587011096e-12
+   -9.922651934227624e-12
+    8.385971333192516e-11
+   -9.887188498837751e-13
+   -1.409814770903482e-12
+   -2.071401758385172e-11
+    8.186811888280008e-11
+ 3.09e+10    
+    8.199976974450366e-11
+   -2.071406291861901e-11
+    8.383660022410291e-11
+   -1.417720430972719e-12
+   -9.924524598288047e-12
+    8.385996573541903e-11
+   -9.907464031529806e-13
+   -1.413130118476896e-12
+   -2.071643187600991e-11
+    8.186531094767109e-11
+ 3.1e+10     
+     8.19969359018246e-11
+    -2.07164987373861e-11
+    8.383686390077696e-11
+   -1.421035268864994e-12
+   -9.926409323271009e-12
+    8.386022223262203e-11
+   -9.927513944960777e-13
+   -1.416441523272289e-12
+   -2.071886168298588e-11
+    8.186249382134023e-11
+ 3.11e+10    
+    8.199409260542712e-11
+   -2.071895001552498e-11
+    8.383713150546352e-11
+   -1.424346045225246e-12
+   -9.928306083083708e-12
+    8.386048271398161e-11
+   -9.947337956778891e-13
+   -1.419748930028508e-12
+   -2.072130697177307e-11
+    8.185966736130809e-11
+ 3.12e+10    
+    8.199123971385774e-11
+   -2.072141672015228e-11
+    8.383740293153558e-11
+   -1.427652704528885e-12
+   -9.930214851568113e-12
+    8.386074707074248e-11
+   -9.966935792840309e-13
+   -1.423052283418978e-12
+   -2.072376770914921e-11
+    8.185683142623418e-11
+ 3.13e+10    
+    8.198837708680807e-11
+   -2.072389881816121e-11
+    8.383767807310189e-11
+   -1.430955191187133e-12
+   -9.932135602507818e-12
+    8.386101519493349e-11
+   -9.986307187053425e-13
+   -1.426351528049612e-12
+   -2.072624386168004e-11
+    8.185398587592457e-11
+ 3.14e+10    
+    8.198550458510232e-11
+   -2.072639627622572e-11
+    8.383795682499615e-11
+   -1.434253449544873e-12
+   -9.934068309634967e-12
+    8.386128697935545e-11
+   -1.000545188122632e-12
+    -1.42964660845666e-12
+   -2.072873539572316e-11
+    8.185113057131951e-11
+ 3.15e+10    
+     8.19826220706847e-11
+   -2.072890906080391e-11
+    8.383823908276462e-11
+   -1.437547423878684e-12
+   -9.936012946636925e-12
+    8.386156231756854e-11
+   -1.002436962491711e-12
+   -1.432937469104786e-12
+   -2.073124227743153e-11
+    8.184826537448041e-11
+ 3.16e+10    
+    8.197972940660679e-11
+   -2.073143713814174e-11
+    8.383852474265513e-11
+   -1.440837058394846e-12
+   -9.937969487162835e-12
+    8.386184110388065e-11
+   -1.004306017528761e-12
+   -1.436224054385236e-12
+   -2.073376447275699e-11
+    8.184539014857837e-11
+ 3.17e+10    
+    8.197682645701606e-11
+    -2.07339804742765e-11
+    8.383881370160584e-11
+    -1.44412229722769e-12
+   -9.939937904829919e-12
+     8.38621232333354e-11
+   -1.006152329695953e-12
+   -1.439506308614134e-12
+   -2.073630194745343e-11
+    8.184250475788111e-11
+ 3.18e+10    
+    8.197391308714286e-11
+      -2.073653903504e-11
+    8.383910585723444e-11
+    -1.44740308443787e-12
+   -9.941918173229887e-12
+    8.386240860170049e-11
+   -1.007975876187382e-12
+    -1.44278417603092e-12
+   -2.073885466708003e-11
+    8.183960906774196e-11
+ 3.19e+10    
+    8.197098916328951e-11
+   -2.073911278606175e-11
+    8.383940110782691e-11
+   -1.450679364010874e-12
+   -9.943910265934895e-12
+    8.386269710545646e-11
+   -1.009776634915304e-12
+   -1.446057600796831e-12
+   -2.074142259700445e-11
+    8.183670294458743e-11
+ 3.2e+10     
+    8.196805455281778e-11
+   -2.074170169277218e-11
+    8.383969935232766e-11
+   -1.453951079855581e-12
+   -9.945914156503624e-12
+    8.386298864178536e-11
+   -1.011554584496631e-12
+   -1.449326526993599e-12
+   -2.074400570240551e-11
+    8.183378625590579e-11
+ 3.21e+10    
+    8.196510912413794e-11
+   -2.074430572040544e-11
+    8.384000049032893e-11
+   -1.457218175802978e-12
+   -9.947929818487079e-12
+    8.386328310856032e-11
+   -1.013309704239736e-12
+   -1.452590898622187e-12
+   -2.074660394827624e-11
+    8.183085887023535e-11
+ 3.22e+10    
+    8.196215274669676e-11
+   -2.074692483400221e-11
+    8.384030442206031e-11
+   -1.460480595604951e-12
+   -9.949957225434283e-12
+    8.386358040433384e-11
+   -1.015041974131527e-12
+   -1.455850659601645e-12
+   -2.074921729942642e-11
+    8.182792065715349e-11
+ 3.23e+10    
+    8.195918529096686e-11
+   -2.074955899841253e-11
+    8.384061104837947e-11
+   -1.463738282933211e-12
+     -9.9519963508979e-12
+    8.386388042832844e-11
+   -1.016751374824808e-12
+   -1.459105753768082e-12
+   -2.075184572048529e-11
+    8.182497148726505e-11
+ 3.24e+10    
+    8.195620662843499e-11
+   -2.075220817829833e-11
+     8.38409202707619e-11
+   -1.466991181378288e-12
+   -9.954047168439669e-12
+    8.386418308042514e-11
+   -1.018437887625907e-12
+   -1.462356124873758e-12
+   -2.075448917590396e-11
+    8.182201123219151e-11
+ 3.25e+10    
+     8.19532166315915e-11
+   -2.075487233813591e-11
+     8.38412319912915e-11
+   -1.470239234448713e-12
+   -9.956109651635719e-12
+    8.386448826115408e-11
+   -1.020101494482558e-12
+   -1.465601716586248e-12
+   -2.075714762995777e-11
+    8.181903976455991e-11
+ 3.26e+10    
+    8.195021517391912e-11
+   -2.075755144221841e-11
+    8.384154611265147e-11
+   -1.473482385570137e-12
+   -9.958183774081805e-12
+    8.386479587168446e-11
+   -1.021742177972116e-12
+   -1.468842472487718e-12
+   -2.075982104674869e-11
+    8.181605695799234e-11
+ 3.27e+10    
+    8.194720212988292e-11
+   -2.076024545465808e-11
+    8.384186253811486e-11
+   -1.476720578084735e-12
+   -9.960269509398416e-12
+    8.386510581381444e-11
+   -1.023359921289969e-12
+   -1.472078336074312e-12
+   -2.076250939020728e-11
+    8.181306268709487e-11
+ 3.28e+10    
+      8.1944177374919e-11
+   -2.076295433938837e-11
+    8.384218117153543e-11
+   -1.479953755250597e-12
+   -9.962366831235682e-12
+    8.386541798996153e-11
+   -1.024954708238249e-12
+   -1.475309250755581e-12
+   -2.076521262409495e-11
+    8.181005682744754e-11
+ 3.29e+10    
+    8.194114078542456e-11
+    -2.07656780601662e-11
+    8.384250191733917e-11
+   -1.483181860241221e-12
+   -9.964475713278321e-12
+    8.386573230315374e-11
+   -1.026526523214787e-12
+    -1.47853515985408e-12
+    -2.07679307120059e-11
+    8.180703925559371e-11
+ 3.3e+10     
+    8.193809223874755e-11
+   -2.076841658057379e-11
+    8.384282468051534e-11
+   -1.486404836145115e-12
+   -9.966596129250328e-12
+    8.386604865701961e-11
+   -1.028075351202353e-12
+   -1.481756006605018e-12
+   -2.077066361736884e-11
+    8.180400984902977e-11
+ 3.31e+10    
+    8.193503161317668e-11
+   -2.077116986402071e-11
+    8.384314936660807e-11
+     -1.4896226259655e-12
+   -9.968728052919627e-12
+    8.386636695577947e-11
+   -1.029601177758131e-12
+   -1.484971734155965e-12
+   -2.077341130344901e-11
+    8.180096848619538e-11
+ 3.32e+10    
+    8.193195878793105e-11
+   -2.077393787374553e-11
+    8.384347588170789e-11
+   -1.492835172620076e-12
+    -9.97087145810261e-12
+    8.386668710423662e-11
+    -1.03110398900342e-12
+   -1.488182285566698e-12
+   -2.077617373334977e-11
+    8.179791504646349e-11
+ 3.33e+10    
+    8.192887364315079e-11
+   -2.077672057281785e-11
+    8.384380413244388e-11
+    -1.49604241894087e-12
+    -9.97302631866856e-12
+    8.386700900776803e-11
+   -1.032583771613646e-12
+   -1.491387603809124e-12
+    -2.07789508700141e-11
+    8.179484941012999e-11
+ 3.34e+10    
+    8.192577605988692e-11
+   -2.077951792413951e-11
+    8.384413402597518e-11
+   -1.499244307674207e-12
+   -9.975192608543992e-12
+    8.386733257231653e-11
+   -1.034040512808571e-12
+   -1.494587631767231e-12
+   -2.078174267622638e-11
+    8.179177145840493e-11
+ 3.35e+10    
+    8.192266592009241e-11
+    -2.07823298904466e-11
+    8.384446546998335e-11
+   -1.502440781480714e-12
+   -9.977370301716816e-12
+    8.386765770438184e-11
+   -1.035474200342752e-12
+   -1.497782312237192e-12
+   -2.078454911461362e-11
+    8.178868107340198e-11
+ 3.36e+10    
+    8.191954310661181e-11
+   -2.078515643431061e-11
+    8.384479837266469e-11
+   -1.505631782935427e-12
+   -9.979559372240529e-12
+    8.386798431101212e-11
+   -1.036884822496266e-12
+   -1.500971587927509e-12
+   -2.078737014764687e-11
+    8.178557813812992e-11
+ 3.37e+10    
+    8.191640750317278e-11
+   -2.078799751814004e-11
+    8.384513264272243e-11
+   -1.508817254527983e-12
+   -9.981759794238199e-12
+    8.386831229979655e-11
+    -1.03827236806563e-12
+   -1.504155401459224e-12
+   -2.079020573764269e-11
+    8.178246253648291e-11
+ 3.38e+10    
+    8.191325899437643e-11
+   -2.079085310418152e-11
+    8.384546818935949e-11
+   -1.511997138662856e-12
+   -9.983971541906347e-12
+    8.386864157885637e-11
+   -1.039636826355001e-12
+   -1.507333695366245e-12
+   -2.079305584676403e-11
+     8.17793341532313e-11
+ 3.39e+10    
+    8.191009746568846e-11
+   -2.079372315452127e-11
+    8.384580492227083e-11
+   -1.515171377659725e-12
+   -9.986194589518878e-12
+     8.38689720568381e-11
+   -1.040978187167568e-12
+    -1.51050641209569e-12
+   -2.079592043702171e-11
+    8.177619287401271e-11
+ 3.4e+10     
+    8.190692280343051e-11
+   -2.079660763108625e-11
+    8.384614275163676e-11
+   -1.518339913753846e-12
+   -9.988428911430717e-12
+    8.386930364290476e-11
+     -1.0422964407972e-12
+   -1.513673494008359e-12
+   -2.079879947027515e-11
+    8.177303858532308e-11
+ 3.41e+10    
+    8.190373489477049e-11
+   -2.079950649564503e-11
+    8.384648158811567e-11
+   -1.521502689096519e-12
+   -9.990674482081566e-12
+    8.386963624672921e-11
+   -1.043591578020298e-12
+   -1.516834883379224e-12
+   -2.080169290823371e-11
+    8.176987117450798e-11
+ 3.42e+10    
+    8.190053362771486e-11
+   -2.080241970980911e-11
+    8.384682134283677e-11
+   -1.524659645755678e-12
+   -9.992931275999308e-12
+    8.386996977848625e-11
+   -1.044863590087892e-12
+   -1.519990522398036e-12
+   -2.080460071245734e-11
+    8.176669052975383e-11
+ 3.43e+10    
+    8.189731889109962e-11
+   -2.080534723503376e-11
+    8.384716192739388e-11
+   -1.527810725716434e-12
+   -9.995199267803614e-12
+      8.3870304148845e-11
+   -1.046112468717941e-12
+   -1.523140353169962e-12
+   -2.080752284435749e-11
+    8.176349654007943e-11
+ 3.44e+10    
+    8.189409057458191e-11
+   -2.080828903261898e-11
+    8.384750325383858e-11
+    -1.53095587088182e-12
+   -9.997478432209311e-12
+    8.387063926896265e-11
+   -1.047338206087845e-12
+   -1.526284317716293e-12
+   -2.081045926519811e-11
+    8.176028909532753e-11
+ 3.45e+10    
+    8.189084856863166e-11
+   -2.081124506371019e-11
+     8.38478452346733e-11
+   -1.534095023073474e-12
+   -9.999768744029554e-12
+    8.387097505047668e-11
+   -1.048540794827191e-12
+   -1.529422357975213e-12
+   -2.081340993609609e-11
+    8.175706808615626e-11
+ 3.46e+10    
+    8.188759276452342e-11
+   -2.081421528929915e-11
+    8.384818778284521e-11
+   -1.537228124032452e-12
+   -1.000207017817918e-11
+    8.387131140549798e-11
+    -1.04972022801071e-12
+   -1.532554415802656e-12
+   -2.081637481802207e-11
+    8.175383340403156e-11
+ 3.47e+10    
+    8.188432305432851e-11
+   -2.081719967022476e-11
+    8.384853081174037e-11
+   -1.540355115420131e-12
+   -1.000438270967782e-11
+    8.387164824660464e-11
+   -1.050876499151401e-12
+   -1.535680432973212e-12
+   -2.081935387180118e-11
+     8.17505849412186e-11
+ 3.48e+10    
+    8.188103933090667e-11
+   -2.082019816717338e-11
+    8.384887423517639e-11
+   -1.543475938819077e-12
+   -1.000670631365284e-11
+    8.387198548683451e-11
+   -1.052009602193923e-12
+   -1.538800351181033e-12
+   -2.082234705811325e-11
+    8.174732259077365e-11
+ 3.49e+10    
+    8.187774148789847e-11
+   -2.082321074067984e-11
+    8.384921796739747e-11
+   -1.546590535734036e-12
+   -1.000904096534245e-11
+     8.38723230396792e-11
+   -1.053119531508153e-12
+   -1.541914112040874e-12
+   -2.082535433749372e-11
+    8.174404624653702e-11
+ 3.5e+10     
+    8.187442941971748e-11
+   -2.082623735112769e-11
+    8.384956192306806e-11
+   -1.549698847592989e-12
+   -1.001138664009852e-11
+    8.387266081907737e-11
+   -1.054206281882924e-12
+   -1.545021657089207e-12
+   -2.082837567033369e-11
+     8.17407558031244e-11
+ 3.51e+10    
+     8.18711030215425e-11
+   -2.082927795874979e-11
+    8.384990601726657e-11
+   -1.552800815748235e-12
+    -1.00137433133894e-11
+    8.387299873940852e-11
+   -1.055269848520017e-12
+   -1.548122927785252e-12
+   -2.083141101688059e-11
+    8.173745115591975e-11
+ 3.52e+10    
+    8.186776218931052e-11
+    -2.08323325236288e-11
+    8.385025016548047e-11
+   -1.555896381477521e-12
+   -1.001611096080275e-11
+    8.387333671548696e-11
+   -1.056310227028312e-12
+   -1.551217865512201e-12
+   -2.083446033723847e-11
+    8.173413220106789e-11
+ 3.53e+10    
+    8.186440681970853e-11
+   -2.083540100569741e-11
+    8.385059428359956e-11
+   -1.558985485985236e-12
+     -1.0018489558048e-11
+    8.387367466255507e-11
+   -1.057327413418123e-12
+   -1.554306411578469e-12
+   -2.083752359136803e-11
+    8.173079883546651e-11
+ 3.54e+10    
+    8.186103681016705e-11
+   -2.083848336473892e-11
+    8.385093828791184e-11
+    -1.56206807040368e-12
+   -1.002087908095927e-11
+    8.387401249627817e-11
+   -1.058321404095738e-12
+   -1.557388507218902e-12
+   -2.084060073908729e-11
+    8.172745095675958e-11
+ 3.55e+10    
+    8.185765205885233e-11
+   -2.084157956038726e-11
+    8.385128209509641e-11
+   -1.565144075794332e-12
+   -1.002327950549752e-11
+    8.387435013273813e-11
+   -1.059292195858159e-12
+   -1.560464093596149e-12
+   -2.084369174007144e-11
+    8.172408846332932e-11
+ 3.56e+10    
+    8.185425246465938e-11
+   -2.084468955212745e-11
+    8.385162562221975e-11
+   -1.568213443149209e-12
+   -1.002569080775334e-11
+    8.387468748842737e-11
+   -1.060239785887992e-12
+   -1.563533111802025e-12
+   -2.084679655385303e-11
+    8.172071125429002e-11
+ 3.57e+10    
+    8.185083792720517e-11
+   -2.084781329929559e-11
+    8.385196878672902e-11
+   -1.571276113392264e-12
+   -1.002811296394909e-11
+    8.387502448024373e-11
+   -1.061164171748533e-12
+    -1.56659550285893e-12
+   -2.084991513982227e-11
+    8.171731922948021e-11
+ 3.58e+10    
+    8.184740834682151e-11
+   -2.085095076107922e-11
+    8.385231150644819e-11
+   -1.574332027380797e-12
+   -1.003054595044137e-11
+    8.387536102548479e-11
+   -1.062065351379066e-12
+   -1.569651207721277e-12
+   -2.085304745722688e-11
+    8.171391228945622e-11
+ 3.59e+10    
+    8.184396362454819e-11
+   -2.085410189651726e-11
+    8.385265369957178e-11
+   -1.577381125906945e-12
+   -1.003298974372317e-11
+    8.387569704184172e-11
+   -1.062943323090267e-12
+   -1.572700167277046e-12
+    -2.08561934651721e-11
+    8.171049033548523e-11
+ 3.6e+10     
+    8.184050366212684e-11
+   -2.085726666450025e-11
+    8.385299528466099e-11
+   -1.580423349699204e-12
+   -1.003544432042615e-11
+    8.387603244739482e-11
+   -1.063798085559859e-12
+     -1.5757423223493e-12
+   -2.085935312262089e-11
+    8.170705326953861e-11
+ 3.61e+10    
+     8.18370283619936e-11
+   -2.086044502377017e-11
+    8.385333618063797e-11
+   -1.583458639424018e-12
+   -1.003790965732268e-11
+    8.387636716060785e-11
+   -1.064629637828373e-12
+   -1.578777613697777e-12
+   -2.086252638839359e-11
+    8.170360099428504e-11
+ 3.62e+10    
+    8.183353762727298e-11
+   -2.086363693292058e-11
+    8.385367630678154e-11
+   -1.586486935687346e-12
+   -1.004038573132789e-11
+    8.387670110032229e-11
+   -1.065437979295119e-12
+   -1.581805982020535e-12
+   -2.086571322116792e-11
+     8.17001334130845e-11
+ 3.63e+10    
+    8.183003136177135e-11
+   -2.086684235039647e-11
+      8.3854015582722e-11
+   -1.589508179036323e-12
+   -1.004287251950177e-11
+    8.387703418575322e-11
+   -1.066223109714314e-12
+   -1.584827367955585e-12
+   -2.086891357947897e-11
+     8.16966504299814e-11
+ 3.64e+10    
+    8.182650946997065e-11
+   -2.087006123449426e-11
+    8.385435392843701e-11
+   -1.592522309960956e-12
+   -1.004536999905098e-11
+    8.387736633648353e-11
+   -1.066985029191358e-12
+    -1.58784171208265e-12
+   -2.087212742171883e-11
+    8.169315194969845e-11
+ 3.65e+10    
+    8.182297185702225e-11
+   -2.087329354336163e-11
+    8.385469126424692e-11
+   -1.595529268895831e-12
+   -1.004787814733079e-11
+    8.387769747245918e-11
+    -1.06772373817928e-12
+   -1.590848954924851e-12
+   -2.087535470613639e-11
+    8.168963787763025e-11
+ 3.66e+10    
+    8.181941842874068e-11
+   -2.087653923499736e-11
+    8.385502751080976e-11
+   -1.598528996221861e-12
+   -1.005039694184682e-11
+    8.387802751398474e-11
+   -1.068439237475374e-12
+   -1.593849036950513e-12
+   -2.087859539083731e-11
+    8.168610811983732e-11
+ 3.67e+10    
+    8.181584909159774e-11
+   -2.087979826725118e-11
+    8.385536258911752e-11
+   -1.601521432268114e-12
+   -1.005292636025692e-11
+    8.387835638171785e-11
+   -1.069131528217915e-12
+   -1.596841898574971e-12
+   -2.088184943378342e-11
+    8.168256258303972e-11
+ 3.68e+10    
+    8.181226375271609e-11
+   -2.088307059782341e-11
+    8.385569642049169e-11
+   -1.604506517313598e-12
+   -1.005546638037274e-11
+    8.387868399666517e-11
+    -1.06980061188313e-12
+   -1.599827480162415e-12
+   -2.088511679279275e-11
+    8.167900117461173e-11
+ 3.69e+10    
+    8.180866231986399e-11
+   -2.088635618426496e-11
+    8.385602892657892e-11
+   -1.607484191589154e-12
+   -1.005801698016145e-11
+    8.387901028017761e-11
+   -1.070446490282214e-12
+   -1.602805722027788e-12
+   -2.088839742553886e-11
+      8.1675423802575e-11
+ 3.7e+10     
+    8.180504470144901e-11
+   -2.088965498397672e-11
+    8.385636002934646e-11
+   -1.610454395279334e-12
+   -1.006057813774722e-11
+    8.387933515394568e-11
+   -1.071069165558586e-12
+   -1.605776564438657e-12
+   -2.089169128955072e-11
+    8.167183037559345e-11
+ 3.71e+10    
+    8.180141080651271e-11
+   -2.089296695420952e-11
+    8.385668965107885e-11
+   -1.613417068524312e-12
+    -1.00631498314129e-11
+    8.387965853999511e-11
+   -1.071668640185244e-12
+   -1.608739947617181e-12
+   -2.089499834221219e-11
+    8.166822080296743e-11
+ 3.72e+10    
+    8.179776054472479e-11
+   -2.089629205206365e-11
+    8.385701771437313e-11
+   -1.616372151421874e-12
+   -1.006573203960133e-11
+    8.387998036068255e-11
+   -1.072244916962265e-12
+   -1.611695811742066e-12
+   -2.089831854076167e-11
+    8.166459499462792e-11
+ 3.73e+10    
+    8.179409382637742e-11
+   -2.089963023448851e-11
+    8.385734414213566e-11
+   -1.619319584029361e-12
+    -1.00683247409169e-11
+      8.3880300538691e-11
+   -1.072797999014461e-12
+   -1.614644096950582e-12
+    -2.09016518422915e-11
+    8.166095286113061e-11
+ 3.74e+10    
+    8.179041056238016e-11
+   -2.090298145828227e-11
+    8.385766885757755e-11
+   -1.622259306365722e-12
+   -1.007092791412682e-11
+    8.388061899702603e-11
+   -1.073327889789174e-12
+   -1.617584743340574e-12
+   -2.090499820374773e-11
+    8.165729431365144e-11
+ 3.75e+10    
+    8.178671066425413e-11
+   -2.090634568009129e-11
+     8.38579917842112e-11
+   -1.625191258413498e-12
+   -1.007354153816246e-11
+    8.388093565901105e-11
+   -1.073834593054203e-12
+   -1.620517690972524e-12
+   -2.090835758192933e-11
+    8.165361926398014e-11
+ 3.76e+10    
+    8.178299404412706e-11
+   -2.090972285640987e-11
+    8.385831284584632e-11
+   -1.628115380120947e-12
+   -1.007616559212064e-11
+     8.38812504482838e-11
+   -1.074318112895869e-12
+   -1.623442879871603e-12
+   -2.091172993348787e-11
+    8.164992762451522e-11
+ 3.77e+10    
+    8.177926061472787e-11
+   -2.091311294357959e-11
+    8.385863196658637e-11
+   -1.631031611404114e-12
+   -1.007880005526479e-11
+    8.388156328879202e-11
+     -1.0747784537172e-12
+   -1.626360250029828e-12
+   -2.091511521492693e-11
+    8.164621930825907e-11
+ 3.78e+10    
+    8.177551028938167e-11
+   -2.091651589778911e-11
+    8.385894907082517e-11
+   -1.633939892148917e-12
+    -1.00814449070262e-11
+    8.388187410478942e-11
+   -1.075215620236283e-12
+   -1.629269741408133e-12
+   -2.091851338260147e-11
+    8.164249422881243e-11
+ 3.79e+10    
+    8.177174298200459e-11
+   -2.091993167507318e-11
+    8.385926408324256e-11
+   -1.636840162213342e-12
+     -1.0084100127005e-11
+    8.388218282083203e-11
+     -1.0756296174847e-12
+   -1.632171293938569e-12
+   -2.092192439271727e-11
+    8.163875230036915e-11
+ 3.8e+10     
+    8.176795860709821e-11
+   -2.092336023131256e-11
+    8.385957692880215e-11
+   -1.639732361429567e-12
+   -1.008676569497139e-11
+    8.388248936177418e-11
+   -1.076020450806108e-12
+   -1.635064847526453e-12
+   -2.092534820133038e-11
+    8.163499343771164e-11
+ 3.81e+10    
+    8.176415707974608e-11
+   -2.092680152223324e-11
+     8.38598875327464e-11
+   -1.642616429606151e-12
+   -1.008944159086652e-11
+    8.388279365276483e-11
+   -1.076388125854981e-12
+   -1.637950342052555e-12
+   -2.092878476434631e-11
+    8.163121755620528e-11
+ 3.82e+10    
+    8.176033831560708e-11
+   -2.093025550340581e-11
+    8.386019582059446e-11
+   -1.645492306530272e-12
+   -1.009212779480356e-11
+    8.388309561924374e-11
+   -1.076732648595388e-12
+   -1.640827717375351e-12
+   -2.093223403751959e-11
+     8.16274245717941e-11
+ 3.83e+10    
+    8.175650223091213e-11
+   -2.093372213024509e-11
+    8.386050171813812e-11
+   -1.648359931969917e-12
+   -1.009482428706857e-11
+     8.38833951869384e-11
+   -1.077054025299996e-12
+   -1.643696913333228e-12
+   -2.093569597645305e-11
+     8.16236144009958e-11
+ 3.84e+10    
+    8.175264874245854e-11
+   -2.093720135800924e-11
+    8.386080515143866e-11
+   -1.651219245676182e-12
+   -1.009753104812137e-11
+    8.388369228185946e-11
+   -1.077352262549093e-12
+   -1.646557869746745e-12
+   -2.093917053659689e-11
+    8.161978696089635e-11
+ 3.85e+10    
+    8.174877776760553e-11
+   -2.094069314179935e-11
+    8.386110604682381e-11
+   -1.654070187385459e-12
+   -1.010024805859644e-11
+    8.388398683029809e-11
+   -1.077627367229809e-12
+   -1.649410526420931e-12
+   -2.094265767324842e-11
+     8.16159421691466e-11
+ 3.86e+10    
+     8.17448892242699e-11
+   -2.094419743655865e-11
+    8.386140433088461e-11
+   -1.656912696821813e-12
+   -1.010297529930373e-11
+    8.388427875882225e-11
+    -1.07787934653538e-12
+   -1.652254823147549e-12
+   -2.094615734155091e-11
+    8.161207994395619e-11
+ 3.87e+10    
+    8.174098303092135e-11
+   -2.094771419707191e-11
+    8.386169993047184e-11
+   -1.659746713699218e-12
+   -1.010571275122924e-11
+    8.388456799427309e-11
+   -1.078108207964595e-12
+   -1.655090699707437e-12
+    -2.09496694964932e-11
+    8.160820020409026e-11
+ 3.88e+10    
+    8.173705910657798e-11
+   -2.095124337796472e-11
+    8.386199277269343e-11
+   -1.662572177723925e-12
+   -1.010846039553592e-11
+    8.388485446376151e-11
+   -1.078313959321284e-12
+   -1.657918095872813e-12
+   -2.095319409290861e-11
+    8.160430286886408e-11
+ 3.89e+10    
+    8.173311737080185e-11
+   -2.095478493370288e-11
+    8.386228278491146e-11
+   -1.665389028596766e-12
+   -1.011121821356431e-11
+    8.388513809466573e-11
+   -1.078496608713956e-12
+   -1.660736951409631e-12
+   -2.095673108547452e-11
+    8.160038785813905e-11
+ 3.9e+10     
+    8.172915774369485e-11
+    -2.09583388185915e-11
+    8.386256989473849e-11
+   -1.668197206015545e-12
+   -1.011398618683303e-11
+    8.388541881462701e-11
+   -1.078656164555544e-12
+   -1.663547206079914e-12
+   -2.096028042871139e-11
+     8.15964550923181e-11
+ 3.91e+10    
+    8.172518014589414e-11
+   -2.096190498677451e-11
+    8.386285403003556e-11
+   -1.670996649677359e-12
+   -1.011676429703949e-11
+    8.388569655154681e-11
+   -1.078792635563232e-12
+   -1.666348799644187e-12
+   -2.096384207698199e-11
+    8.159250449234172e-11
+ 3.92e+10    
+     8.17211844985683e-11
+   -2.096548339223379e-11
+    8.386313511890887e-11
+   -1.673787299281009e-12
+    -1.01195525260604e-11
+    8.388597123358386e-11
+   -1.078906030758389e-12
+   -1.669141671863797e-12
+   -2.096741598449055e-11
+    8.158853597968306e-11
+ 3.93e+10    
+    8.171717072341272e-11
+   -2.096907398878841e-11
+    8.386341308970681e-11
+   -1.676569094529411e-12
+   -1.012235085595229e-11
+    8.388624278915124e-11
+   -1.078996359466624e-12
+    -1.67192576250335e-12
+   -2.097100210528221e-11
+    8.158454947634474e-11
+ 3.94e+10    
+    8.171313874264588e-11
+   -2.097267673009394e-11
+     8.38636878710176e-11
+   -1.679341975131981e-12
+   -1.012515926895194e-11
+    8.388651114691254e-11
+   -1.079063631317912e-12
+   -1.674701011333115e-12
+   -2.097460039324186e-11
+     8.15805449048536e-11
+ 3.95e+10    
+    8.170908847900532e-11
+   -2.097629156964164e-11
+    8.386395939166592e-11
+   -1.682105880807057e-12
+   -1.012797774747679e-11
+    8.388677623577967e-11
+   -1.079107856246831e-12
+    -1.67746735813145e-12
+   -2.097821080209349e-11
+    8.157652218825751e-11
+ 3.96e+10    
+    8.170501985574326e-11
+   -2.097991846075763e-11
+    8.386422758071086e-11
+   -1.684860751284354e-12
+   -1.013080627412543e-11
+    8.388703798490971e-11
+   -1.079129044492895e-12
+   -1.680224742687236e-12
+   -2.098183328539934e-11
+    8.157248125012078e-11
+ 3.97e+10    
+    8.170093279662317e-11
+   -2.098355735660223e-11
+    8.386449236744309e-11
+   -1.687606526307393e-12
+   -1.013364483167784e-11
+    8.388729632370154e-11
+   -1.079127206600976e-12
+   -1.682973104802333e-12
+     -2.0985467796559e-11
+     8.15684220145208e-11
+ 3.98e+10    
+    8.169682722591558e-11
+   -2.098720821016907e-11
+    8.386475368138192e-11
+   -1.690343145635958e-12
+   -1.013649340309577e-11
+    8.388755118179402e-11
+   -1.079102353421797e-12
+   -1.685712384294016e-12
+   -2.098911428880859e-11
+    8.156434440604333e-11
+ 3.99e+10    
+    8.169270306839421e-11
+   -2.099087097428416e-11
+    8.386501145227315e-11
+   -1.693070549048569e-12
+     -1.0139351971523e-11
+    8.388780248906206e-11
+   -1.079054496112554e-12
+   -1.688442520997472e-12
+   -2.099277271521986e-11
+    8.156024834977915e-11
+ 4e+10       
+    8.168856024933281e-11
+   -2.099454560160547e-11
+    8.386526561008631e-11
+   -1.695788676344943e-12
+   -1.014222052028558e-11
+     8.38880501756144e-11
+   -1.078983646137602e-12
+   -1.691163454768246e-12
+   -2.099644302869928e-11
+    8.155613377132053e-11
+ 4.01e+10    
+    8.168439869450044e-11
+   -2.099823204462153e-11
+    8.386551608501219e-11
+   -1.698497467348514e-12
+   -1.014509903289207e-11
+    8.388829417179139e-11
+    -1.07888981526921e-12
+   -1.693875125484733e-12
+   -2.100012518198734e-11
+    8.155200059675672e-11
+ 4.02e+10    
+    8.168021833015867e-11
+   -2.100193025565114e-11
+    8.386576280746046e-11
+   -1.701196861908866e-12
+   -1.014798749303363e-11
+    8.388853440816109e-11
+   -1.078773015588435e-12
+     -1.6965774730507e-12
+   -2.100381912765736e-11
+    8.154784875267091e-11
+ 4.03e+10    
+    8.167601908305764e-11
+   -2.100564018684217e-11
+     8.38660057080573e-11
+   -1.703886799904292e-12
+    -1.01508858845843e-11
+    8.388877081551781e-11
+   -1.078633259486056e-12
+   -1.699270437397729e-12
+    -2.10075248181149e-11
+    8.154367816613627e-11
+ 4.04e+10    
+     8.16718008804325e-11
+    -2.10093617901709e-11
+    8.386624471764296e-11
+   -1.706567221244258e-12
+   -1.015379419160097e-11
+    8.388900332487885e-11
+   -1.078470559663584e-12
+   -1.701953958487768e-12
+   -2.101124220559663e-11
+    8.153948876471235e-11
+ 4.05e+10    
+    8.166756364999994e-11
+   -2.101309501744109e-11
+    8.386647976726903e-11
+   -1.709238065871957e-12
+    -1.01567123983235e-11
+    8.388923186748235e-11
+   -1.078284929134368e-12
+   -1.704627976315629e-12
+   -2.101497124216956e-11
+    8.153528047644175e-11
+ 4.06e+10    
+    8.166330731995471e-11
+   -2.101683982028315e-11
+    8.386671078819712e-11
+   -1.711899273766796e-12
+   -1.015964048917482e-11
+    8.388945637478449e-11
+   -1.078076381224754e-12
+   -1.707292430911494e-12
+   -2.101871187973011e-11
+    8.153105322984633e-11
+ 4.07e+10    
+    8.165903181896636e-11
+   -2.102059615015332e-11
+    8.386693771189569e-11
+   -1.714550784946927e-12
+   -1.016257844876087e-11
+    8.388967677845695e-11
+    -1.07784492957535e-12
+   -1.709947262343483e-12
+   -2.102246407000306e-11
+    8.152680695392406e-11
+ 4.08e+10    
+    8.165473707617537e-11
+   -2.102436395833266e-11
+    8.386716047003806e-11
+   -1.717192539471791e-12
+   -1.016552626187059e-11
+    8.388989301038486e-11
+   -1.077590588142332e-12
+   -1.712592410720102e-12
+   -2.102622776454088e-11
+    8.152254157814528e-11
+ 4.09e+10    
+    8.165042302119044e-11
+   -2.102814319592636e-11
+    8.386737899450045e-11
+   -1.719824477444646e-12
+   -1.016848391347588e-11
+    8.389010500266422e-11
+   -1.077313371198834e-12
+   -1.715227816192856e-12
+   -2.103000291472261e-11
+    8.151825703244956e-11
+ 4.1e+10     
+    8.164608958408506e-11
+    -2.10319338138628e-11
+    8.386759321735948e-11
+   -1.722446539015117e-12
+   -1.017145138873154e-11
+    8.389031268759946e-11
+   -1.077013293336426e-12
+   -1.717853418958722e-12
+     -2.1033789471753e-11
+    8.151395324724228e-11
+ 4.11e+10    
+    8.164173669539383e-11
+   -2.103573576289254e-11
+    8.386780307089034e-11
+    -1.72505866438172e-12
+   -1.017442867297506e-11
+    8.389051599770091e-11
+   -1.076690369466627e-12
+   -1.720469159262752e-12
+   -2.103758738666156e-11
+    8.150963015339159e-11
+ 4.12e+10    
+    8.163736428610988e-11
+   -2.103954899358775e-11
+     8.38680084875644e-11
+   -1.727660793794416e-12
+    -1.01774157517266e-11
+    8.389071486568324e-11
+   -1.076344614822503e-12
+   -1.723074977400551e-12
+    -2.10413966103017e-11
+    8.150528768222465e-11
+ 4.13e+10    
+     8.16329722876813e-11
+   -2.104337345634097e-11
+    8.386820940004742e-11
+    -1.73025286755718e-12
+   -1.018041261068875e-11
+    8.389090922446251e-11
+   -1.075976044960334e-12
+   -1.725670813720859e-12
+   -2.104521709334979e-11
+    8.150092576552516e-11
+ 4.14e+10    
+    8.162856063200824e-11
+   -2.104720910136453e-11
+    8.386840574119735e-11
+   -1.732834826030519e-12
+   -1.018341923574634e-11
+    8.389109900715407e-11
+   -1.075584675761328e-12
+    -1.72825660862809e-12
+   -2.104904878630406e-11
+    8.149654433552937e-11
+ 4.15e+10    
+    8.162412925143981e-11
+   -2.105105587868948e-11
+    8.386859744406237e-11
+   -1.735406609634042e-12
+   -1.018643561296618e-11
+    8.389128414707067e-11
+   -1.075170523433427e-12
+   -1.730832302584884e-12
+   -2.105289163948394e-11
+    8.149214332492391e-11
+ 4.16e+10    
+    8.161967807877108e-11
+   -2.105491373816473e-11
+    8.386878444187887e-11
+   -1.737968158849037e-12
+   -1.018946172859685e-11
+    8.389146457771995e-11
+   -1.074733604513114e-12
+   -1.733397836114644e-12
+   -2.105674560302889e-11
+    8.148772266684189e-11
+ 4.17e+10    
+    8.161520704723978e-11
+   -2.105878262945628e-11
+    8.386896666806932e-11
+   -1.740519414220995e-12
+   -1.019249756906841e-11
+    8.389164023280281e-11
+   -1.074273935867357e-12
+    -1.73595314980408e-12
+   -2.106061062689769e-11
+    8.148328229486038e-11
+ 4.18e+10    
+    8.161071609052372e-11
+   -2.106266250204618e-11
+    8.386914405624099e-11
+   -1.743060316362151e-12
+   -1.019554312099205e-11
+    8.389181104621053e-11
+   -1.073791534695543e-12
+   -1.738498184305805e-12
+   -2.106448666086725e-11
+    8.147882214299713e-11
+ 4.19e+10    
+    8.160620514273804e-11
+   -2.106655330523181e-11
+    8.386931654018337e-11
+   -1.745590805954107e-12
+   -1.019859837115977e-11
+    8.389197695202344e-11
+   -1.073286418531514e-12
+   -1.741032880340813e-12
+   -2.106837365453184e-11
+    8.147434214570784e-11
+ 4.2e+10     
+    8.160167413843169e-11
+   -2.107045498812475e-11
+    8.386948405386643e-11
+   -1.748110823750325e-12
+   -1.020166330654402e-11
+    8.389213788450893e-11
+    -1.07275860524561e-12
+   -1.743557178701094e-12
+   -2.107227155730228e-11
+    8.146984223788333e-11
+ 4.21e+10    
+    8.159712301258515e-11
+   -2.107436749965018e-11
+    8.386964653143915e-11
+   -1.750620310578714e-12
+   -1.020473791429731e-11
+    8.389229377811846e-11
+   -1.072208113046819e-12
+   -1.746071020252137e-12
+   -2.107618031840467e-11
+    8.146532235484613e-11
+ 4.22e+10    
+    8.159255170060738e-11
+   -2.107829078854577e-11
+    8.386980390722728e-11
+   -1.753119207344169e-12
+   -1.020782218175178e-11
+    8.389244456748685e-11
+   -1.071634960484925e-12
+   -1.748574345935498e-12
+   -2.108009988687978e-11
+    8.146078243234808e-11
+ 4.23e+10    
+    8.158796013833329e-11
+   -2.108222480336099e-11
+    8.386995611573179e-11
+   -1.755607455031142e-12
+   -1.021091609641873e-11
+    8.389259018742968e-11
+   -1.071039166452754e-12
+    -1.75106709677135e-12
+   -2.108403021158195e-11
+     8.14562224065677e-11
+ 4.24e+10    
+    8.158334826202031e-11
+     -2.1086169492456e-11
+    8.387010309162718e-11
+   -1.758084994706157e-12
+   -1.021401964598825e-11
+    8.389273057294106e-11
+   -1.070420750188417e-12
+   -1.753549213861008e-12
+   -2.108797124117818e-11
+    8.145164221410671e-11
+ 4.25e+10    
+    8.157871600834708e-11
+   -2.109012480400104e-11
+    8.387024476975942e-11
+    -1.76055176752043e-12
+   -1.021713281832862e-11
+    8.389286565919279e-11
+   -1.069779731277654e-12
+   -1.756020638389483e-12
+   -2.109192292414736e-11
+    8.144704179198818e-11
+ 4.26e+10    
+    8.157406331440908e-11
+   -2.109409068597532e-11
+    8.387038108514471e-11
+   -1.763007714712329e-12
+   -1.022025560148585e-11
+     8.38929953815313e-11
+   -1.069116129656169e-12
+   -1.758481311628016e-12
+   -2.109588520877915e-11
+    8.144242107765298e-11
+ 4.27e+10    
+    8.156939011771736e-11
+   -2.109806708616617e-11
+    8.387051197296703e-11
+   -1.765452777609976e-12
+   -1.022338798368311e-11
+    8.389311967547669e-11
+   -1.068429965612053e-12
+   -1.760931174936597e-12
+   -2.109985804317317e-11
+    8.143778000895776e-11
+ 4.28e+10    
+    8.156469635619511e-11
+   -2.110205395216842e-11
+    8.387063736857761e-11
+   -1.767886897633766e-12
+   -1.022652995332025e-11
+    8.389323847672062e-11
+   -1.067721259788216e-12
+   -1.763370169766531e-12
+   -2.110384137523811e-11
+    8.143311852417196e-11
+ 4.29e+10    
+    8.155998196817577e-11
+   -2.110605123138324e-11
+    8.387075720749219e-11
+   -1.770310016298913e-12
+   -1.022968149897307e-11
+    8.389335172112424e-11
+   -1.066990033184886e-12
+   -1.765798237662949e-12
+   -2.110783515269064e-11
+    8.142843656197526e-11
+ 4.3e+10     
+    8.155524689239969e-11
+   -2.111005887101737e-11
+    8.387087142538983e-11
+   -1.772722075217972e-12
+   -1.023284260939285e-11
+    8.389345934471715e-11
+   -1.066236307162126e-12
+   -1.768215320267295e-12
+   -2.111183932305489e-11
+    8.142373406145505e-11
+ 4.31e+10    
+    8.155049106801234e-11
+    -2.11140768180823e-11
+    8.387097995811183e-11
+   -1.775123016103379e-12
+   -1.023601327350566e-11
+    8.389356128369485e-11
+   -1.065460103442396e-12
+    -1.77062135931991e-12
+    -2.11158538336611e-11
+    8.141901096210379e-11
+ 4.32e+10    
+    8.154571443456138e-11
+   -2.111810501939339e-11
+    8.387108274165899e-11
+   -1.777512780769959e-12
+   -1.023919348041168e-11
+    8.389365747441762e-11
+   -1.064661444113165e-12
+   -1.773016296662491e-12
+     -2.1119878631645e-11
+    8.141426720381666e-11
+ 4.33e+10    
+    8.154091693199449e-11
+   -2.112214342156897e-11
+    8.387117971219113e-11
+   -1.779891311137462e-12
+   -1.024238321938458e-11
+    8.389374785340846e-11
+   -1.063840351629527e-12
+   -1.775400074240624e-12
+   -2.112391366394686e-11
+    8.140950272688896e-11
+ 4.34e+10    
+    8.153609850065678e-11
+    -2.11261919710296e-11
+    8.387127080602512e-11
+   -1.782258549233072e-12
+   -1.024558247987083e-11
+    8.389383235735186e-11
+   -1.062996848816886e-12
+   -1.777772634106291e-12
+   -2.112795887731063e-11
+    8.140471747201362e-11
+ 4.35e+10    
+    8.153125908128855e-11
+   -2.113025061399718e-11
+    8.387135595963371e-11
+    -1.78461443719389e-12
+   -1.024879125148897e-11
+    8.389391092309173e-11
+   -1.062130958873644e-12
+   -1.780133918420358e-12
+   -2.113201421828292e-11
+    8.139991138027871e-11
+ 4.36e+10    
+    8.152639861502257e-11
+   -2.113431929649398e-11
+    8.387143510964297e-11
+   -1.786958917269498e-12
+   -1.025200952402881e-11
+    8.389398348763005e-11
+   -1.061242705373937e-12
+   -1.782483869455045e-12
+   -2.113607963321236e-11
+     8.13950843931652e-11
+ 4.37e+10    
+    8.152151704338227e-11
+   -2.113839796434196e-11
+    8.387150819283211e-11
+   -1.789291931824381e-12
+   -1.025523728745078e-11
+    8.389404998812538e-11
+   -1.060332112270394e-12
+   -1.784822429596456e-12
+   -2.114015506824855e-11
+    8.139023645254454e-11
+ 4.38e+10    
+     8.15166143082789e-11
+   -2.114248656316195e-11
+    8.387157514613156e-11
+   -1.791613423340451e-12
+   -1.025847453188509e-11
+    8.389411036189043e-11
+   -1.059399203896931e-12
+   -1.787149541347022e-12
+   -2.114424046934113e-11
+    8.138536750067614e-11
+ 4.39e+10    
+    8.151169035200961e-11
+   -2.114658503837279e-11
+    8.387163590662129e-11
+    -1.79392333441955e-12
+   -1.026172124763099e-11
+    8.389416454639207e-11
+   -1.058444004971552e-12
+   -1.789465147327997e-12
+    -2.11483357822393e-11
+    8.138047748020547e-11
+ 4.4e+10     
+    8.150674511725527e-11
+   -2.115069333519041e-11
+    8.387169041152974e-11
+   -1.796221607785886e-12
+   -1.026497742515588e-11
+    8.389421247924823e-11
+   -1.057466540599207e-12
+    -1.79176919028189e-12
+   -2.115244095249042e-11
+    8.137556633416099e-11
+ 4.41e+10    
+     8.15017785470775e-11
+   -2.115481139862717e-11
+    8.387173859823197e-11
+   -1.798508186288531e-12
+   -1.026824305509455e-11
+     8.38942540982275e-11
+   -1.056466836274638e-12
+   -1.794061613074936e-12
+   -2.115655592543965e-11
+    8.137063400595264e-11
+ 4.42e+10    
+    8.149679058491745e-11
+   -2.115893917349102e-11
+      8.3871780404249e-11
+   -1.800783012903852e-12
+    -1.02715181282483e-11
+    8.389428934124713e-11
+   -1.055444917885286e-12
+   -1.796342358699565e-12
+   -2.116068064622884e-11
+    8.136568043936921e-11
+ 4.43e+10    
+    8.149178117459289e-11
+    -2.11630766043846e-11
+    8.387181576724579e-11
+   -1.803046030737999e-12
+   -1.027480263558406e-11
+    8.389431814637154e-11
+   -1.054400811714188e-12
+   -1.798611370276815e-12
+    -2.11648150597958e-11
+    8.136070557857614e-11
+ 4.44e+10    
+    8.148675026029644e-11
+   -2.116722363570466e-11
+    8.387184462503016e-11
+   -1.805297183029323e-12
+   -1.027809656823354e-11
+    8.389434045181102e-11
+   -1.053334544442897e-12
+   -1.800868591058768e-12
+   -2.116895911087348e-11
+    8.135570936811346e-11
+ 4.45e+10    
+    8.148169778659315e-11
+   -2.117138021164101e-11
+    8.387186691555152e-11
+   -1.807536413150822e-12
+   -1.028139991749228e-11
+    8.389435619592039e-11
+   -1.052246143154464e-12
+   -1.803113964430987e-12
+   -2.117311274398906e-11
+    8.135069175289336e-11
+ 4.46e+10    
+    8.147662369841855e-11
+   -2.117554627617599e-11
+    8.387188257689951e-11
+   -1.809763664612568e-12
+   -1.028471267481881e-11
+    8.389436531719737e-11
+   -1.051135635336356e-12
+   -1.805347433914914e-12
+   -2.117727590346322e-11
+    8.134565267819809e-11
+ 4.47e+10    
+    8.147152794107653e-11
+   -2.117972177308357e-11
+    8.387189154730272e-11
+   -1.811978881064136e-12
+   -1.028803483183361e-11
+    8.389436775428147e-11
+   -1.050003048883481e-12
+   -1.807568943170292e-12
+   -2.118144853340946e-11
+    8.134059208967818e-11
+ 4.48e+10    
+    8.146641046023701e-11
+   -2.118390664592854e-11
+    8.387189376512719e-11
+    -1.81418200629697e-12
+   -1.029136638031822e-11
+    8.389436344595223e-11
+   -1.048848412101163e-12
+   -1.809778435997559e-12
+   -2.118563057773299e-11
+    8.133550993334981e-11
+ 4.49e+10    
+    8.146127120193452e-11
+   -2.118810083806589e-11
+    8.387188916887552e-11
+   -1.816372984246855e-12
+   -1.029470731221422e-11
+    8.389435233112796e-11
+   -1.047671753708159e-12
+   -1.811975856340206e-12
+   -2.118982198013025e-11
+    8.133040615559294e-11
+ 4.5e+10     
+     8.14561101125651e-11
+      -2.119230429264e-11
+    8.387187769718562e-11
+   -1.818551758996231e-12
+   -1.029805761962242e-11
+    8.389433434886511e-11
+   -1.046473102839675e-12
+   -1.814161148287201e-12
+   -2.119402268408799e-11
+    8.132528070314915e-11
+ 4.51e+10    
+    8.145092713888552e-11
+   -2.119651695258393e-11
+    8.387185928882897e-11
+   -1.820718274776644e-12
+   -1.030141729480158e-11
+    8.389430943835574e-11
+   -1.045252489050417e-12
+    -1.81633425607531e-12
+   -2.119823263288254e-11
+    8.132013352311981e-11
+ 4.52e+10    
+    8.144572222801033e-11
+   -2.120073876061864e-11
+    8.387183388270993e-11
+   -1.822872475971049e-12
+   -1.030478633016756e-11
+    8.389427753892701e-11
+    -1.04400994231763e-12
+   -1.818495124091501e-12
+   -2.120245176957905e-11
+    8.131496456296385e-11
+ 4.53e+10    
+    8.144049532741026e-11
+   -2.120496965925231e-11
+     8.38718014178647e-11
+   -1.825014307116231e-12
+   -1.030816471829236e-11
+    8.389423859003999e-11
+   -1.042745493044147e-12
+   -1.820643696875257e-12
+   -2.120668003703069e-11
+    8.130977377049557e-11
+ 4.54e+10    
+    8.143524638491021e-11
+   -2.120920959077959e-11
+    8.387176183345927e-11
+   -1.827143712905119e-12
+   -1.031155245190287e-11
+     8.38941925312878e-11
+   -1.041459172061453e-12
+   -1.822779919120909e-12
+   -2.121091737787802e-11
+    8.130456109388307e-11
+ 4.55e+10    
+    8.142997534868722e-11
+   -2.121345849728096e-11
+    8.387171506878895e-11
+   -1.829260638189116e-12
+   -1.031494952387998e-11
+    8.389413930239488e-11
+   -1.040151010632768e-12
+   -1.824903735679981e-12
+   -2.121516373454818e-11
+    8.129932648164591e-11
+ 4.56e+10    
+    8.142468216726886e-11
+   -2.121771632062199e-11
+    8.387166106327743e-11
+   -1.831365027980479e-12
+   -1.031835592725742e-11
+    8.389407884321539e-11
+   -1.038821040456102e-12
+   -1.827015091563508e-12
+   -2.121941904925415e-11
+    8.129406988265326e-11
+ 4.57e+10    
+    8.141936678953085e-11
+   -2.122198300245274e-11
+     8.38715997564749e-11
+   -1.833456827454565e-12
+   -1.032177165522075e-11
+    8.389401109373241e-11
+    -1.03746929366735e-12
+   -1.829113931944306e-12
+   -2.122368326399414e-11
+    8.128879124612197e-11
+ 4.58e+10    
+    8.141402916469523e-11
+    -2.12262584842068e-11
+    8.387153108805737e-11
+   -1.835535981952196e-12
+   -1.032519670110614e-11
+    8.389393599405623e-11
+   -1.036095802843365e-12
+   -1.831200202159307e-12
+    -2.12279563205507e-11
+    8.128349052161454e-11
+ 4.59e+10    
+    8.140866924232907e-11
+   -2.123054270710112e-11
+     8.38714549978256e-11
+   -1.837602436981923e-12
+   -1.032863105839937e-11
+    8.389385348442341e-11
+   -1.034700601005044e-12
+   -1.833273847711792e-12
+   -2.123223816049029e-11
+    8.127816765903744e-11
+ 4.6e+10     
+    8.140328697234178e-11
+   -2.123483561213488e-11
+    8.387137142570378e-11
+   -1.839656138222321e-12
+   -1.033207472073465e-11
+    8.389376350519582e-11
+   -1.033283721620417e-12
+   -1.835334814273711e-12
+    -2.12365287251624e-11
+    8.127282260863899e-11
+ 4.61e+10    
+    8.139788230498391e-11
+   -2.123913714008911e-11
+    8.387128031173863e-11
+   -1.841697031524236e-12
+   -1.033552768189344e-11
+    8.389366599685902e-11
+   -1.031845198607729e-12
+   -1.837383047687895e-12
+    -2.12408279556988e-11
+    8.126745532100719e-11
+ 4.62e+10    
+    8.139245519084488e-11
+   -2.124344723152597e-11
+    8.387118159609828e-11
+   -1.843725062913089e-12
+   -1.033898993580342e-11
+    8.389356090002158e-11
+   -1.030385066338523e-12
+   -1.839418493970327e-12
+   -2.124513579301334e-11
+     8.12620657470689e-11
+ 4.63e+10    
+     8.13870055808513e-11
+    -2.12477658267881e-11
+    8.387107521907099e-11
+   -1.845740178591074e-12
+   -1.034246147653717e-11
+    8.389344815541339e-11
+   -1.028903359640718e-12
+   -1.841441099312351e-12
+   -2.124945217780064e-11
+    8.125665383808661e-11
+ 4.64e+10    
+    8.138153342626543e-11
+   -2.125209286599817e-11
+     8.38709611210647e-11
+   -1.847742324939427e-12
+   -1.034594229831116e-11
+    8.389332770388538e-11
+   -1.027400113801692e-12
+   -1.843450810082928e-12
+   -2.125377705053599e-11
+    8.125121954565766e-11
+ 4.65e+10    
+    8.137603867868305e-11
+   -2.125642828905804e-11
+    8.387083924260516e-11
+   -1.849731448520614e-12
+   -1.034943239548435e-11
+    8.389319948640723e-11
+   -1.025875364571352e-12
+   -1.845447572830811e-12
+    -2.12581103514744e-11
+    8.124576282171185e-11
+ 4.66e+10    
+    8.137052129003158e-11
+   -2.126077203564824e-11
+    8.387070952433555e-11
+   -1.851707496080586e-12
+   -1.035293176255724e-11
+    8.389306344406764e-11
+   -1.024329148165196e-12
+    -1.84743133428673e-12
+   -2.126245202065018e-11
+    8.124028361850981e-11
+ 4.67e+10    
+    8.136498121256883e-11
+   -2.126512404522752e-11
+    8.387057190701518e-11
+   -1.853670414550924e-12
+   -1.035644039417042e-11
+    8.389291951807195e-11
+   -1.022761501267374e-12
+   -1.849402041365625e-12
+   -2.126680199787619e-11
+     8.12347818886413e-11
+ 4.68e+10    
+    8.135941839888074e-11
+   -2.126948425703217e-11
+    8.387042633151876e-11
+   -1.855620151051048e-12
+   -1.035995828510353e-11
+    8.389276764974221e-11
+   -1.021172461033745e-12
+   -1.851359641168763e-12
+   -2.127116022274335e-11
+    8.122925758502323e-11
+ 4.69e+10    
+    8.135383280187993e-11
+    -2.12738526100754e-11
+    8.387027273883499e-11
+   -1.857556652890413e-12
+   -1.036348543027393e-11
+    8.389260778051526e-11
+   -1.019562065094905e-12
+   -1.853304080985903e-12
+   -2.127552663461995e-11
+    8.122371066089792e-11
+ 4.7e+10     
+    8.134822437480393e-11
+   -2.127822904314691e-11
+    8.387011107006581e-11
+   -1.859479867570596e-12
+   -1.036702182473547e-11
+    8.389243985194208e-11
+   -1.017930351559241e-12
+   -1.855235308297465e-12
+    -2.12799011726512e-11
+    8.121814106983159e-11
+ 4.71e+10    
+    8.134259307121333e-11
+   -2.128261349481227e-11
+     8.38699412664257e-11
+   -1.861389742787493e-12
+   -1.037056746367729e-11
+    8.389226380568687e-11
+   -1.016277359015924e-12
+   -1.857153270776632e-12
+   -2.128428377575858e-11
+    8.121254876571227e-11
+ 4.72e+10    
+    8.133693884499006e-11
+   -2.128700590341245e-11
+    8.386976326924004e-11
+   -1.863286226433453e-12
+   -1.037412234242242e-11
+    8.389207958352576e-11
+   -1.014603126537931e-12
+   -1.859057916291467e-12
+   -2.128867438263929e-11
+    8.120693370274825e-11
+ 4.73e+10    
+    8.133126165033626e-11
+    -2.12914062070633e-11
+    8.386957701994522e-11
+    -1.86516926659936e-12
+   -1.037768645642675e-11
+    8.389188712734584e-11
+   -1.012907693685045e-12
+   -1.860949192907023e-12
+   -2.129307293176579e-11
+    8.120129583546636e-11
+ 4.74e+10    
+    8.132556144177161e-11
+   -2.129581434365494e-11
+    8.386938246008651e-11
+   -1.867038811576739e-12
+   -1.038125980127746e-11
+    8.389168637914449e-11
+   -1.011191100506818e-12
+   -1.862827048887432e-12
+   -2.129747936138512e-11
+    8.119563511871007e-11
+ 4.75e+10    
+    8.131983817413251e-11
+   -2.130023025085144e-11
+    8.386917953131787e-11
+   -1.868894809859872e-12
+   -1.038484237269195e-11
+    8.389147728102811e-11
+   -1.009453387545544e-12
+   -1.864691432697963e-12
+   -2.130189360951867e-11
+    8.118995150763827e-11
+ 4.76e+10    
+    8.131409180257003e-11
+   -2.130465386609018e-11
+     8.38689681754009e-11
+   -1.870737210147842e-12
+    -1.03884341665164e-11
+    8.389125977521078e-11
+   -1.007694595839214e-12
+   -1.866542293007089e-12
+   -2.130631561396121e-11
+    8.118424495772267e-11
+ 4.77e+10    
+    8.130832228254821e-11
+   -2.130908512658147e-11
+    8.386874833420387e-11
+   -1.872565961346609e-12
+   -1.039203517872456e-11
+    8.389103380401436e-11
+   -1.005914766924426e-12
+   -1.868379578688542e-12
+   -2.131074531228098e-11
+    8.117851542474745e-11
+ 4.78e+10    
+     8.13025295698429e-11
+   -2.131352396930813e-11
+      8.3868519949701e-11
+    -1.87438101257105e-12
+   -1.039564540541637e-11
+    8.389079930986661e-11
+   -1.004113942839314e-12
+   -1.870203238823314e-12
+   -2.131518264181874e-11
+    8.117276286480613e-11
+ 4.79e+10    
+    8.129671362053936e-11
+   -2.131797033102487e-11
+     8.38682829639714e-11
+    -1.87618231314699e-12
+   -1.039926484281666e-11
+    8.389055623530037e-11
+   -1.002292166126426e-12
+   -1.872013222701732e-12
+    -2.13196275396875e-11
+    8.116698723430104e-11
+ 4.8e+10     
+    8.129087439103132e-11
+    -2.13224241482581e-11
+    8.386803731919796e-11
+   -1.877969812613205e-12
+    -1.04028934872738e-11
+    8.389030452295324e-11
+   -1.000449479835604e-12
+   -1.873809479825372e-12
+   -2.132407994277211e-11
+    8.116118848994111e-11
+ 4.81e+10    
+    8.128501183801897e-11
+   -2.132688535730531e-11
+    8.386778295766728e-11
+   -1.879743460723443e-12
+    -1.04065313352584e-11
+    8.389004411556598e-11
+   -9.985859275268285e-13
+   -1.875591959909128e-12
+   -2.132853978772874e-11
+    8.115536658874052e-11
+ 4.82e+10    
+    8.127912591850756e-11
+   -2.133135389423476e-11
+    8.386751982176789e-11
+   -1.881503207448403e-12
+   -1.041017838336187e-11
+    8.388977495598182e-11
+   -9.967015532730435e-13
+   -1.877360612883132e-12
+   -2.133300701098439e-11
+    8.114952148801653e-11
+ 4.83e+10    
+    8.127321658980573e-11
+   -2.133582969488508e-11
+    8.386724785398995e-11
+   -1.883249002977715e-12
+   -1.041383462829514e-11
+    8.388949698714587e-11
+   -9.947964016629514e-13
+   -1.879115388894745e-12
+   -2.133748154873668e-11
+    8.114365314538864e-11
+ 4.84e+10    
+    8.126728380952399e-11
+   -2.134031269486489e-11
+    8.386696699692439e-11
+   -1.884980797721859e-12
+   -1.041750006688731e-11
+    8.388921015210372e-11
+   -9.928705178038157e-13
+    -1.88085623831046e-12
+   -2.134196333695326e-11
+    8.113776151877641e-11
+ 4.85e+10    
+    8.126132753557271e-11
+   -2.134480282955228e-11
+    8.386667719326173e-11
+   -1.886698542314171e-12
+   -1.042117469608421e-11
+    8.388891439400087e-11
+   -9.909239473241748e-13
+   -1.882583111717883e-12
+   -2.134645231137144e-11
+    8.113184656639788e-11
+ 4.86e+10    
+    8.125534772616165e-11
+    -2.13493000340948e-11
+    8.386637838579186e-11
+   -1.888402187612706e-12
+   -1.042485851294706e-11
+    8.388860965608217e-11
+   -9.889567363766047e-13
+   -1.884295959927585e-12
+   -2.135094840749799e-11
+    8.112590824676833e-11
+ 4.87e+10    
+    8.124934433979689e-11
+   -2.135380424340875e-11
+    8.386607051740252e-11
+   -1.890091684702185e-12
+   -1.042855151465109e-11
+    8.388829588169024e-11
+   -9.869689316403923e-13
+    -1.88599473397505e-12
+   -2.135545156060854e-11
+    8.111994651869832e-11
+ 4.88e+10    
+    8.124331733528054e-11
+   -2.135831539217906e-11
+     8.38657535310792e-11
+    -1.89176698489588e-12
+   -1.043225369848414e-11
+    8.388797301426525e-11
+   -9.849605803242106e-13
+    -1.88767938512252e-12
+   -2.135996170574748e-11
+    8.111396134129251e-11
+ 4.89e+10    
+    8.123726667170843e-11
+   -2.136283341485888e-11
+    8.386542736990379e-11
+   -1.893428039737506e-12
+   -1.043596506184528e-11
+    8.388764099734371e-11
+   -9.829317301687634e-13
+   -1.889349864860887e-12
+   -2.136447877772728e-11
+    8.110795267394735e-11
+ 4.9e+10     
+    8.123119230846898e-11
+   -2.136735824566937e-11
+    8.386509197705419e-11
+   -1.895074801003058e-12
+   -1.043968560224337e-11
+     8.38872997745578e-11
+   -9.808824294493847e-13
+   -1.891006124911533e-12
+   -2.136900271112852e-11
+    8.110192047635037e-11
+ 4.91e+10    
+    8.122509420524151e-11
+   -2.137188981859931e-11
+    8.386474729580314e-11
+   -1.896707220702694e-12
+   -1.044341531729566e-11
+    8.388694928963469e-11
+   -9.788127269786343e-13
+   -1.892648117228157e-12
+   -2.137353344029947e-11
+    8.109586470847813e-11
+ 4.92e+10    
+    8.121897232199457e-11
+   -2.137642806740487e-11
+    8.386439326951789e-11
+   -1.898325251082552e-12
+   -1.044715420472644e-11
+    8.388658948639552e-11
+   -9.767226721088188e-13
+   -1.894275793998609e-12
+   -2.137807089935568e-11
+    8.108978533059482e-11
+ 4.93e+10    
+    8.121282661898482e-11
+   -2.138097292560938e-11
+    8.386402984165921e-11
+   -1.899928844626563e-12
+   -1.045090226236554e-11
+    8.388622030875458e-11
+    -9.74612314734525e-13
+   -1.895889107646699e-12
+   -2.138261502217981e-11
+    8.108368230325046e-11
+ 4.94e+10    
+    8.120665705675494e-11
+   -2.138552432650296e-11
+     8.38636569557806e-11
+   -1.901517954058259e-12
+   -1.045465948814695e-11
+    8.388584170071885e-11
+   -9.724817052950825e-13
+   -1.897488010833961e-12
+   -2.138716574242137e-11
+    8.107755558727978e-11
+ 4.95e+10    
+    8.120046359613273e-11
+   -2.139008220314246e-11
+    8.386327455552757e-11
+   -1.903092532342577e-12
+   -1.045842588010733e-11
+    8.388545360638654e-11
+   -9.703308947770274e-13
+    -1.89907245646146e-12
+   -2.139172299349635e-11
+    8.107140514380039e-11
+ 4.96e+10    
+    8.119424619822921e-11
+   -2.139464648835107e-11
+    8.386288258463703e-11
+   -1.904652532687588e-12
+    -1.04622014363847e-11
+    8.388505596994743e-11
+   -9.681599347164909e-13
+   -1.900642397671502e-12
+   -2.139628670858717e-11
+    8.106523093421118e-11
+ 4.97e+10    
+    8.118800482443699e-11
+   -2.139921711471822e-11
+    8.386248098693663e-11
+   -1.906197908546299e-12
+   -1.046598615521689e-11
+    8.388464873568086e-11
+    -9.65968877201574e-13
+   -1.902197787849444e-12
+   -2.140085682064232e-11
+    8.105903292019122e-11
+ 4.98e+10    
+    8.118173943642936e-11
+   -2.140379401459938e-11
+    8.386206970634359e-11
+   -1.907728613618375e-12
+   -1.046978003494013e-11
+     8.38842318479558e-11
+   -9.637577748746882e-13
+   -1.903738580625345e-12
+   -2.140543326237612e-11
+    8.105281106369763e-11
+ 4.99e+10    
+    8.117544999615821e-11
+   -2.140837712011577e-11
+    8.386164868686453e-11
+    -1.90924460185183e-12
+   -1.047358307398764e-11
+    8.388380525122997e-11
+   -9.615266809348466e-13
+   -1.905264729875725e-12
+   -2.141001596626868e-11
+    8.104656532696465e-11
+ 5e+10       
+     8.11691364658527e-11
+   -2.141296636315431e-11
+    8.386121787259451e-11
+   -1.910745827444786e-12
+   -1.047739527088808e-11
+    8.388336889004885e-11
+   -9.592756491399134e-13
+   -1.906776189725254e-12
+    -2.14146048645656e-11
+    8.104029567250183e-11
+ 5.01e+10    
+    8.116279880801808e-11
+   -2.141756167536746e-11
+    8.386077720771619e-11
+    -1.91223224484713e-12
+   -1.048121662426423e-11
+     8.38829227090451e-11
+   -9.570047338088355e-13
+   -1.908272914548407e-12
+   -2.141919988927771e-11
+    8.103400206309224e-11
+ 5.02e+10    
+     8.11564369854338e-11
+   -2.142216298817299e-11
+    8.386032663649941e-11
+   -1.913703808762206e-12
+   -1.048504713283144e-11
+     8.38824666529379e-11
+   -9.547139898237971e-13
+   -1.909754858971145e-12
+   -2.142380097218117e-11
+    8.102768446179181e-11
+ 5.03e+10    
+    8.115005096115239e-11
+   -2.142677023275399e-11
+    8.385986610330073e-11
+   -1.915160474148454e-12
+    -1.04888867953962e-11
+    8.388200066653224e-11
+   -9.524034726323702e-13
+   -1.911221977872568e-12
+   -2.142840804481721e-11
+     8.10213428319271e-11
+ 5.04e+10    
+    8.114364069849757e-11
+   -2.143138334005863e-11
+    8.385939555256174e-11
+    -1.91660219622108e-12
+   -1.049273561085467e-11
+    8.388152469471808e-11
+   -9.500732382495883e-13
+   -1.912674226386505e-12
+   -2.143302103849184e-11
+    8.101497713709375e-11
+ 5.05e+10    
+    8.113720616106316e-11
+   -2.143600224080011e-11
+    8.385891492880972e-11
+   -1.918028930453661e-12
+   -1.049659357819121e-11
+    8.388103868246983e-11
+   -9.477233432600042e-13
+   -1.914111559903195e-12
+   -2.143763988427599e-11
+    8.100858734115573e-11
+ 5.06e+10    
+    8.113074731271144e-11
+   -2.144062686545663e-11
+    8.385842417665608e-11
+   -1.919440632579758e-12
+   -1.050046069647693e-11
+    8.388054257484541e-11
+    -9.45353844819692e-13
+   -1.915533934070816e-12
+   -2.144226451300533e-11
+    8.100217340824318e-11
+ 5.07e+10    
+    8.112426411757201e-11
+   -2.144525714427129e-11
+    8.385792324079598e-11
+   -1.920837258594525e-12
+   -1.050433696486818e-11
+    8.388003631698585e-11
+   -9.429648006581985e-13
+   -1.916941304797092e-12
+    -2.14468948552801e-11
+      8.0995735302751e-11
+ 5.08e+10    
+    8.111775654003945e-11
+   -2.144989300725195e-11
+    8.385741206600777e-11
+   -1.922218764756261e-12
+   -1.050822238260509e-11
+    8.387951985411444e-11
+   -9.405562690804581e-13
+   -1.918333628250901e-12
+   -2.145153084146516e-11
+    8.098927298933785e-11
+ 5.09e+10    
+    8.111122454477315e-11
+   -2.145453438417139e-11
+     8.38568905971523e-11
+   -1.923585107588001e-12
+   -1.051211694901014e-11
+    8.387899313153612e-11
+   -9.381283089686565e-13
+   -1.919710860863765e-12
+   -2.145617240168986e-11
+    8.098278643292413e-11
+ 5.1e+10     
+    8.110466809669491e-11
+   -2.145918120456706e-11
+     8.38563587791719e-11
+   -1.924936243879045e-12
+   -1.051602066348659e-11
+    8.387845609463692e-11
+   -9.356809797840549e-13
+   -1.921072959331389e-12
+   -2.146081946584814e-11
+    8.097627559869092e-11
+ 5.11e+10    
+    8.109808716098765e-11
+   -2.146383339774128e-11
+    8.385581655709067e-11
+   -1.926272130686472e-12
+   -1.051993352551711e-11
+    8.387790868888304e-11
+   -9.332143415687422e-13
+   -1.922419880615225e-12
+   -2.146547196359827e-11
+    8.096974045207819e-11
+ 5.12e+10    
+     8.10914817030942e-11
+   -2.146849089276102e-11
+    8.385526387601276e-11
+   -1.927592725336698e-12
+   -1.052385553466215e-11
+    8.387735085982047e-11
+   -9.307284549473752e-13
+   -1.923751581943928e-12
+   -2.147012982436305e-11
+    8.096318095878351e-11
+ 5.13e+10    
+    8.108485168871599e-11
+   -2.147315361845819e-11
+    8.385470068112264e-11
+   -1.928897985426915e-12
+   -1.052778669055862e-11
+    8.387678255307427e-11
+   -9.282233811288421e-13
+   -1.925068020814851e-12
+   -2.147479297732973e-11
+    8.095659708476066e-11
+ 5.14e+10    
+    8.107819708381086e-11
+   -2.147782150342945e-11
+    8.385412691768401e-11
+   -1.930187868826605e-12
+   -1.053172699291829e-11
+    8.387620371434791e-11
+   -9.256991819078749e-13
+   -1.926369154995531e-12
+   -2.147946135145011e-11
+    8.094998879621797e-11
+ 5.15e+10    
+    8.107151785459276e-11
+   -2.148249447603636e-11
+    8.385354253103942e-11
+   -1.931462333679024e-12
+   -1.053567644152632e-11
+    8.387561428942257e-11
+   -9.231559196666225e-13
+   -1.927654942525128e-12
+   -2.148413487544039e-11
+    8.094335605961702e-11
+ 5.16e+10    
+    8.106481396752921e-11
+   -2.148717246440545e-11
+    8.385294746660963e-11
+   -1.932721338402599e-12
+   -1.053963503623983e-11
+    8.387501422415689e-11
+   -9.205936573761801e-13
+   -1.928925341715859e-12
+   -2.148881347778155e-11
+    8.093669884167137e-11
+ 5.17e+10    
+    8.105808538934067e-11
+   -2.149185539642827e-11
+    8.385234166989272e-11
+    -1.93396484169239e-12
+   -1.054360277698635e-11
+    8.387440346448577e-11
+   -9.180124585980403e-13
+   -1.930180311154419e-12
+     -2.1493497086719e-11
+    8.093001710934454e-11
+ 5.18e+10    
+    8.105133208699863e-11
+   -2.149654319976149e-11
+    8.385172508646405e-11
+   -1.935192802521515e-12
+   -1.054757966376231e-11
+     8.38737819564203e-11
+   -9.154123874855009e-13
+   -1.931419809703401e-12
+   -2.149818563026307e-11
+    8.092331082984915e-11
+ 5.19e+10    
+     8.10445540277244e-11
+     -2.1501235801827e-11
+    8.385109766197547e-11
+     -1.9364051801425e-12
+   -1.055156569663166e-11
+    8.387314964604679e-11
+   -9.127935087850473e-13
+   -1.932643796502661e-12
+    -2.15028790361888e-11
+    8.091657997064525e-11
+ 5.2e+10     
+    8.103775117898785e-11
+   -2.150593312981215e-11
+    8.385045934215442e-11
+   -1.937601934088733e-12
+   -1.055556087572425e-11
+    8.387250647952659e-11
+   -9.101558878376204e-13
+   -1.933852230970704e-12
+   -2.150757723203625e-11
+    8.090982449943891e-11
+ 5.21e+10    
+    8.103092350850542e-11
+   -2.151063511066969e-11
+    8.384981007280388e-11
+   -1.938783024175757e-12
+   -1.055956520123442e-11
+     8.38718524030951e-11
+      -9.074995905799e-13
+   -1.935045072806036e-12
+   -2.151228014511059e-11
+    8.090304438418066e-11
+ 5.22e+10    
+    8.102407098423935e-11
+   -2.151534167111805e-11
+    8.384914979980142e-11
+   -1.939948410502681e-12
+   -1.056357867341947e-11
+    8.387118736306141e-11
+   -9.048246835454671e-13
+   -1.936222281988505e-12
+   -2.151698770248214e-11
+    8.089623959306431e-11
+ 5.23e+10    
+    8.101719357439591e-11
+    -2.15200527376416e-11
+    8.384847846909902e-11
+   -1.941098053453469e-12
+   -1.056760129259818e-11
+    8.387051130580767e-11
+   -9.021312338659558e-13
+   -1.937383818780635e-12
+   -2.152169983098662e-11
+    8.088941009452517e-11
+ 5.24e+10    
+    8.101029124742404e-11
+   -2.152476823649056e-11
+    8.384779602672203e-11
+   -1.942231913698293e-12
+    -1.05716330591493e-11
+    8.386982417778845e-11
+   -8.994193092721306e-13
+   -1.938529643728909e-12
+   -2.152641645722534e-11
+    8.088255585723913e-11
+ 5.25e+10    
+    8.100336397201403e-11
+    -2.15294880936815e-11
+    8.384710241876925e-11
+   -1.943349952194804e-12
+   -1.057567397351013e-11
+    8.386912592553048e-11
+   -8.966889780949003e-13
+   -1.939659717665087e-12
+   -2.153113750756538e-11
+    8.087567685012073e-11
+ 5.26e+10    
+    8.099641171709593e-11
+   -2.153421223499743e-11
+    8.384639759141193e-11
+    -1.94445213018943e-12
+   -1.057972403617491e-11
+    8.386841649563177e-11
+    -8.93940309266283e-13
+   -1.940774001707464e-12
+   -2.153586290813973e-11
+    8.086877304232189e-11
+ 5.27e+10    
+    8.098943445183836e-11
+   -2.153894058598799e-11
+    8.384568149089322e-11
+    -1.94553840921866e-12
+   -1.058378324769342e-11
+    8.386769583476123e-11
+   -8.911733723203087e-13
+    -1.94187245726214e-12
+    -2.15405925848476e-11
+    8.086184440323069e-11
+ 5.28e+10    
+    8.098243214564696e-11
+   -2.154367307196983e-11
+    8.384495406352819e-11
+    -1.94660875111026e-12
+   -1.058785160866951e-11
+    8.386696388965806e-11
+   -8.883882373938689e-13
+   -1.942955046024259e-12
+   -2.154532646335461e-11
+    8.085489090246968e-11
+ 5.29e+10    
+    8.097540476816285e-11
+   -2.154840961802662e-11
+    8.384421525570262e-11
+   -1.947663117984554e-12
+   -1.059192911975947e-11
+    8.386622060713128e-11
+    -8.85584975227483e-13
+    -1.94402172997924e-12
+   -2.155006446909303e-11
+    8.084791250989464e-11
+ 5.3e+10     
+    8.096835228926148e-11
+   -2.155315014900955e-11
+    8.384346501387277e-11
+   -1.948701472255614e-12
+   -1.059601578167069e-11
+    8.386546593405924e-11
+   -8.827636571660416e-13
+   -1.945072471403983e-12
+   -2.155480652726216e-11
+    8.084090919559311e-11
+ 5.31e+10    
+    8.096127467905135e-11
+   -2.155789458953777e-11
+    8.384270328456532e-11
+   -1.949723776632466e-12
+   -1.060011159516013e-11
+    8.386469981738912e-11
+   -8.799243551594497e-13
+   -1.946107232868086e-12
+   -2.155955256282844e-11
+    8.083388092988285e-11
+ 5.32e+10    
+    8.095417190787205e-11
+   -2.156264286399824e-11
+    8.384193001437621e-11
+   -1.950729994120305e-12
+    -1.06042165610328e-11
+    8.386392220413609e-11
+   -8.770671417632311e-13
+   -1.947125977234988e-12
+   -2.156430250052588e-11
+    8.082682768331073e-11
+ 5.33e+10    
+    8.094704394629325e-11
+   -2.156739489654646e-11
+     8.38411451499702e-11
+   -1.951720088021641e-12
+   -1.060833068014029e-11
+    8.386313304138338e-11
+   -8.741920901390711e-13
+   -1.948128667663169e-12
+    -2.15690562648563e-11
+    8.081974942665084e-11
+ 5.34e+10    
+     8.09398907651135e-11
+   -2.157215061110669e-11
+    8.384034863808126e-11
+   -1.952694021937459e-12
+   -1.061245395337933e-11
+    8.386233227628115e-11
+   -8.712992740552801e-13
+   -1.949115267607302e-12
+   -2.157381378008975e-11
+    8.081264613090377e-11
+ 5.35e+10    
+    8.093271233535823e-11
+    -2.15769099313721e-11
+    8.383954042551058e-11
+   -1.953651759768379e-12
+    -1.06165863816902e-11
+    8.386151985604659e-11
+   -8.683887678872128e-13
+   -1.950085740819342e-12
+   -2.157857497026477e-11
+    8.080551776729438e-11
+ 5.36e+10    
+    8.092550862827905e-11
+   -2.158167278080562e-11
+    8.383872045912774e-11
+   -1.954593265715765e-12
+    -1.06207279660554e-11
+      8.3860695727963e-11
+   -8.654606466176014e-13
+   -1.951040051349698e-12
+   -2.158333975918879e-11
+    8.079836430727111e-11
+ 5.37e+10    
+    8.091827961535162e-11
+   -2.158643908263976e-11
+    8.383788868586892e-11
+   -1.955518504282843e-12
+   -1.062487870749806e-11
+    8.385985983937953e-11
+   -8.625149858368479e-13
+   -1.951978163548304e-12
+   -2.158810807043854e-11
+     8.07911857225041e-11
+ 5.38e+10    
+    8.091102526827482e-11
+   -2.159120875987746e-11
+    8.383704505273716e-11
+   -1.956427440275779e-12
+   -1.062903860708048e-11
+    8.385901213771057e-11
+    -8.59551861743239e-13
+   -1.952900042065708e-12
+   -2.159287982736034e-11
+    8.078398198488403e-11
+ 5.39e+10    
+    8.090374555896916e-11
+   -2.159598173529226e-11
+    8.383618950680183e-11
+   -1.957320038804787e-12
+   -1.063320766590273e-11
+    8.385815257043556e-11
+    -8.56571351143089e-13
+   -1.953805651854172e-12
+   -2.159765495307068e-11
+    8.077675306652066e-11
+ 5.4e+10     
+    8.089644045957545e-11
+   -2.160075793142886e-11
+    8.383532199519781e-11
+   -1.958196265285171e-12
+   -1.063738588510106e-11
+    8.385728108509808e-11
+   -8.535735314508324e-13
+   -1.954694958168672e-12
+   -2.160243337045646e-11
+    8.076949893974136e-11
+ 5.41e+10    
+    8.088910994245323e-11
+   -2.160553727060351e-11
+    8.383444246512538e-11
+   -1.959056085438367e-12
+    -1.06415732658465e-11
+    8.385639762930553e-11
+   -8.505584806890433e-13
+   -1.955567926568009e-12
+   -2.160721500217556e-11
+    8.076221957708984e-11
+ 5.42e+10    
+    8.088175398017941e-11
+   -2.161031967490442e-11
+     8.38335508638498e-11
+   -1.959899465293005e-12
+   -1.064576980934344e-11
+    8.385550215072925e-11
+   -8.475262774883651e-13
+   -1.956424522915778e-12
+   -2.161199977065722e-11
+     8.07549149513245e-11
+ 5.43e+10    
+    8.087437254554715e-11
+   -2.161510506619248e-11
+    8.383264713870081e-11
+   -1.960726371185874e-12
+   -1.064997551682807e-11
+    8.385459459710308e-11
+   -8.444770010874381e-13
+   -1.957264713381406e-12
+   -2.161678759810265e-11
+    8.074758503541751e-11
+ 5.44e+10    
+    8.086696561156432e-11
+   -2.161989336610144e-11
+    8.383173123707197e-11
+   -1.961536769762993e-12
+   -1.065419038956697e-11
+    8.385367491622396e-11
+   -8.414107313326701e-13
+   -1.958088464441144e-12
+   -2.162157840648532e-11
+    8.074022980255276e-11
+ 5.45e+10    
+    8.085953315145164e-11
+   -2.162468449603854e-11
+    8.383080310642034e-11
+   -1.962330627980535e-12
+   -1.065841442885559e-11
+    8.385274305595038e-11
+   -8.383275486780086e-13
+    -1.95889574287905e-12
+   -2.162637211755154e-11
+    8.073284922612502e-11
+ 5.46e+10    
+    8.085207513864236e-11
+   -2.162947837718532e-11
+    8.382986269426658e-11
+   -1.963107913105822e-12
+   -1.066264763601699e-11
+    8.385179896420315e-11
+   -8.352275341846213e-13
+   -1.959686515787933e-12
+   -2.163116865282114e-11
+    8.072544327973829e-11
+ 5.47e+10    
+    8.084459154677962e-11
+   -2.163427493049758e-11
+    8.382890994819359e-11
+    -1.96386859271829e-12
+   -1.066689001240007e-11
+    8.385084258896399e-11
+   -8.321107695204957e-13
+   -1.960460750570344e-12
+   -2.163596793358776e-11
+    8.071801193720449e-11
+ 5.48e+10    
+    8.083708234971609e-11
+   -2.163907407670656e-11
+     8.38279448158471e-11
+   -1.964612634710417e-12
+   -1.067114155937839e-11
+    8.384987387827551e-11
+   -8.289773369599893e-13
+   -1.961218414939485e-12
+   -2.164076988091954e-11
+    8.071055517254202e-11
+ 5.49e+10    
+    8.082954752151202e-11
+    -2.16438757363191e-11
+    8.382696724493429e-11
+   -1.965340007288647e-12
+   -1.067540227834863e-11
+    8.384889278024113e-11
+    -8.25827319383301e-13
+   -1.961959476920089e-12
+   -2.164557441565967e-11
+    8.070307295997419e-11
+ 5.5e+10     
+    8.082198703643393e-11
+   -2.164867982961833e-11
+    8.382597718322435e-11
+   -1.966050678974306e-12
+   -1.067967217072911e-11
+    8.384789924302386e-11
+   -8.226608002758681e-13
+   -1.962683904849441e-12
+   -2.165038145842697e-11
+    8.069556527392839e-11
+ 5.51e+10    
+    8.081440086895337e-11
+   -2.165348627666438e-11
+    8.382497457854721e-11
+   -1.966744618604501e-12
+   -1.068395123795842e-11
+    8.384689321484676e-11
+   -8.194778637276958e-13
+   -1.963391667378142e-12
+   -2.165519092961649e-11
+    8.068803208903394e-11
+ 5.52e+10    
+    8.080678899374542e-11
+   -2.165829499729492e-11
+    8.382395937879382e-11
+   -1.967421795332991e-12
+   -1.068823948149389e-11
+    8.384587464399187e-11
+   -8.162785944326322e-13
+   -1.964082733471079e-12
+   -2.166000274940006e-11
+    8.068047338012142e-11
+ 5.53e+10    
+    8.079915138568741e-11
+   -2.166310591112583e-11
+    8.382293153191564e-11
+   -1.968082178631055e-12
+   -1.069253690281032e-11
+    8.384484347880032e-11
+   -8.130630776875453e-13
+   -1.964757072408227e-12
+   -2.166481683772709e-11
+    8.067288912222079e-11
+ 5.54e+10    
+    8.079148801985747e-11
+    -2.16679189375518e-11
+    8.382189098592362e-11
+   -1.968725738288361e-12
+   -1.069684350339834e-11
+     8.38437996676717e-11
+   -8.098313993914389e-13
+   -1.965414653785533e-12
+   -2.166963311432503e-11
+    8.066527929056017e-11
+ 5.55e+10    
+    8.078379887153299e-11
+   -2.167273399574703e-11
+    8.382083768888887e-11
+   -1.969352444413758e-12
+   -1.070115928476318e-11
+    8.384274315906349e-11
+   -8.065836460445231e-13
+   -1.966055447515721e-12
+   -2.167445149870014e-11
+    8.065764386056456e-11
+ 5.56e+10    
+    8.077608391618973e-11
+   -2.167755100466595e-11
+    8.381977158894154e-11
+   -1.969962267436172e-12
+   -1.070548424842311e-11
+    8.384167390149123e-11
+   -8.033199047471582e-13
+   -1.966679423829152e-12
+   -2.167927191013811e-11
+    8.064998280785432e-11
+ 5.57e+10    
+     8.07683431294999e-11
+   -2.168236988304395e-11
+    8.381869263427064e-11
+   -1.970555178105326e-12
+   -1.070981839590812e-11
+    8.384059184352763e-11
+   -8.000402631987836e-13
+   -1.967286553274578e-12
+   -2.168409426770483e-11
+    8.064229610824372e-11
+ 5.58e+10    
+    8.076057648733091e-11
+   -2.168719054939787e-11
+    8.381760077312382e-11
+   -1.971131147492601e-12
+   -1.071416172875846e-11
+    8.383949693380252e-11
+   -7.967448096967347e-13
+   -1.967876806719966e-12
+   -2.168891849024705e-11
+     8.06345837377399e-11
+ 5.59e+10    
+    8.075278396574415e-11
+   -2.169201292202706e-11
+    8.381649595380696e-11
+   -1.971690146991781e-12
+   -1.071851424852322e-11
+    8.383838912100231e-11
+   -7.934336331350078e-13
+    -1.96845015535328e-12
+   -2.169374449639303e-11
+      8.0626845672541e-11
+ 5.6e+10     
+    8.074496554099369e-11
+   -2.169683691901391e-11
+    8.381537812468379e-11
+   -1.972232148319841e-12
+   -1.072287595675895e-11
+    8.383726835386973e-11
+   -7.901068230029458e-13
+   -1.969006570683224e-12
+    -2.16985722045535e-11
+    8.061908188903536e-11
+ 5.61e+10    
+    8.073712118952469e-11
+   -2.170166245822469e-11
+    8.381424723417532e-11
+   -1.972757123517662e-12
+   -1.072724685502827e-11
+    8.383613458120337e-11
+   -7.867644693838519e-13
+   -1.969546024539978e-12
+   -2.170340153292214e-11
+    8.061129236379954e-11
+ 5.62e+10    
+    8.072925088797206e-11
+   -2.170648945731029e-11
+    8.381310323076019e-11
+   -1.973265044950801e-12
+   -1.073162694489848e-11
+    8.383498775185777e-11
+   -7.834066629535274e-13
+   -1.970068489075974e-12
+    -2.17082323994766e-11
+    8.060347707359741e-11
+ 5.63e+10    
+    8.072135461315929e-11
+   -2.171131783370717e-11
+    8.381194606297359e-11
+     -1.9737558853102e-12
+   -1.073601622794016e-11
+    8.383382781474233e-11
+   -7.800334949787403e-13
+   -1.970573936766593e-12
+   -2.171306472197914e-11
+     8.05956359953787e-11
+ 5.64e+10    
+    8.071343234209643e-11
+   -2.171614750463772e-11
+    8.381077567940709e-11
+   -1.974229617612902e-12
+   -1.074041470572571e-11
+    8.383265471882165e-11
+   -7.766450573156189e-13
+    -1.97106234041085e-12
+   -2.171789841797742e-11
+    8.058776910627723e-11
+ 5.65e+10    
+    8.070548405197981e-11
+   -2.172097838711173e-11
+    8.380959202870892e-11
+   -1.974686215202728e-12
+   -1.074482237982814e-11
+    8.383146841311488e-11
+   -7.732414424079697e-13
+    -1.97153367313215e-12
+   -2.172273340480543e-11
+    8.057987638361013e-11
+ 5.66e+10    
+    8.069750972018983e-11
+   -2.172581039792679e-11
+    8.380839505958278e-11
+   -1.975125651750982e-12
+   -1.074923925181953e-11
+    8.383026884669553e-11
+    -7.69822743285529e-13
+   -1.971987908378894e-12
+   -2.172756959958426e-11
+    8.057195780487612e-11
+ 5.67e+10    
+    8.068950932428963e-11
+   -2.173064345366919e-11
+    8.380718472078807e-11
+    -1.97554790125708e-12
+   -1.075366532326976e-11
+    8.382905596869107e-11
+   -7.663890535621326e-13
+   -1.972425019925191e-12
+   -2.173240691922298e-11
+    8.056401334775416e-11
+ 5.68e+10    
+    8.068148284202431e-11
+   -2.173547747071497e-11
+    8.380596096113967e-11
+   -1.975952938049266e-12
+   -1.075810059574509e-11
+    8.382782972828258e-11
+    -7.62940467433801e-13
+   -1.972844981871517e-12
+   -2.173724528041942e-11
+    8.055604299010228e-11
+ 5.69e+10    
+    8.067343025131885e-11
+   -2.174031236523062e-11
+     8.38047237295073e-11
+   -1.976340736785173e-12
+   -1.076254507080685e-11
+    8.382659007470468e-11
+   -7.594770796768019e-13
+   -1.973247768645328e-12
+   -2.174208459966117e-11
+    8.054804670995611e-11
+ 5.7e+10     
+    8.066535153027739e-11
+   -2.174514805317415e-11
+    8.380347297481528e-11
+    -1.97671127245253e-12
+   -1.076699875001008e-11
+      8.3825336957245e-11
+   -7.559989856455507e-13
+   -1.973633355001684e-12
+   -2.174692479322645e-11
+     8.05400244855273e-11
+ 5.71e+10    
+    8.065724665718134e-11
+   -2.174998445029581e-11
+    8.380220864604238e-11
+   -1.977064520369715e-12
+   -1.077146163490206e-11
+     8.38240703252439e-11
+   -7.525062812705191e-13
+   -1.974001716023907e-12
+   -2.175176577718488e-11
+    8.053197629520251e-11
+ 5.72e+10    
+    8.064911561048828e-11
+   -2.175482147213925e-11
+    8.380093069222152e-11
+   -1.977400456186367e-12
+   -1.077593372702118e-11
+    8.382279012809425e-11
+    -7.48999063056036e-13
+   -1.974352827124123e-12
+    -2.17566074673986e-11
+    8.052390211754194e-11
+ 5.73e+10    
+    8.064095836883078e-11
+   -2.175965903404229e-11
+    8.379963906243949e-11
+   -1.977719055884008e-12
+   -1.078041502789544e-11
+    8.382149631524124e-11
+   -7.454774280780027e-13
+   -1.974686664043894e-12
+   -2.176144977952317e-11
+    8.051580193127786e-11
+ 5.74e+10    
+     8.06327749110145e-11
+   -2.176449705113796e-11
+    8.379833370583677e-11
+   -1.978020295776567e-12
+    -1.07849055390412e-11
+    8.382018883618189e-11
+   -7.419414739815478e-13
+   -1.975003202854787e-12
+   -2.176629262900842e-11
+    8.050767571531353e-11
+ 5.75e+10    
+    8.062456521601731e-11
+   -2.176933543835543e-11
+    8.379701457160652e-11
+   -1.978304152510972e-12
+   -1.078940526196177e-11
+    8.381886764046511e-11
+   -7.383912989786234e-13
+   -1.975302419958882e-12
+   -2.177113593109957e-11
+    8.049952344872146e-11
+ 5.76e+10    
+    8.061632926298814e-11
+   -2.177417411042116e-11
+    8.379568160899581e-11
+   -1.978570603067702e-12
+   -1.079391419814621e-11
+    8.381753267769084e-11
+   -7.348270018454877e-13
+   -1.975584292089419e-12
+   -2.177597960083806e-11
+    8.049134511074239e-11
+ 5.77e+10    
+    8.060806703124487e-11
+   -2.177901298185966e-11
+    8.379433476730393e-11
+   -1.978819624761282e-12
+    -1.07984323490679e-11
+     8.38161838975105e-11
+   -7.312486819201479e-13
+   -1.975848796311252e-12
+   -2.178082355306274e-11
+    8.048314068078385e-11
+ 5.78e+10    
+    8.059977850027353e-11
+   -2.178385196699472e-11
+    8.379297399588264e-11
+   -1.979051195240856e-12
+   -1.080295971618327e-11
+    8.381482124962623e-11
+   -7.276564390997174e-13
+   -1.976095910021413e-12
+   -2.178566770241071e-11
+    8.047491013841877e-11
+ 5.79e+10    
+    8.059146364972691e-11
+   -2.178869097995034e-11
+    8.379159924413639e-11
+    -1.97926529249066e-12
+   -1.080749630093057e-11
+    8.381344468379094e-11
+   -7.240503738376889e-13
+   -1.976325610949592e-12
+   -2.179051196331847e-11
+    8.046665346338414e-11
+ 5.8e+10     
+    8.058312245942304e-11
+   -2.179352993465183e-11
+    8.379021046152126e-11
+   -1.979461894830543e-12
+   -1.081204210472844e-11
+    8.381205414980781e-11
+   -7.204305871411551e-13
+   -1.976537877158687e-12
+   -2.179535625002297e-11
+    8.045837063557983e-11
+ 5.81e+10    
+    8.057475490934421e-11
+   -2.179836874482694e-11
+    8.378880759754546e-11
+    -1.97964098091642e-12
+   -1.081659712897475e-11
+    8.381064959753011e-11
+   -7.167971805679321e-13
+   -1.976732687045243e-12
+   -2.180020047656255e-11
+    8.045006163506702e-11
+ 5.82e+10    
+    8.056636097963504e-11
+   -2.180320732400673e-11
+    8.378739060176829e-11
+   -1.979802529740785e-12
+   -1.082116137504522e-11
+    8.380923097686136e-11
+   -7.131502562236271e-13
+   -1.976910019339948e-12
+   -2.180504455677818e-11
+    8.044172644206708e-11
+ 5.83e+10    
+    8.055794065060187e-11
+   -2.180804558552697e-11
+    8.378595942380092e-11
+   -1.979946520633136e-12
+   -1.082573484429217e-11
+    8.380779823775439e-11
+   -7.094899167586214e-13
+   -1.977069853108101e-12
+   -2.180988840431449e-11
+    8.043336503696013e-11
+ 5.84e+10    
+    8.054949390271064e-11
+     -2.1812883442529e-11
+    8.378451401330525e-11
+   -1.980072933260431e-12
+   -1.083031753804329e-11
+    8.380635133021147e-11
+   -7.058162653649813e-13
+   -1.977212167750045e-12
+   -2.181473193262078e-11
+     8.04249774002837e-11
+ 5.85e+10    
+    8.054102071658637e-11
+   -2.181772080796098e-11
+    8.378305431999425e-11
+   -1.980181747627544e-12
+   -1.083490945760032e-11
+    8.380489020428461e-11
+   -7.021294057733033e-13
+    -1.97733694300162e-12
+   -2.181957505495241e-11
+    8.041656351273164e-11
+ 5.86e+10    
+    8.053252107301118e-11
+   -2.182255759457908e-11
+    8.378158029363157e-11
+   -1.980272944077648e-12
+   -1.083951060423782e-11
+    8.380341481007433e-11
+   -6.984294422494704e-13
+   -1.977444158934595e-12
+   -2.182441768437157e-11
+    8.040812335515235e-11
+ 5.87e+10    
+    8.052399495292325e-11
+   -2.182739371494843e-11
+     8.37800918840313e-11
+   -1.980346503292662e-12
+   -1.084412097920192e-11
+     8.38019250977302e-11
+   -6.947164795913515e-13
+   -1.977533795957067e-12
+   -2.182925973374874e-11
+    8.039965690854765e-11
+ 5.88e+10    
+    8.051544233741561e-11
+   -2.183222908144457e-11
+     8.37785890410576e-11
+   -1.980402406293645e-12
+   -1.084874058370904e-11
+    8.380042101745032e-11
+   -6.909906231254232e-13
+   -1.977605834813859e-12
+   -2.183410111576376e-11
+    8.039116415407213e-11
+ 5.89e+10    
+    8.050686320773471e-11
+   -2.183706360625446e-11
+    8.377707171462512e-11
+   -1.980440634441168e-12
+   -1.085336941894469e-11
+    8.379890251948135e-11
+   -6.872519787033038e-13
+   -1.977660256586952e-12
+   -2.183894174290699e-11
+    8.038264507303067e-11
+ 5.9e+10     
+    8.049825754527886e-11
+   -2.184189720137772e-11
+    8.377553985469812e-11
+   -1.980461169435676e-12
+   -1.085800748606226e-11
+    8.379736955411804e-11
+   -6.835006526982403e-13
+   -1.977697042695831e-12
+   -2.184378152748046e-11
+    8.037409964687793e-11
+ 5.91e+10    
+    8.048962533159742e-11
+   -2.184672977862782e-11
+    8.377399341129055e-11
+   -1.980463993317904e-12
+   -1.086265478618171e-11
+    8.379582207170329e-11
+   -6.797367520015059e-13
+   -1.977716174897842e-12
+   -2.184862038159924e-11
+    8.036552785721694e-11
+ 5.92e+10    
+    8.048096654838889e-11
+   -2.185156124963339e-11
+    8.377243233446603e-11
+   -1.980449088469175e-12
+    -1.08673113203884e-11
+    8.379426002262761e-11
+   -6.759603840187196e-13
+   -1.977717635288603e-12
+   -2.185345821719246e-11
+    8.035692968579756e-11
+ 5.93e+10    
+    8.047228117750046e-11
+   -2.185639152583943e-11
+    8.377085657433726e-11
+   -1.980416437611787e-12
+   -1.087197708973193e-11
+    8.379268335732943e-11
+   -6.721716566661206e-13
+   -1.977701406302283e-12
+   -2.185829494600476e-11
+    8.034830511451541e-11
+ 5.94e+10    
+    8.046356920092572e-11
+    -2.18612205185085e-11
+    8.376926608106636e-11
+   -1.980366023809292e-12
+   -1.087665209522486e-11
+    8.379109202629474e-11
+   -6.683706783667339e-13
+   -1.977667470711991e-12
+   -2.186313047959743e-11
+    8.033965412541054e-11
+ 5.95e+10    
+    8.045483060080407e-11
+   -2.186604813872216e-11
+    8.376766080486445e-11
+   -1.980297830466849e-12
+   -1.088133633784153e-11
+     8.37894859800565e-11
+   -6.645575580464981e-13
+     -1.9776158116301e-12
+    -2.18679647293496e-11
+    8.033097670066613e-11
+ 5.96e+10    
+    8.044606535941914e-11
+     -2.1870874297382e-11
+    8.376604069599122e-11
+   -1.980211841331542e-12
+   -1.088602981851685e-11
+    8.378786516919517e-11
+    -6.60732405130306e-13
+   -1.977546412508494e-12
+   -2.187279760645971e-11
+    8.032227282260694e-11
+ 5.97e+10    
+     8.04372734591975e-11
+   -2.187569890521121e-11
+    8.376440570475539e-11
+   -1.980108040492621e-12
+   -1.089073253814525e-11
+    8.378622954433824e-11
+   -6.568953295379668e-13
+   -1.977459257138962e-12
+   -2.187762902194682e-11
+    8.031354247369879e-11
+ 5.98e+10    
+    8.042845488270767e-11
+   -2.188052187275578e-11
+    8.376275578151392e-11
+   -1.979986412381852e-12
+   -1.089544449757927e-11
+    8.378457905615975e-11
+   -6.530464416801227e-13
+   -1.977354329653421e-12
+   -2.188245888665155e-11
+    8.030478563654627e-11
+ 5.99e+10    
+    8.041960961265834e-11
+   -2.188534311038578e-11
+    8.376109087667238e-11
+   -1.979846941773747e-12
+   -1.090016569762861e-11
+     8.37829136553808e-11
+   -6.491858524540589e-13
+   -1.977231614524243e-12
+   -2.188728711123791e-11
+    8.029600229389236e-11
+ 6e+10       
+    8.041073763189748e-11
+   -2.189016252829678e-11
+    8.375941094068433e-11
+   -1.979689613785834e-12
+   -1.090489613905885e-11
+    8.378123329276891e-11
+   -6.453136732394893e-13
+   -1.977091096564465e-12
+   -2.189211360619436e-11
+    8.028719242861648e-11
+ 6.01e+10    
+    8.040183892341101e-11
+   -2.189498003651119e-11
+    8.375771592405181e-11
+   -1.979514413878929e-12
+   -1.090963582259031e-11
+    8.377953791913803e-11
+   -6.414300158942244e-13
+   -1.976932760928137e-12
+   -2.189693828183515e-11
+    8.027835602373389e-11
+ 6.02e+10    
+    8.039291347032147e-11
+   -2.189979554487965e-11
+    8.375600577732437e-11
+   -1.979321327857356e-12
+   -1.091438474889694e-11
+    8.377782748534833e-11
+   -6.375349927498128e-13
+   -1.976756593110482e-12
+   -2.190176104830175e-11
+    8.026949306239382e-11
+ 6.03e+10    
+     8.03839612558868e-11
+   -2.190460896308238e-11
+    8.375428045109995e-11
+   -1.979110341869175e-12
+   -1.091914291860519e-11
+    8.377610194230642e-11
+   -6.336287166070818e-13
+   -1.976562578948195e-12
+   -2.190658181556432e-11
+     8.02606035278786e-11
+ 6.04e+10    
+    8.037498226349879e-11
+   -2.190942020063053e-11
+     8.37525398960237e-11
+   -1.978881442406419e-12
+   -1.092391033229278e-11
+    8.377436124096472e-11
+   -6.297113007316323e-13
+   -1.976350704619624e-12
+   -2.191140049342295e-11
+     8.02516874036022e-11
+ 6.05e+10    
+    8.036597647668249e-11
+    -2.19142291668678e-11
+    8.375078406278886e-11
+   -1.978634616305294e-12
+    -1.09286869904877e-11
+    8.377260533232169e-11
+   -6.257828588492415e-13
+   -1.976120956645054e-12
+   -2.191621699150915e-11
+    8.024274467310936e-11
+ 6.06e+10    
+    8.035694387909431e-11
+   -2.191903577097154e-11
+    8.374901290213575e-11
+   -1.978369850746384e-12
+   -1.093347289366703e-11
+    8.377083416742178e-11
+   -6.218435051412296e-13
+   -1.975873321886834e-12
+   -2.192103121928735e-11
+    8.023377532007394e-11
+ 6.07e+10    
+    8.034788445452113e-11
+   -2.192383992195459e-11
+    8.374722636485239e-11
+   -1.978087133254811e-12
+   -1.093826804225582e-11
+    8.376904769735478e-11
+   -6.178933542397356e-13
+   -1.975607787549636e-12
+   -2.192584308605604e-11
+    8.022477932829767e-11
+ 6.08e+10    
+    8.033879818687893e-11
+    -2.19286415286663e-11
+    8.374542440177401e-11
+   -1.977786451700467e-12
+   -1.094307243662601e-11
+    8.376724587325639e-11
+   -6.139325212229307e-13
+   -1.975324341180616e-12
+    -2.19306525009496e-11
+    8.021575668170935e-11
+ 6.09e+10    
+    8.032968506021158e-11
+   -2.193344049979434e-11
+    8.374360696378298e-11
+   -1.977467794298125e-12
+   -1.094788607709536e-11
+    8.376542864630789e-11
+   -6.099611216101667e-13
+   -1.975022970669591e-12
+   -2.193545937293957e-11
+    8.020670736436333e-11
+ 6.1e+10     
+    8.032054505868987e-11
+   -2.193823674386608e-11
+    8.374177400180894e-11
+   -1.977131149607638e-12
+   -1.095270896392632e-11
+    8.376359596773583e-11
+   -6.059792713570747e-13
+   -1.974703664249236e-12
+    -2.19402636108361e-11
+    8.019763136043843e-11
+ 6.11e+10    
+    8.031137816660972e-11
+      -2.194303016925e-11
+    8.373992546682849e-11
+   -1.976776506534057e-12
+   -1.095754109732501e-11
+    8.376174778881233e-11
+   -6.019870868505645e-13
+   -1.974366410495158e-12
+   -2.194506512328948e-11
+    8.018852865423633e-11
+ 6.12e+10    
+    8.030218436839146e-11
+   -2.194782068415722e-11
+    8.373806130986506e-11
+   -1.976403854327796e-12
+   -1.096238247744004e-11
+    8.375988406085446e-11
+   -5.979846849037866e-13
+   -1.974011198326177e-12
+    -2.19498638187917e-11
+    8.017939923018106e-11
+ 6.13e+10    
+    8.029296364857848e-11
+   -2.195260819664313e-11
+    8.373618148198916e-11
+   -1.976013182584722e-12
+    -1.09672331043616e-11
+     8.37580047352246e-11
+   -5.939721827510385e-13
+   -1.973638017004335e-12
+   -2.195465960567788e-11
+    8.017024307281743e-11
+ 6.14e+10    
+    8.028371599183591e-11
+    -2.19573926146088e-11
+    8.373428593431802e-11
+   -1.975604481246329e-12
+   -1.097209297812029e-11
+    8.375610976333062e-11
+   -5.899496980425583e-13
+   -1.973246856135101e-12
+   -2.195945239212781e-11
+    8.016106016680945e-11
+ 6.15e+10    
+    8.027444138294959e-11
+   -2.196217384580259e-11
+     8.37323746180156e-11
+   -1.975177740599779e-12
+   -1.097696209868614e-11
+    8.375419909662502e-11
+   -5.859173488393269e-13
+   -1.972837705667459e-12
+   -2.196424208616754e-11
+    8.015185049694003e-11
+ 6.16e+10    
+    8.026513980682503e-11
+   -2.196695179782172e-11
+    8.373044748429273e-11
+    -1.97473295127806e-12
+   -1.098184046596749e-11
+    8.375227268660543e-11
+   -5.818752536077342e-13
+   -1.972410555894047e-12
+   -2.196902859567094e-11
+    8.014261404810914e-11
+ 6.17e+10    
+    8.025581124848554e-11
+   -2.197172637811368e-11
+    8.372850448440656e-11
+   -1.974270104260037e-12
+   -1.098672807981009e-11
+    8.375033048481465e-11
+   -5.778235312142425e-13
+   -1.971965397451196e-12
+   -2.197381182836115e-11
+    8.013335080533276e-11
+ 6.18e+10    
+    8.024645569307188e-11
+   -2.197649749397812e-11
+    8.372654556966101e-11
+   -1.973789190870541e-12
+   -1.099162493999596e-11
+    8.374837244284017e-11
+   -5.737623009199553e-13
+   -1.971502221319092e-12
+   -2.197859169181233e-11
+    8.012406075374179e-11
+ 6.19e+10    
+    8.023707312584066e-11
+   -2.198126505256813e-11
+     8.37245706914066e-11
+   -1.973290202780438e-12
+    -1.09965310462424e-11
+    8.374639851231436e-11
+   -5.696916823751394e-13
+   -1.971021018821822e-12
+   -2.198336809345108e-11
+    8.011474387858092e-11
+ 6.2e+10     
+    8.022766353216319e-11
+   -2.198602896089206e-11
+    8.372257980104029e-11
+    -1.97277313200669e-12
+   -1.100144639820107e-11
+    8.374440864491446e-11
+   -5.656117956136714e-13
+   -1.970521781627434e-12
+   -2.198814094055816e-11
+    8.010540016520753e-11
+ 6.21e+10    
+    8.021822689752434e-11
+   -2.199078912581498e-11
+    8.372057285000539e-11
+    -1.97223797091241e-12
+   -1.100637099545689e-11
+    8.374240279236249e-11
+     -5.6152276104745e-13
+    -1.97000450174802e-12
+   -2.199291014027011e-11
+    8.009602959909034e-11
+ 6.22e+10    
+    8.020876320752161e-11
+   -2.199554545406046e-11
+    8.371854978979176e-11
+   -1.971684712206908e-12
+   -1.101130483752706e-11
+    8.374038090642526e-11
+   -5.574246994607274e-13
+   -1.969469171539766e-12
+    -2.19976755995808e-11
+    8.008663216580843e-11
+ 6.23e+10    
+     8.01992724478636e-11
+    -2.20002978522122e-11
+    8.371651057193595e-11
+   -1.971113348945681e-12
+   -1.101624792386023e-11
+    8.373834293891437e-11
+   -5.533177320043856e-13
+   -1.968915783702989e-12
+   -2.200243722534312e-11
+    8.007720785105016e-11
+ 6.24e+10    
+    8.018975460436912e-11
+   -2.200504622671549e-11
+    8.371445514802041e-11
+   -1.970523874530489e-12
+   -1.102120025383526e-11
+    8.373628884168599e-11
+   -5.492019801901723e-13
+   -1.968344331282182e-12
+   -2.200719492427062e-11
+    8.006775664061182e-11
+ 6.25e+10    
+    8.018020966296602e-11
+   -2.200979048387912e-11
+    8.371238346967435e-11
+   -1.969916282709343e-12
+   -1.102616182676053e-11
+    8.373421856664114e-11
+   -5.450775658848566e-13
+   -1.967754807666026e-12
+   -2.201194860293916e-11
+    8.005827852039669e-11
+ 6.26e+10    
+     8.01706376096901e-11
+   -2.201453052987695e-11
+    8.371029548857318e-11
+   -1.969290567576504e-12
+   -1.103113264187276e-11
+    8.373213206572549e-11
+   -5.409446113043449e-13
+   -1.967147206587419e-12
+   -2.201669816778865e-11
+    8.004877347641393e-11
+ 6.27e+10    
+    8.016103843068405e-11
+   -2.201926627074961e-11
+    8.370819115643886e-11
+   -1.968646723572504e-12
+   -1.103611269833625e-11
+    8.373002929092952e-11
+    -5.36803239007733e-13
+   -1.966521522123484e-12
+   -2.202144352512469e-11
+    8.003924149477763e-11
+ 6.28e+10    
+    8.015141211219589e-11
+   -2.202399761240617e-11
+    8.370607042503954e-11
+   -1.967984745484096e-12
+   -1.104110199524184e-11
+     8.37279101942883e-11
+   -5.326535718913062e-13
+   -1.965877748695558e-12
+    -2.20261845811202e-11
+    8.002968256170518e-11
+ 6.29e+10    
+    8.014175864057854e-11
+   -2.202872446062593e-11
+    8.370393324618991e-11
+   -1.967304628444244e-12
+   -1.104610053160596e-11
+    8.372577472788168e-11
+   -5.284957331824889e-13
+   -1.965215881069193e-12
+   -2.203092124181731e-11
+    8.002009666351682e-11
+ 6.3e+10     
+    8.013207800228849e-11
+   -2.203344672106012e-11
+    8.370177957175095e-11
+   -1.966606367932117e-12
+   -1.105110830636973e-11
+    8.372362284383401e-11
+   -5.243298464337341e-13
+   -1.964535914354141e-12
+   -2.203565341312887e-11
+    8.001048378663419e-11
+ 6.31e+10    
+    8.012237018388429e-11
+   -2.203816429923356e-11
+    8.369960935363028e-11
+   -1.965889959772994e-12
+   -1.105612531839819e-11
+    8.372145449431481e-11
+    -5.20156035516367e-13
+   -1.963837844004316e-12
+   -2.204038100084034e-11
+    8.000084391757937e-11
+ 6.32e+10    
+    8.011263517202605e-11
+   -2.204287710054653e-11
+    8.369742254378173e-11
+   -1.965155400138286e-12
+   -1.106115156647914e-11
+    8.371926963153815e-11
+   -5.159744246143656e-13
+   -1.963121665817754e-12
+   -2.204510391061151e-11
+    7.999117704297386e-11
+ 6.33e+10    
+    8.010287295347405e-11
+   -2.204758503027645e-11
+    8.369521909420572e-11
+   -1.964402685545393e-12
+   -1.106618704932243e-11
+    8.371706820776269e-11
+   -5.117851382181118e-13
+   -1.962387375936585e-12
+   -2.204982204797814e-11
+    7.998148314953732e-11
+ 6.34e+10    
+    8.009308351508789e-11
+   -2.205228799357968e-11
+    8.369299895694918e-11
+    -1.96363181285772e-12
+   -1.107123176555903e-11
+    8.371485017529243e-11
+   -5.075883011180622e-13
+   -1.961634970846988e-12
+   -2.205453531835393e-11
+    7.997176222408698e-11
+ 6.35e+10    
+    8.008326684382512e-11
+   -2.205698589549322e-11
+    8.369076208410549e-11
+   -1.962842779284531e-12
+   -1.107628571374011e-11
+     8.37126154864757e-11
+   -5.033840383984046e-13
+   -1.960864447379083e-12
+   -2.205924362703207e-11
+    7.996201425353605e-11
+ 6.36e+10    
+     8.00734229267407e-11
+   -2.206167864093672e-11
+    8.368850842781496e-11
+   -1.962035582380918e-12
+   -1.108134889233626e-11
+    8.371036409370609e-11
+   -4.991724754306226e-13
+   -1.960075802706928e-12
+   -2.206394687918726e-11
+    7.995223922489302e-11
+ 6.37e+10    
+    8.006355175098536e-11
+   -2.206636613471401e-11
+    8.368623794026399e-11
+   -1.961210220047671e-12
+   -1.108642129973652e-11
+    8.370809594942213e-11
+   -4.949537378670623e-13
+   -1.959269034348377e-12
+   -2.206864497987727e-11
+    7.994243712526049e-11
+ 6.38e+10    
+    8.005365330380481e-11
+   -2.207104828151504e-11
+    8.368395057368617e-11
+   -1.960366690531187e-12
+   -1.109150293424758e-11
+     8.37058110061072e-11
+   -4.907279516344117e-13
+   -1.958444140165046e-12
+   -2.207333783404497e-11
+    7.993260794183455e-11
+ 6.39e+10    
+    8.004372757253912e-11
+   -2.207572498591781e-11
+    8.368164628036159e-11
+   -1.959504992423377e-12
+   -1.109659379409301e-11
+    8.370350921628995e-11
+   -4.864952429271502e-13
+   -1.957601118362179e-12
+      -2.207802534652e-11
+    7.992275166190313e-11
+ 6.4e+10     
+    8.003377454462116e-11
+   -2.208039615238997e-11
+    8.367932501261732e-11
+   -1.958625124661513e-12
+    -1.11016938774123e-11
+    8.370119053254411e-11
+   -4.822557382009535e-13
+   -1.956739967488567e-12
+   -2.208270742202065e-11
+    7.991286827284545e-11
+ 6.41e+10    
+     8.00237942075758e-11
+   -2.208506168529089e-11
+    8.367698672282704e-11
+   -1.957727086528135e-12
+   -1.110680318226008e-11
+     8.36988549074886e-11
+    -4.78009564166052e-13
+   -1.955860686436432e-12
+   -2.208738396515577e-11
+    7.990295776213117e-11
+ 6.42e+10    
+    8.001378654901898e-11
+   -2.208972148887335e-11
+    8.367463136341194e-11
+   -1.956810877650877e-12
+    -1.11119217066054e-11
+    8.369650229378762e-11
+   -4.737568477805376e-13
+   -1.954963274441304e-12
+   -2.209205488042643e-11
+    7.989302011731871e-11
+ 6.43e+10    
+    8.000375155665664e-11
+   -2.209437546728553e-11
+    8.367225888683969e-11
+    -1.95587649800238e-12
+   -1.111704944833076e-11
+    8.369413264415088e-11
+   -4.694977162436455e-13
+   -1.954047731081893e-12
+   -2.209672007222803e-11
+    7.988305532605514e-11
+ 6.44e+10    
+    7.999368921828383e-11
+   -2.209902352457278e-11
+    8.366986924562549e-11
+   -1.954923947900052e-12
+   -1.112218640523139e-11
+    8.369174591133333e-11
+   -4.652322969889828e-13
+   -1.953114056279951e-12
+   -2.210137944485197e-11
+    7.987306337607488e-11
+ 6.45e+10    
+     7.99835995217837e-11
+   -2.210366556467949e-11
+    8.366746239233125e-11
+   -1.953953228006027e-12
+   -1.112733257501449e-11
+    8.368934204813558e-11
+   -4.609607176777055e-13
+   -1.952162250300145e-12
+   -2.210603290248762e-11
+    7.986304425519853e-11
+ 6.46e+10    
+    7.997348245512641e-11
+   -2.210830149145121e-11
+    8.366503827956693e-11
+   -1.952964339326865e-12
+    -1.11324879552985e-11
+      8.3686921007404e-11
+   -4.566831061916732e-13
+    -1.95119231374987e-12
+   -2.211068034922427e-11
+    7.985299795133212e-11
+ 6.47e+10    
+    7.996333800636848e-11
+   -2.211293120863626e-11
+    8.366259685998942e-11
+   -1.951957283213461e-12
+    -1.11376525436121e-11
+    8.368448274203053e-11
+    -4.52399590626565e-13
+   -1.950204247579126e-12
+   -2.211532168905281e-11
+    7.984292445246622e-11
+ 6.48e+10    
+    7.995316616365174e-11
+   -2.211755461988772e-11
+    8.366013808630314e-11
+   -1.950932061360847e-12
+   -1.114282633739372e-11
+    8.368202720495308e-11
+   -4.481102992849388e-13
+   -1.949198053080317e-12
+   -2.211995682586798e-11
+     7.98328237466752e-11
+ 6.49e+10    
+    7.994296691520215e-11
+   -2.212217162876557e-11
+    8.365766191126034e-11
+   -1.949888675807964e-12
+   -1.114800933399061e-11
+    8.367955434915529e-11
+   -4.438153606692683e-13
+   -1.948173731888111e-12
+   -2.212458566346987e-11
+    7.982269582211571e-11
+ 6.5e+10     
+    7.993274024932916e-11
+   -2.212678213873828e-11
+    8.365516828766087e-11
+   -1.948827128937487e-12
+   -1.115320153065817e-11
+    8.367706412766731e-11
+   -4.395149034749437e-13
+   -1.947131285979204e-12
+   -2.212920810556629e-11
+    7.981254066702654e-11
+ 6.51e+10    
+    7.992248615442497e-11
+   -2.213138605318506e-11
+    8.365265716835261e-11
+   -1.947747423475623e-12
+   -1.115840292455922e-11
+    8.367455649356515e-11
+   -4.352090565832192e-13
+   -1.946070717672177e-12
+   -2.213382405577435e-11
+    7.980235826972726e-11
+ 6.52e+10    
+    7.991220461896291e-11
+   -2.213598327539754e-11
+    8.365012850623123e-11
+   -1.946649562491857e-12
+   -1.116361351276323e-11
+    8.367203139997125e-11
+   -4.308979490541562e-13
+   -1.944992029627274e-12
+   -2.213843341762264e-11
+    7.979214861861748e-11
+ 6.53e+10    
+    7.990189563149756e-11
+   -2.214057370858198e-11
+    8.364758225424081e-11
+   -1.945533549398746e-12
+   -1.116883329224563e-11
+    8.366948880005442e-11
+   -4.265817101195041e-13
+   -1.943895224846187e-12
+   -2.214303609455299e-11
+     7.97819117021759e-11
+ 6.54e+10    
+    7.989155918066308e-11
+   -2.214515725586105e-11
+    8.364501836537348e-11
+   -1.944399387951702e-12
+   -1.117406225988712e-11
+    8.366692864703022e-11
+   -4.222604691755574e-13
+    -1.94278030667185e-12
+   -2.214763198992263e-11
+    7.977164750895966e-11
+ 6.55e+10    
+    7.988119525517281e-11
+   -2.214973382027587e-11
+    8.364243679266976e-11
+   -1.943247082248724e-12
+   -1.117930041247292e-11
+    8.366435089416079e-11
+   -4.179343557759969e-13
+   -1.941647278788199e-12
+   -2.215222100700601e-11
+    7.976135602760313e-11
+ 6.56e+10    
+    7.987080384381802e-11
+   -2.215430330478804e-11
+    8.363983748921877e-11
+   -1.942076636730143e-12
+   -1.118454774669213e-11
+    8.366175549475536e-11
+   -4.136034996246711e-13
+   -1.940496145219963e-12
+   -2.215680304899689e-11
+    7.975103724681758e-11
+ 6.57e+10    
+    7.986038493546747e-11
+   -2.215886561228157e-11
+    8.363722040815858e-11
+   -1.940888056178375e-12
+   -1.118980425913707e-11
+    8.365914240216999e-11
+   -4.092680305683695e-13
+   -1.939326910332404e-12
+   -2.216137801901025e-11
+    7.974069115538989e-11
+ 6.58e+10    
+    7.984993851906613e-11
+   -2.216342064556482e-11
+    8.363458550267576e-11
+   -1.939681345717666e-12
+   -1.119506994630251e-11
+    8.365651156980799e-11
+   -4.049280785895559e-13
+   -1.938139578831086e-12
+   -2.216594582008428e-11
+    7.973031774218196e-11
+ 6.59e+10    
+    7.983946458363492e-11
+   -2.216796830737275e-11
+    8.363193272600611e-11
+   -1.938456510813787e-12
+    -1.12003448045851e-11
+    8.365386295112004e-11
+   -4.005837737990892e-13
+   -1.936934155761596e-12
+    -2.21705063551825e-11
+    7.971991699612993e-11
+ 6.6e+10     
+    7.982896311826946e-11
+   -2.217250850036862e-11
+    8.362926203143449e-11
+   -1.937213557273775e-12
+    -1.12056288302827e-11
+    8.365119649960441e-11
+   -3.962352464288966e-13
+   -1.935710646509284e-12
+   -2.217505952719564e-11
+    7.970948890624328e-11
+ 6.61e+10    
+    7.981843411213938e-11
+    -2.21770411271463e-11
+    8.362657337229521e-11
+   -1.935952491245624e-12
+   -1.121092201959372e-11
+    8.364851216880697e-11
+   -3.918826268246287e-13
+   -1.934469056799015e-12
+   -2.217960523894376e-11
+    7.969903346160408e-11
+ 6.62e+10    
+    7.980787755448752e-11
+   -2.218156609023205e-11
+    8.362386670197223e-11
+   -1.934673319217994e-12
+   -1.121622436861649e-11
+    8.364580991232133e-11
+   -3.875260454382944e-13
+   -1.933209392694872e-12
+   -2.218414339317819e-11
+    7.968855065136637e-11
+ 6.63e+10    
+    7.979729343462924e-11
+   -2.218608329208673e-11
+    8.362114197389891e-11
+   -1.933376048019937e-12
+   -1.122153587334865e-11
+    8.364308968378957e-11
+   -3.831656328208656e-13
+   -1.931931660599843e-12
+   -2.218867389258364e-11
+    7.967804046475499e-11
+ 6.64e+10    
+    7.978668174195166e-11
+   -2.219059263510791e-11
+    8.361839914155903e-11
+   -1.932060684820485e-12
+   -1.122685652968653e-11
+    8.364035143690153e-11
+   -3.788015196148744e-13
+   -1.930635867255583e-12
+   -2.219319663978023e-11
+    7.966750289106552e-11
+ 6.65e+10    
+    7.977604246591267e-11
+   -2.219509402163163e-11
+    8.361563815848593e-11
+   -1.930727237128445e-12
+   -1.123218633342453e-11
+    8.363759512539578e-11
+   -3.744338365469533e-13
+   -1.929322019742046e-12
+   -2.219771153732551e-11
+    7.965693791966264e-11
+ 6.66e+10    
+    7.976537559604063e-11
+   -2.219958735393478e-11
+    8.361285897826354e-11
+   -1.929375712791987e-12
+   -1.123752528025453e-11
+    8.363482070305948e-11
+   -3.700627144204014e-13
+    -1.92799012547722e-12
+   -2.220221848771658e-11
+    7.964634553998036e-11
+ 6.67e+10    
+    7.975468112193297e-11
+     -2.2204072534237e-11
+    8.361006155452615e-11
+   -1.928006119998343e-12
+   -1.124287336576529e-11
+     8.36320281237284e-11
+   -3.656882841076815e-13
+   -1.926640192216801e-12
+   -2.220671739339204e-11
+    7.963572574152058e-11
+ 6.68e+10    
+    7.974395903325625e-11
+    -2.22085494647028e-11
+    8.360724584095899e-11
+   -1.926618467273428e-12
+   -1.124823058544194e-11
+    8.362921734128766e-11
+    -3.61310676542942e-13
+   -1.925272228053842e-12
+   -2.221120815673423e-11
+    7.962507851385265e-11
+ 6.69e+10    
+    7.973320931974478e-11
+   -2.221301804744361e-11
+    8.360441179129798e-11
+   -1.925212763481527e-12
+    -1.12535969346653e-11
+    8.362638830967121e-11
+   -3.569300227144956e-13
+   -1.923886241418433e-12
+    -2.22156906800711e-11
+    7.961440384661283e-11
+ 6.7e+10     
+    7.972243197120021e-11
+   -2.221747818451992e-11
+    8.360155935933017e-11
+   -1.923789017824887e-12
+   -1.125897240871145e-11
+    8.362354098286309e-11
+   -3.525464536572794e-13
+   -1.922482241077362e-12
+   -2.222016486567861e-11
+    7.960370172950336e-11
+ 6.71e+10    
+    7.971162697749118e-11
+   -2.222192977794345e-11
+    8.359868849889419e-11
+   -1.922347239843382e-12
+   -1.126435700275108e-11
+     8.36206753148966e-11
+    -3.48160100445321e-13
+   -1.921060236133757e-12
+   -2.222463061578249e-11
+    7.959297215229189e-11
+ 6.72e+10    
+    7.970079432855173e-11
+   -2.222637272967894e-11
+    8.359579916387998e-11
+   -1.920887439414108e-12
+   -1.126975071184896e-11
+    8.361779125985472e-11
+   -3.437710941841622e-13
+    -1.91962023602673e-12
+    -2.22290878325604e-11
+    7.958221510481074e-11
+ 6.73e+10    
+    7.968993401438166e-11
+   -2.223080694164674e-11
+    8.359289130822959e-11
+   -1.919409626751007e-12
+   -1.127515353096349e-11
+    8.361488877187112e-11
+   -3.393795660032903e-13
+   -1.918162250531007e-12
+   -2.223353641814442e-11
+    7.957143057695673e-11
+ 6.74e+10    
+    7.967904602504529e-11
+   -2.223523231572446e-11
+    8.358996488593674e-11
+   -1.917913812404495e-12
+   -1.128056545494604e-11
+    8.361196780512961e-11
+   -3.349856470485464e-13
+   -1.916686289756566e-12
+   -2.223797627462255e-11
+    7.956061855868964e-11
+ 6.75e+10    
+    7.966813035067072e-11
+    -2.22396487537494e-11
+    8.358701985104774e-11
+   -1.916400007260994e-12
+   -1.128598647854061e-11
+    8.360902831386438e-11
+    -3.30589468474525e-13
+   -1.915192364148233e-12
+   -2.224240730404125e-11
+    7.954977904003236e-11
+ 6.76e+10    
+    7.965718698144981e-11
+   -2.224405615752059e-11
+    8.358405615766135e-11
+   -1.914868222542597e-12
+   -1.129141659638319e-11
+    8.360607025236099e-11
+   -3.261911614369647e-13
+   -1.913680484485304e-12
+   -2.224682940840761e-11
+    7.953891201107006e-11
+ 6.77e+10    
+    7.964621590763687e-11
+   -2.224845442880084e-11
+    8.358107375992915e-11
+   -1.913318469806592e-12
+   -1.129685580300132e-11
+    8.360309357495561e-11
+   -3.217908570851178e-13
+   -1.912150661881156e-12
+   -2.225124248969103e-11
+    7.952801746194949e-11
+ 6.78e+10    
+    7.963521711954862e-11
+   -2.225284346931904e-11
+    8.357807261205569e-11
+   -1.911750760945071e-12
+   -1.130230409281363e-11
+    8.360009823603625e-11
+   -3.173886865541285e-13
+   -1.910602907782828e-12
+   -2.225564644982593e-11
+    7.951709538287859e-11
+ 6.79e+10    
+    7.962419060756287e-11
+   -2.225722318077209e-11
+    8.357505266829887e-11
+   -1.910165108184459e-12
+   -1.130776146012929e-11
+    8.359708419004196e-11
+   -3.129847809573992e-13
+   -1.909037233970597e-12
+   -2.226004119071339e-11
+    7.950614576412547e-11
+ 6.8e+10     
+     7.96131363621192e-11
+   -2.226159346482739e-11
+    8.357201388297028e-11
+    -1.90856152408513e-12
+   -1.131322789914765e-11
+    8.359405139146436e-11
+   -3.085792713789282e-13
+   -1.907453652557592e-12
+   -2.226442661422377e-11
+    7.949516859601863e-11
+ 6.81e+10    
+    7.960205437371676e-11
+   -2.226595422312449e-11
+    8.356895621043499e-11
+   -1.906940021540879e-12
+   -1.131870340395768e-11
+    8.359099979484688e-11
+   -3.041722888656871e-13
+   -1.905852175989314e-12
+   -2.226880262219842e-11
+    7.948416386894565e-11
+ 6.82e+10    
+    7.959094463291512e-11
+   -2.227030535727787e-11
+     8.35658796051126e-11
+   -1.905300613778518e-12
+   -1.132418796853761e-11
+    8.358792935478542e-11
+   -2.997639644199428e-13
+   -1.904232817043244e-12
+   -2.227316911645214e-11
+    7.947313157335306e-11
+ 6.83e+10    
+     7.95798071303328e-11
+   -2.227464676887854e-11
+    8.356278402147689e-11
+   -1.903643314357389e-12
+   -1.132968158675447e-11
+    8.358484002592852e-11
+   -2.953544289916138e-13
+   -1.902595588828374e-12
+   -2.227752599877519e-11
+    7.946207169974557e-11
+ 6.84e+10    
+    7.956864185664753e-11
+   -2.227897835949658e-11
+     8.35596694140564e-11
+   -1.901968137168903e-12
+    -1.13351842523636e-11
+    8.358173176297796e-11
+   -2.909438134706093e-13
+   -1.900940504784753e-12
+   -2.228187317093548e-11
+    7.945098423868585e-11
+ 6.85e+10    
+    7.955744880259482e-11
+   -2.228330003068312e-11
+    8.355653573743449e-11
+   -1.900275096436028e-12
+   -1.134069595900833e-11
+    8.357860452068867e-11
+   -2.865322486791638e-13
+    -1.89926757868303e-12
+   -2.228621053468088e-11
+    7.943986918079394e-11
+ 6.86e+10    
+    7.954622795896832e-11
+   -2.228761168397274e-11
+    8.355338294625009e-11
+   -1.898564206712819e-12
+   -1.134621670021954e-11
+    8.357545825386926e-11
+   -2.821198653641831e-13
+   -1.897576824623988e-12
+   -2.229053799174122e-11
+    7.942872651674655e-11
+ 6.87e+10    
+    7.953497931661881e-11
+   -2.229191322088533e-11
+    8.355021099519745e-11
+   -1.896835482883923e-12
+   -1.135174646941519e-11
+    8.357229291738202e-11
+   -2.777067941895728e-13
+   -1.895868257038065e-12
+   -2.229485544383053e-11
+    7.941755623727689e-11
+ 6.88e+10    
+    7.952370286645359e-11
+   -2.229620454292849e-11
+    8.354701983902668e-11
+   -1.895088940164051e-12
+   -1.135728525990007e-11
+    8.356910846614377e-11
+   -2.732931657285995e-13
+   -1.894141890684836e-12
+    -2.22991627926493e-11
+    7.940635833317382e-11
+ 6.89e+10    
+    7.951239859943664e-11
+   -2.230048555159986e-11
+    8.354380943254433e-11
+   -1.893324594097477e-12
+    -1.13628330648653e-11
+    8.356590485512567e-11
+   -2.688791104562164e-13
+   -1.892397740652587e-12
+    -2.23034599398866e-11
+    7.939513279528197e-11
+ 6.9e+10     
+    7.950106650658758e-11
+   -2.230475614838893e-11
+    8.354057973061292e-11
+   -1.891542460557517e-12
+   -1.136838987738798e-11
+    8.356268203935351e-11
+   -2.644647587414245e-13
+   -1.890635822357737e-12
+   -2.230774678722221e-11
+    7.938387961450061e-11
+ 6.91e+10    
+    7.948970657898158e-11
+   -2.230901623477965e-11
+    8.353733068815235e-11
+   -1.889742555745976e-12
+   -1.137395569043092e-11
+    8.355943997390855e-11
+   -2.600502408396257e-13
+   -1.888856151544395e-12
+   -2.231202323632902e-11
+    7.937259878178403e-11
+ 6.92e+10    
+    7.947831880774868e-11
+   -2.231326571225243e-11
+    8.353406226013948e-11
+   -1.887924896192623e-12
+   -1.137953049684219e-11
+    8.355617861392731e-11
+   -2.556356868849744e-13
+   -1.887058744283786e-12
+   -2.231628918887501e-11
+    7.936129028814014e-11
+ 6.93e+10    
+    7.946690318407332e-11
+   -2.231750448228623e-11
+    8.353077440160842e-11
+   -1.886089498754649e-12
+    -1.13851142893548e-11
+    8.355289791460211e-11
+   -2.512212268827533e-13
+   -1.885243616973754e-12
+   -2.232054454652561e-11
+    7.934995412463098e-11
+ 6.94e+10    
+    7.945545969919448e-11
+    -2.23217324463611e-11
+    8.352746706765113e-11
+   -1.884236380616093e-12
+   -1.139070706058642e-11
+    8.354959783118152e-11
+   -2.468069907017472e-13
+   -1.883410786338231e-12
+   -2.232478921094588e-11
+    7.933859028237199e-11
+ 6.95e+10    
+    7.944398834440446e-11
+    -2.23259495059601e-11
+    8.352414021341809e-11
+   -1.882365559287285e-12
+   -1.139630880303902e-11
+    8.354627831897039e-11
+   -2.423931080666279e-13
+    -1.88156026942667e-12
+   -2.232902308380263e-11
+     7.93271987525314e-11
+ 6.96e+10    
+    7.943248911104926e-11
+   -2.233015556257174e-11
+    8.352079379411774e-11
+   -1.880477052604277e-12
+   -1.140191950909852e-11
+     8.35429393333305e-11
+   -2.379797085503487e-13
+   -1.879692083613521e-12
+   -2.233324606676686e-11
+     7.93157795263303e-11
+ 6.97e+10    
+     7.94209619905277e-11
+   -2.233435051769204e-11
+    8.351742776501762e-11
+   -1.878570878728261e-12
+   -1.140753917103459e-11
+     8.35395808296808e-11
+   -2.335669215665471e-13
+    -1.87780624659764e-12
+   -2.233745806151571e-11
+    7.930433259504187e-11
+ 6.98e+10    
+    7.940940697429119e-11
+   -2.233853427282677e-11
+    8.351404208144424e-11
+   -1.876647056144954e-12
+   -1.141316778100018e-11
+    8.353620276349734e-11
+   -2.291548763619728e-13
+   -1.875902776401769e-12
+   -2.234165896973475e-11
+    7.929285794999126e-11
+ 6.99e+10    
+     7.93978240538438e-11
+   -2.234270672949397e-11
+    8.351063669878398e-11
+   -1.874705603664034e-12
+   -1.141880533103153e-11
+    8.353280509031467e-11
+   -2.247437020089124e-13
+   -1.873981691371899e-12
+   -2.234584869312049e-11
+    7.928135558255544e-11
+ 7e+10       
+    7.938621322074103e-11
+   -2.234686778922564e-11
+    8.350721157248263e-11
+   -1.872746540418529e-12
+   -1.142445181304755e-11
+    8.352938776572516e-11
+   -2.203335273976321e-13
+   -1.872043010176729e-12
+   -2.235002713338225e-11
+     7.92698254841625e-11
* NOTE: Solution at 1e+08 Hz used as DC point.

.ends
