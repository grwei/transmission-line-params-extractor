* begin ansoft header
* node 1 Diff1
* node 2 Comm1
* node 3 Diff2
* node 4 Comm2
* node 5 Diff3
* node 6 Comm3
* node 7 Diff4
* node 8 Comm4
* node 9 Diff5
* node 10 Comm5
* node 11 Diff6
* node 12 Comm6
* node 13 Diff7
* node 14 Comm7
* node 15 Diff8
* node 16 Comm8
* node 17 Diff9
* node 18 Comm9
* node 19 Diff10
* node 20 Comm10
* node 21 Diff11
* node 22 Comm11
* node 23 Diff12
* node 24 Comm12
* node 25 Diff13
* node 26 Comm13
* node 27 Diff14
* node 28 Comm14
* node 29 Diff15
* node 30 Comm15
* node 31 Diff16
* node 32 Comm16
* 
* created by ElectronicsDesktop
* end ansoft header

.subckt m16lines_port_lfws 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 
v2_3 2 33 dc 0.0
v2_4 2 34 dc 0.0
v2_7 2 35 dc 0.0
v2_8 2 36 dc 0.0
v2_9 2 37 dc 0.0
v2_10 2 38 dc 0.0
v2_11 2 39 dc 0.0
v2_14 2 40 dc 0.0
v2_15 2 41 dc 0.0
v2_16 2 42 dc 0.0
v3_4 3 43 dc 0.0
v3_5 3 44 dc 0.0
v3_6 3 45 dc 0.0
v3_7 3 46 dc 0.0
v3_8 3 47 dc 0.0
v3_9 3 48 dc 0.0
v3_10 3 49 dc 0.0
v3_11 3 50 dc 0.0
v3_12 3 51 dc 0.0
v3_13 3 52 dc 0.0
v3_15 3 53 dc 0.0
v3_16 3 54 dc 0.0
v4_5 4 55 dc 0.0
v4_6 4 56 dc 0.0
v4_7 4 57 dc 0.0
v4_8 4 58 dc 0.0
v4_9 4 59 dc 0.0
v4_10 4 60 dc 0.0
v4_11 4 61 dc 0.0
v4_12 4 62 dc 0.0
v4_13 4 63 dc 0.0
v4_14 4 64 dc 0.0
v5_6 5 65 dc 0.0
v5_7 5 66 dc 0.0
v5_8 5 67 dc 0.0
v5_9 5 68 dc 0.0
v5_10 5 69 dc 0.0
v5_11 5 70 dc 0.0
v5_12 5 71 dc 0.0
v5_13 5 72 dc 0.0
v5_14 5 73 dc 0.0
v5_15 5 74 dc 0.0
v6_7 6 75 dc 0.0
v6_8 6 76 dc 0.0
v6_9 6 77 dc 0.0
v6_10 6 78 dc 0.0
v6_11 6 79 dc 0.0
v6_12 6 80 dc 0.0
v6_13 6 81 dc 0.0
v6_14 6 82 dc 0.0
v6_15 6 83 dc 0.0
v6_16 6 84 dc 0.0
v7_8 7 85 dc 0.0
v7_9 7 86 dc 0.0
v7_10 7 87 dc 0.0
v7_11 7 88 dc 0.0
v7_12 7 89 dc 0.0
v7_13 7 90 dc 0.0
v7_14 7 91 dc 0.0
v7_15 7 92 dc 0.0
v7_16 7 93 dc 0.0
v8_9 8 94 dc 0.0
v8_10 8 95 dc 0.0
v8_11 8 96 dc 0.0
v8_12 8 97 dc 0.0
v8_13 8 98 dc 0.0
v8_14 8 99 dc 0.0
v8_15 8 100 dc 0.0
v8_16 8 101 dc 0.0
v9_10 9 102 dc 0.0
v9_11 9 103 dc 0.0
v9_12 9 104 dc 0.0
v9_13 9 105 dc 0.0
v9_14 9 106 dc 0.0
v9_15 9 107 dc 0.0
v9_16 9 108 dc 0.0
v10_11 10 109 dc 0.0
v10_12 10 110 dc 0.0
v10_13 10 111 dc 0.0
v10_14 10 112 dc 0.0
v10_15 10 113 dc 0.0
v10_16 10 114 dc 0.0
v11_12 11 115 dc 0.0
v11_13 11 116 dc 0.0
v11_14 11 117 dc 0.0
v11_15 11 118 dc 0.0
v11_16 11 119 dc 0.0
v12_13 12 120 dc 0.0
v12_14 12 121 dc 0.0
v12_15 12 122 dc 0.0
v12_16 12 123 dc 0.0
v13_14 13 124 dc 0.0
v13_15 13 125 dc 0.0
v13_16 13 126 dc 0.0
v14_15 14 127 dc 0.0
v14_16 14 128 dc 0.0
v15_16 15 129 dc 0.0
v18_19 18 130 dc 0.0
v18_20 18 131 dc 0.0
v18_21 18 132 dc 0.0
v18_23 18 133 dc 0.0
v18_24 18 134 dc 0.0
v18_25 18 135 dc 0.0
v18_26 18 136 dc 0.0
v18_27 18 137 dc 0.0
v18_30 18 138 dc 0.0
v18_31 18 139 dc 0.0
v18_32 18 140 dc 0.0
v19_20 19 141 dc 0.0
v19_21 19 142 dc 0.0
v19_22 19 143 dc 0.0
v19_23 19 144 dc 0.0
v19_24 19 145 dc 0.0
v19_25 19 146 dc 0.0
v19_26 19 147 dc 0.0
v19_27 19 148 dc 0.0
v19_28 19 149 dc 0.0
v19_29 19 150 dc 0.0
v19_30 19 151 dc 0.0
v19_32 19 152 dc 0.0
v20_21 20 153 dc 0.0
v20_22 20 154 dc 0.0
v20_23 20 155 dc 0.0
v20_24 20 156 dc 0.0
v20_25 20 157 dc 0.0
v20_26 20 158 dc 0.0
v20_27 20 159 dc 0.0
v20_28 20 160 dc 0.0
v20_29 20 161 dc 0.0
v20_30 20 162 dc 0.0
v20_31 20 163 dc 0.0
v21_22 21 164 dc 0.0
v21_23 21 165 dc 0.0
v21_24 21 166 dc 0.0
v21_25 21 167 dc 0.0
v21_26 21 168 dc 0.0
v21_27 21 169 dc 0.0
v21_28 21 170 dc 0.0
v21_29 21 171 dc 0.0
v21_30 21 172 dc 0.0
v21_31 21 173 dc 0.0
v22_23 22 174 dc 0.0
v22_24 22 175 dc 0.0
v22_25 22 176 dc 0.0
v22_26 22 177 dc 0.0
v22_27 22 178 dc 0.0
v22_28 22 179 dc 0.0
v22_29 22 180 dc 0.0
v22_30 22 181 dc 0.0
v22_31 22 182 dc 0.0
v23_17 23 183 dc 0.0
v23_24 23 184 dc 0.0
v23_25 23 185 dc 0.0
v23_26 23 186 dc 0.0
v23_27 23 187 dc 0.0
v23_28 23 188 dc 0.0
v23_29 23 189 dc 0.0
v23_30 23 190 dc 0.0
v23_31 23 191 dc 0.0
v23_32 23 192 dc 0.0
v24_25 24 193 dc 0.0
v24_26 24 194 dc 0.0
v24_27 24 195 dc 0.0
v24_28 24 196 dc 0.0
v24_29 24 197 dc 0.0
v24_30 24 198 dc 0.0
v24_31 24 199 dc 0.0
v24_32 24 200 dc 0.0
v25_26 25 201 dc 0.0
v25_27 25 202 dc 0.0
v25_28 25 203 dc 0.0
v25_29 25 204 dc 0.0
v25_30 25 205 dc 0.0
v25_31 25 206 dc 0.0
v25_32 25 207 dc 0.0
v26_27 26 208 dc 0.0
v26_28 26 209 dc 0.0
v26_29 26 210 dc 0.0
v26_30 26 211 dc 0.0
v26_31 26 212 dc 0.0
v26_32 26 213 dc 0.0
v27_28 27 214 dc 0.0
v27_29 27 215 dc 0.0
v27_30 27 216 dc 0.0
v27_31 27 217 dc 0.0
v27_32 27 218 dc 0.0
v28_29 28 219 dc 0.0
v28_30 28 220 dc 0.0
v28_31 28 221 dc 0.0
v28_32 28 222 dc 0.0
v29_30 29 223 dc 0.0
v29_31 29 224 dc 0.0
v29_32 29 225 dc 0.0
v30_31 30 226 dc 0.0
v30_32 30 227 dc 0.0
v31_32 31 228 dc 0.0
v1_0 1 229 dc 0.0
v2_0 2 230 dc 0.0
v3_0 3 231 dc 0.0
v4_0 4 232 dc 0.0
v5_0 5 233 dc 0.0
v6_0 6 234 dc 0.0
v7_0 7 235 dc 0.0
v8_0 8 236 dc 0.0
v9_0 9 237 dc 0.0
v10_0 10 238 dc 0.0
v11_0 11 239 dc 0.0
v12_0 12 240 dc 0.0
v13_0 13 241 dc 0.0
v14_0 14 242 dc 0.0
v15_0 15 243 dc 0.0
v16_0 16 244 dc 0.0
v17_0 17 245 dc 0.0
v18_0 18 246 dc 0.0
v19_0 19 247 dc 0.0
v20_0 20 248 dc 0.0
v21_0 21 249 dc 0.0
v22_0 22 250 dc 0.0
v23_0 23 251 dc 0.0
v24_0 24 252 dc 0.0
v25_0 25 253 dc 0.0
v26_0 26 254 dc 0.0
v27_0 27 255 dc 0.0
v28_0 28 256 dc 0.0
v29_0 29 257 dc 0.0
v30_0 30 258 dc 0.0
v31_0 31 259 dc 0.0
v32_0 32 260 dc 0.0
rc1_2to1 2 261 1e-05
cs1_2to1 261 1 0.022709950613374p
rp_2to1 2 1 55.052874804299
rl1_2to3 33 262 4.5707764709967
ls1_2to3 262 3 0.0099840045033175n
rl1_2to4 34 263 0.81990806623954
ls1_2to4 263 4 0.0019121977798303n
rc1_2to5 2 264 1e-05
cs1_2to5 264 5 4.0551794102895p
rp_2to5 2 5 0.2398483832036
rc1_2to6 2 265 1e-05
cs1_2to6 265 6 142.25535476535p
rp_2to6 2 6 0.081195869294773
rl1_2to7 35 266 0.027813484343015
ls1_2to7 266 7 4.714313216976e-05n
rl1_2to8 36 267 0.0095401065754837
ls1_2to8 267 8 3.2547475810405e-05n
rl1_2to9 37 268 0.0027055301932368
ls1_2to9 268 9 2.5121147106576e-05n
rl1_2to10 38 269 10.183205526566
ls1_2to10 269 10 0.00066760332467876n
rl1_2to11 39 270 1.4841134687625
ls1_2to11 270 11 0.0027505976901978n
rc1_2to12 2 271 1e-05
cs1_2to12 271 12 24.964681121352p
rp_2to12 2 12 0.35842710534024
rc1_2to13 2 272 1e-05
cs1_2to13 272 13 123.76220069235p
rp_2to13 2 13 0.11962758767993
rl1_2to14 40 273 0.041115922034354
ls1_2to14 273 14 4.3401209353191e-05n
rl1_2to15 41 274 0.014170411451887
ls1_2to15 274 15 2.4665002427688e-05n
rl1_2to16 42 275 0.0044377283478624
ls1_2to16 275 16 2.2315529829239e-05n
rc1_3to1 3 276 1e-05
cs1_3to1 276 1 0.0064730580322975p
rp_3to1 3 1 62.743373144645
rl1_3to4 43 277 5.47711821005
ls1_3to4 277 4 0.01739914038108n
rl1_3to5 44 278 1.0941980340492
ls1_3to5 278 5 0.0041479772577017n
rl1_3to6 45 279 0.30795421606978
ls1_3to6 279 6 0.0027594763829868n
rl1_3to7 46 280 0.10744523826476
ls1_3to7 280 7 0.00021099854512102n
rl1_3to8 47 281 0.037379114648727
ls1_3to8 281 8 0.00012059143658524n
rl1_3to9 48 282 0.012829217927753
ls1_3to9 282 9 6.5726164240924e-05n
rl1_3to10 49 283 23.633512884239
ls1_3to10 283 10 0.061239065810127n
rl1_3to11 50 284 12.632330631258
ls1_3to11 284 11 0.019114396558035n
rl1_3to12 51 285 1.7980838423889
ls1_3to12 285 12 0.0046820570474152n
rl1_3to13 52 286 0.47471640328827
ls1_3to13 286 13 0.0029169751023032n
rc1_3to14 3 287 1e-05
cs1_3to14 287 14 8.2224840090124p
rp_3to14 3 14 0.15819724234047
rl1_3to15 53 288 0.054049782205702
ls1_3to15 288 15 0.00011793200024701n
rl1_3to16 54 289 0.019091816932722
ls1_3to16 289 16 6.1629052176463e-05n
rc1_4to1 4 290 1e-05
cs1_4to1 290 1 0.0049708788137995p
rp_4to1 4 1 63.758196885758
rl1_4to5 55 291 6.0474297742881
ls1_4to5 291 5 0.021728794442956n
rl1_4to6 56 292 1.0913728386974
ls1_4to6 292 6 0.0041116580777319n
rl1_4to7 57 293 0.31411203829878
ls1_4to7 293 7 0.0035098553289707n
rl1_4to8 58 294 0.11096712444768
ls1_4to8 294 8 0.00065183721669702n
rl1_4to9 59 295 0.042081430975488
ls1_4to9 295 9 0.00019226465384724n
rl1_4to10 60 296 2.8272766034206
ls1_4to10 296 10 0.0054501565922518n
rs2_4to10 60 297 78.662634711701
ls2_4to10 297 10 54.861402418091n
rl1_4to11 61 298 22.418359973864
ls1_4to11 298 11 0.054017527768045n
rl1_4to12 62 299 12.285279738552
ls1_4to12 299 12 0.016026358965936n
rl1_4to13 63 300 1.9025048337655
ls1_4to13 300 13 0.0060517495920729n
rl1_4to14 64 301 0.48671459046189
ls1_4to14 301 14 0.0042386645825967n
rc1_4to15 4 302 1e-05
cs1_4to15 302 15 7.2123538308188p
rp_4to15 4 15 0.15980147609686
rc1_4to16 4 303 1e-05
cs1_4to16 303 16 82.018548612799p
rp_4to16 4 16 0.059807174731739
rc1_5to1 5 304 1e-05
cs1_5to1 304 1 0.0090085066416436p
rp_5to1 5 1 61.24134840515
rl1_5to6 65 305 5.5334874795765
ls1_5to6 305 6 0.016812570146982n
rl1_5to7 66 306 1.0575223364608
ls1_5to7 306 7 0.003623304078051n
rl1_5to8 67 307 0.31165140627942
ls1_5to8 307 8 0.0032960609614604n
rl1_5to9 68 308 0.11053544330595
ls1_5to9 308 9 0.0007543150619179n
rl1_5to10 69 309 0.66297555866631
ls1_5to10 309 10 0.0029288341501355n
rl1_5to11 70 310 2.9529527326667
ls1_5to11 310 11 0.005888896958691n
rs2_5to11 70 311 78.73016644146
ls2_5to11 311 11 55.721634121077n
rl1_5to12 71 312 25.274130714186
ls1_5to12 312 12 0.070730853635153n
rl1_5to13 72 313 12.294402306634
ls1_5to13 313 13 0.0152945763397n
rl1_5to14 73 314 1.8562017536388
ls1_5to14 314 14 0.0052415736236279n
rl1_5to15 74 315 0.46974739032455
ls1_5to15 315 15 0.0016962548200732n
rc1_5to16 5 316 1e-05
cs1_5to16 316 16 14.151727300032p
rp_5to16 5 16 0.16008667116934
rc1_6to1 6 317 1e-05
cs1_6to1 317 1 0.0054373734131884p
rp_6to1 6 1 63.405349773286
rl1_6to7 75 318 5.5800842444851
ls1_6to7 318 7 0.019016181357439n
rl1_6to8 76 319 1.0927255646091
ls1_6to8 319 8 0.0043799545581632n
rl1_6to9 77 320 0.32025257933671
ls1_6to9 320 9 0.0055771816816188n
rl1_6to10 78 321 0.20264539661748
ls1_6to10 321 10 0.0027436629241564n
rl1_6to11 79 322 0.6513932265888
ls1_6to11 322 11 0.0026498139777078n
rl1_6to12 80 323 2.9262041339747
ls1_6to12 323 12 0.0059348987936003n
rs2_6to12 80 324 77.144836738923
ls2_6to12 324 12 53.521041638913n
rl1_6to13 81 325 23.200703069106
ls1_6to13 325 13 0.057034559785324n
rl1_6to14 82 326 12.685418949222
ls1_6to14 326 14 0.021158444709377n
rl1_6to15 83 327 1.8455859068135
ls1_6to15 327 15 0.0053853464907585n
rl1_6to16 84 328 0.48785769832151
ls1_6to16 328 16 0.0042289913645955n
rc1_7to1 7 329 1e-05
cs1_7to1 329 1 0.0047951762826714p
rp_7to1 7 1 64.568489942435
rl1_7to8 85 330 5.9331228096839
ls1_7to8 330 8 0.0090808564433888n
rs2_7to8 85 331 204.96428709027
ls2_7to8 331 8 129.24839408891n
rl1_7to9 86 332 1.1292941935342
ls1_7to9 332 9 0.0026740642789721n
rs2_7to9 86 333 34.259326444637
ls2_7to9 333 9 27.365771949966n
rl1_7to10 87 334 0.072954154244444
ls1_7to10 334 10 0.00051901758967552n
rl1_7to11 88 335 0.20561459677425
ls1_7to11 335 11 0.0026139529611354n
rl1_7to12 89 336 0.66584436804716
ls1_7to12 336 12 0.0029028148211041n
rl1_7to13 90 337 2.8687068863596
ls1_7to13 337 13 0.0056197946952356n
rs2_7to13 90 338 79.521693954388
ls2_7to13 338 13 57.054473367365n
rl1_7to14 91 339 22.625107750035
ls1_7to14 339 14 0.054644152330224n
rl1_7to15 92 340 12.611852418067
ls1_7to15 340 15 0.016883013813522n
rl1_7to16 93 341 1.9345625011406
ls1_7to16 341 16 0.006106366097213n
rc1_8to1 8 342 1e-05
cs1_8to1 342 1 0.0081702364908477p
rp_8to1 8 1 62.221159035399
rl1_8to9 94 343 5.763391958284
ls1_8to9 343 9 0.0092399808850521n
rs2_8to9 94 344 185.41667265204
ls2_8to9 344 9 115.03238368477n
rl1_8to10 95 345 0.024858850279847
ls1_8to10 345 10 0.00010937606659599n
rl1_8to11 96 346 0.075200110242627
ls1_8to11 346 11 0.00062396418579027n
rl1_8to12 97 347 0.21244854168621
ls1_8to12 347 12 0.0037147892855716n
rl1_8to13 98 348 0.66896218290624
ls1_8to13 348 13 0.0029492286241133n
rl1_8to14 99 349 2.910188097808
ls1_8to14 349 14 0.0058846513885886n
rs2_8to14 99 350 76.408832468648
ls2_8to14 350 14 53.76789344094n
rl1_8to15 100 351 24.37141312484
ls1_8to15 351 15 0.066314092449275n
rl1_8to16 101 352 12.593543919797
ls1_8to16 352 16 0.013805050028611n
rc1_9to1 9 353 1e-05
cs1_9to1 353 1 0.007723812542579p
rp_9to1 9 1 61.698867586247
rl1_9to10 102 354 0.008115694243794
ls1_9to10 354 10 5.9706056804292e-05n
rl1_9to11 103 355 0.025738928752625
ls1_9to11 355 11 0.00012004698455434n
rl1_9to12 104 356 0.077775731293454
ls1_9to12 356 12 0.0011169581911561n
rl1_9to13 105 357 0.21375233642938
ls1_9to13 357 13 0.0042950748259696n
rl1_9to14 106 358 0.67871819076653
ls1_9to14 358 14 0.0017319090943815n
rs2_9to14 106 359 24.790224620912
ls2_9to14 359 14 13.484591097934n
rl1_9to15 107 360 3.0153186831549
ls1_9to15 360 15 0.0067129898487208n
rs2_9to15 107 361 66.03047990001
ls2_9to15 361 15 45.471600982101n
rl1_9to16 108 362 23.587083025226
ls1_9to16 362 16 0.074519430848421n
rc1_10to1 10 363 1e-05
cs1_10to1 363 1 0.0055351520797547p
rp_10to1 10 1 62.354424100289
rl1_10to11 109 364 5.8323594857209
ls1_10to11 364 11 0.01973924021548n
rl1_10to12 110 365 1.042158384415
ls1_10to12 365 12 0.003575885106908n
rl1_10to13 111 366 0.30564324291169
ls1_10to13 366 13 0.0033256391809023n
rl1_10to14 112 367 0.1064836979379
ls1_10to14 367 14 0.00039703625163842n
rl1_10to15 113 368 0.036226823666415
ls1_10to15 368 15 0.00010963567281598n
rl1_10to16 114 369 0.012397869705905
ls1_10to16 369 16 5.8571638481794e-05n
rc1_11to1 11 370 1e-05
cs1_11to1 370 1 0.0048208025624361p
rp_11to1 11 1 63.43096354788
rl1_11to12 115 371 5.4054065700146
ls1_11to12 371 12 0.015936267975915n
rl1_11to13 116 372 1.0706179698045
ls1_11to13 372 13 0.0039141344968398n
rl1_11to14 117 373 0.3105248168073
ls1_11to14 373 14 0.0031596026475636n
rl1_11to15 118 374 0.10731966841944
ls1_11to15 374 15 0.0001227892576036n
rl1_11to16 119 375 0.037516637691349
ls1_11to16 375 16 0.00011516049151949n
rc1_12to1 12 376 1e-05
cs1_12to1 376 1 0.0085684515128475p
rp_12to1 12 1 61.547529177675
rl1_12to13 120 377 5.7911750095015
ls1_12to13 377 13 0.02101620606954n
rl1_12to14 121 378 1.1043756410546
ls1_12to14 378 14 0.0043887549206535n
rl1_12to15 122 379 0.31336806223061
ls1_12to15 379 15 0.0034260930650563n
rl1_12to16 123 380 0.11164629213925
ls1_12to16 380 16 0.00058711894728338n
rc1_13to1 13 381 1e-05
cs1_13to1 381 1 0.0049052033759043p
rp_13to1 13 1 63.756760870664
rl1_13to14 124 382 5.7887101834028
ls1_13to14 382 14 0.019307513453654n
rl1_13to15 125 383 1.0716529640353
ls1_13to15 383 15 0.0037808172888378n
rl1_13to16 126 384 0.31781600828225
ls1_13to16 384 16 0.0036718147053263n
rc1_14to1 14 385 1e-05
cs1_14to1 385 1 0.0049337530691287p
rp_14to1 14 1 63.705010733893
rl1_14to15 127 386 5.5722104734831
ls1_14to15 386 15 0.016744613485289n
rl1_14to16 128 387 1.0924024077164
ls1_14to16 387 16 0.0039479787254241n
rc1_15to1 15 388 1e-05
cs1_15to1 388 1 0.0074609962349815p
rp_15to1 15 1 62.386878639183
rl1_15to16 129 389 5.9629240639603
ls1_15to16 389 16 0.01966599652423n
rc1_16to1 16 390 1e-05
cs1_16to1 390 1 0.0090702484046234p
rp_16to1 16 1 62.152013211255
rc1_18to17 18 391 1e-05
cs1_18to17 391 17 0.021694525809104p
rp_18to17 18 17 55.652617226743
rl1_18to19 130 392 4.7833367020265
ls1_18to19 392 19 0.011479906623241n
rl1_18to20 131 393 0.84266299072837
ls1_18to20 393 20 0.0020189708865579n
rl1_18to21 132 394 0.24544556490159
ls1_18to21 394 21 0.00016707203657462n
rc1_18to22 18 395 1e-05
cs1_18to22 395 22 38.049600660081p
rp_18to22 18 22 0.085522518493605
rl1_18to23 133 396 0.028257705415655
ls1_18to23 396 23 5.1371527348292e-05n
rl1_18to24 134 397 0.0097753873797185
ls1_18to24 397 24 3.5390429501168e-05n
rl1_18to25 135 398 0.002786991202182
ls1_18to25 398 25 2.5335597105923e-05n
rl1_18to26 136 399 10.715583847081
ls1_18to26 399 26 0.0081048479311411n
rl1_18to27 137 400 1.5246448138922
ls1_18to27 400 27 0.0030858351968548n
rc1_18to28 18 401 1e-05
cs1_18to28 401 28 18.930249391497p
rp_18to28 18 28 0.36692920801763
rc1_18to29 18 402 1e-05
cs1_18to29 402 29 126.24308649673p
rp_18to29 18 29 0.12073485611967
rl1_18to30 138 403 0.04304577587796
ls1_18to30 403 30 6.8314000150837e-05n
rl1_18to31 139 404 0.014760910447221
ls1_18to31 404 31 3.218952855409e-05n
rl1_18to32 140 405 0.0045455008590457
ls1_18to32 405 32 2.4242702818792e-05n
rc1_19to17 19 406 1e-05
cs1_19to17 406 17 0.0040979507853953p
rp_19to17 19 17 63.979024471582
rl1_19to20 141 407 5.4810838370727
ls1_19to20 407 20 0.015976604356902n
rl1_19to21 142 408 1.0875453970754
ls1_19to21 408 21 0.0039552030745397n
rl1_19to22 143 409 0.31719609515907
ls1_19to22 409 22 0.004748551985814n
rl1_19to23 144 410 0.10645841926142
ls1_19to23 410 23 2.988033655155e-05n
rl1_19to24 145 411 0.037134513063019
ls1_19to24 411 24 0.00011858356143666n
rl1_19to25 146 412 0.012698394633427
ls1_19to25 412 25 6.0228488329403e-05n
rl1_19to26 147 413 23.402004021416
ls1_19to26 413 26 0.054508812453068n
rl1_19to27 148 414 12.591564412649
ls1_19to27 414 27 0.019213537547286n
rl1_19to28 149 415 1.7863234730664
ls1_19to28 415 28 0.0044211120914756n
rl1_19to29 150 416 0.46588520451968
ls1_19to29 416 29 0.0011852560822052n
rl1_19to30 151 417 0.16087470388418
ls1_19to30 417 30 0.00038184095939732n
rc1_19to31 19 418 1e-05
cs1_19to31 418 31 115.28755423068p
rp_19to31 19 31 0.058119360166013
rl1_19to32 152 419 0.018933296352198
ls1_19to32 419 32 6.1125026537859e-05n
rc1_20to17 20 420 1e-05
cs1_20to17 420 17 0.0020932367039147p
rp_20to17 20 17 65.772866765019
rl1_20to21 153 421 6.0890388948827
ls1_20to21 421 21 0.022302992609449n
rl1_20to22 154 422 1.1620221308753
ls1_20to22 422 22 0.0028351373028725n
rs2_20to22 154 423 34.062322257045
ls2_20to22 423 22 26.979183411084n
rl1_20to23 155 424 0.31385548912773
ls1_20to23 424 23 0.0036324987813466n
rl1_20to24 156 425 0.11097907364222
ls1_20to24 425 24 0.0007864899679622n
rl1_20to25 157 426 0.041966771799232
ls1_20to25 426 25 9.531043550698e-05n
rl1_20to26 158 427 2.7772309901499
ls1_20to26 427 26 0.0047799424959444n
rs2_20to26 158 428 92.470105694787
ls2_20to26 428 26 63.584448744907n
rl1_20to27 159 429 22.322066598202
ls1_20to27 429 27 0.052631449999738n
rl1_20to28 160 430 12.4065656937
ls1_20to28 430 28 0.018219341522347n
rl1_20to29 161 431 1.8740465418611
ls1_20to29 431 29 0.0055549773903491n
rl1_20to30 162 432 0.50072839233771
ls1_20to30 432 30 0.0076431405806905n
rl1_20to31 163 433 0.1627452632471
ls1_20to31 433 31 0.00038680233126405n
rc1_20to32 20 434 1e-05
cs1_20to32 434 32 62.977316250069p
rp_20to32 20 32 0.059786369911815
rc1_21to17 21 435 1e-05
cs1_21to17 435 17 0.0093507024155968p
rp_21to17 21 17 61.13070861743
rl1_21to22 164 436 6.0652347926053
ls1_21to22 436 22 0.0098301672680765n
rs2_21to22 164 437 189.21111115978
ls2_21to22 437 22 118.23347891922n
rl1_21to23 165 438 1.0640200529346
ls1_21to23 438 23 0.0037544811488554n
rl1_21to24 166 439 0.31210592213861
ls1_21to24 439 24 0.0036328329910767n
rl1_21to25 167 440 0.11011930409589
ls1_21to25 440 25 0.00043939491379711n
rl1_21to26 168 441 0.6537559433489
ls1_21to26 441 26 0.0025954660829749n
rl1_21to27 169 442 2.9322042808006
ls1_21to27 442 27 0.0057523585918024n
rs2_21to27 169 443 80.00986695377
ls2_21to27 443 27 56.510126135665n
rl1_21to28 170 444 25.335776694416
ls1_21to28 444 28 0.069597169346499n
rl1_21to29 171 445 11.970485137216
ls1_21to29 445 29 0.010553261155799n
rl1_21to30 172 446 1.942492152568
ls1_21to30 446 30 0.007169730352712n
rl1_21to31 173 447 0.48050927336708
ls1_21to31 447 31 0.0035455906860294n
rc1_21to32 21 448 1e-05
cs1_21to32 448 32 9.1483469823938p
rp_21to32 21 32 0.15984802531917
rc1_22to17 22 449 1e-05
cs1_22to17 449 17 0.012464056347394p
rp_22to17 22 17 60.209907038618
rl1_22to23 174 450 5.1912697278032
ls1_22to23 450 23 0.011554943818135n
rl1_22to24 175 451 1.0375191214498
ls1_22to24 451 24 0.0031535801356728n
rl1_22to25 176 452 0.3066303112459
ls1_22to25 452 25 0.0014760695323775n
rl1_22to26 177 453 0.20731320079752
ls1_22to26 453 26 0.0034816308361724n
rl1_22to27 178 454 0.68562172187576
ls1_22to27 454 27 0.0017538097231848n
rs2_22to27 178 455 26.166582982564
ls2_22to27 455 27 12.14979854591n
rl1_22to28 179 456 3.1497470078395
ls1_22to28 456 28 0.0072072251682141n
rs2_22to28 179 457 66.254582232843
ls2_22to28 457 28 45.788217602591n
rl1_22to29 180 458 26.408553638154
ls1_22to29 458 29 0.081852674104936n
rl1_22to30 181 459 12.133000997934
ls1_22to30 459 30 0.015370050024938n
rl1_22to31 182 460 1.7868248530921
ls1_22to31 460 31 0.0039292646455602n
rc1_22to32 22 461 1e-05
cs1_22to32 461 32 0.76601782337465p
rp_22to32 22 32 0.4662614947082
rl1_23to17 183 462 64.61640100423
ls1_23to17 462 17 0.022920292717633n
rl1_23to24 184 463 5.876895552006
ls1_23to24 463 24 0.0091718935398184n
rs2_23to24 184 464 198.23599690585
ls2_23to24 464 24 125.40373098666n
rl1_23to25 185 465 1.0966814431528
ls1_23to25 465 25 0.0041498877674375n
rl1_23to26 186 466 0.071950771649096
ls1_23to26 466 26 0.00022622958927316n
rl1_23to27 187 467 0.2042661216075
ls1_23to27 467 27 0.0023578597892727n
rl1_23to28 188 468 0.66817595881371
ls1_23to28 468 28 0.0029279849940588n
rl1_23to29 189 469 2.9560392011312
ls1_23to29 469 29 0.0058336410223418n
rs2_23to29 189 470 80.415395221445
ls2_23to29 470 29 57.019919967646n
rl1_23to30 190 471 21.539257945471
ls1_23to30 471 30 0.039990355420503n
rl1_23to31 191 472 13.003626017128
ls1_23to31 472 31 0.023723554895002n
rl1_23to32 192 473 1.8921363838992
ls1_23to32 473 32 0.0057095614521659n
rc1_24to17 24 474 1e-05
cs1_24to17 474 17 0.0040729598926934p
rp_24to17 24 17 64.894426390273
rl1_24to25 193 475 5.4951150418127
ls1_24to25 475 25 0.016441768198408n
rl1_24to26 194 476 0.024613510804178
ls1_24to26 476 26 9.9964654322386e-05n
rl1_24to27 195 477 0.074861299566852
ls1_24to27 477 27 0.00060667228734876n
rl1_24to28 196 478 0.21272333638266
ls1_24to28 478 28 0.0038402147014638n
rl1_24to29 197 479 0.68094265873168
ls1_24to29 479 29 0.0031350917554485n
rl1_24to30 198 480 2.7825410504468
ls1_24to30 480 30 0.0051454148286459n
rs2_24to30 198 481 86.561949085166
ls2_24to30 481 30 61.494759249269n
rl1_24to31 199 482 23.051704010031
ls1_24to31 482 31 0.063276089835864n
rl1_24to32 200 483 12.145603704948
ls1_24to32 483 32 0.014136130279517n
rc1_25to17 25 484 1e-05
cs1_25to17 484 17 0.0025872358567055p
rp_25to17 25 17 63.371790692028
rl1_25to26 201 485 0.0080348048046001
ls1_25to26 485 26 5.2500622382984e-05n
rl1_25to27 202 486 0.025549395001484
ls1_25to27 486 27 0.00010800722468768n
rl1_25to28 203 487 0.077554461503487
ls1_25to28 487 28 0.00086845347736479n
rl1_25to29 204 488 0.21527249554961
ls1_25to29 488 29 0.0037673804603938n
rl1_25to30 205 489 0.64569512735998
ls1_25to30 489 30 0.0023227635943516n
rl1_25to31 206 490 2.8134479939312
ls1_25to31 490 31 0.0052384056624615n
rs2_25to31 206 491 83.62093647763
ls2_25to31 491 31 57.483710906825n
rl1_25to32 207 492 22.717769618
ls1_25to32 492 32 0.063468008490505n
rc1_26to17 26 493 1e-05
cs1_26to17 493 17 0.0052866275092728p
rp_26to17 26 17 63.304595690127
rl1_26to27 208 494 5.6886412779647
ls1_26to27 494 27 0.017051625087106n
rl1_26to28 209 495 1.025711154075
ls1_26to28 495 28 0.0030692434961921n
rl1_26to29 210 496 0.29856046148997
ls1_26to29 496 29 0.0014564534943413n
rl1_26to30 211 497 0.10771597313396
ls1_26to30 497 30 0.00052987873668443n
rl1_26to31 212 498 0.036482394978191
ls1_26to31 498 31 0.00010791458762474n
rl1_26to32 213 499 0.012261933549486
ls1_26to32 499 32 5.503102572465e-05n
rc1_27to17 27 500 1e-05
cs1_27to17 500 17 0.0024247650561559p
rp_27to17 27 17 65.290298765432
rl1_27to28 214 501 5.3606346231851
ls1_27to28 501 28 0.015580873337424n
rl1_27to29 215 502 1.0477395109317
ls1_27to29 502 29 0.0034511947631553n
rl1_27to30 216 503 0.31704767034438
ls1_27to30 503 30 0.0046813842024596n
rl1_27to31 217 504 0.10871824385598
ls1_27to31 504 31 0.00034461389714203n
rl1_27to32 218 505 0.03733854081386
ls1_27to32 505 32 0.00011570155816175n
rc1_28to17 28 506 1e-05
cs1_28to17 506 17 0.0084637072154121p
rp_28to17 28 17 61.973152800531
rl1_28to29 219 507 5.6718868164847
ls1_28to29 507 29 0.018548962062866n
rl1_28to30 220 508 1.1586122008336
ls1_28to30 508 30 0.0028317191073257n
rs2_28to30 220 509 34.598193928849
ls2_28to30 509 30 27.241143873145n
rl1_28to31 221 510 0.32008436874817
ls1_28to31 510 31 0.0044818516382859n
rl1_28to32 222 511 0.11158642051158
ls1_28to32 511 32 0.00062946735271935n
rc1_29to17 29 512 1e-05
cs1_29to17 512 17 0.012433147798463p
rp_29to17 29 17 60.075224853704
rl1_29to30 223 513 6.312470758803
ls1_29to30 513 30 0.010614406817802n
rs2_29to30 223 514 185.59643366615
ls2_29to30 514 30 118.61849175783n
rl1_29to31 224 515 1.1208733742112
ls1_29to31 515 31 0.0044761899884717n
rl1_29to32 225 516 0.32085726399312
ls1_29to32 516 32 0.0041073667978246n
rc1_30to17 30 517 1e-05
cs1_30to17 517 17 0.0021566516187104p
rp_30to17 30 17 64.844453196884
rl1_30to31 226 518 5.4678412354981
ls1_30to31 518 31 0.015201039341144n
rl1_30to32 227 519 1.0467029445858
ls1_30to32 519 32 0.0031054418214491n
rc1_31to17 31 520 1e-05
cs1_31to17 520 17 0.0048855120737811p
rp_31to17 31 17 63.996242229957
rl1_31to32 228 521 5.5206940704434
ls1_31to32 521 32 0.016653613011085n
rc1_32to17 32 522 1e-05
cs1_32to17 522 17 0.003609899103506p
rp_32to17 32 17 65.07684216048
rl1_1to0 229 523 88.100694676763
ls1_1to0 523 0 0.051696217462194n
rl1_2to0 230 524 116.21494333378
ls1_2to0 524 0 0.12327277036118n
rl1_3to0 231 525 119.0718859071
ls1_3to0 525 0 0.12758589350584n
rl1_4to0 232 526 119.09833970003
ls1_4to0 526 0 0.12203295140613n
rl1_5to0 233 527 119.84369306294
ls1_5to0 527 0 0.12574866202615n
rl1_6to0 234 528 119.38362820766
ls1_6to0 528 0 0.12723015273376n
rl1_7to0 235 529 121.04644388416
ls1_7to0 529 0 0.13276653400931n
rl1_8to0 236 530 117.97203817224
ls1_8to0 530 0 0.12698905767876n
rl1_9to0 237 531 88.158704601506
ls1_9to0 531 0 0.053003775239735n
rl1_10to0 238 532 117.61473864952
ls1_10to0 532 0 0.12819248651544n
rl1_11to0 239 533 118.52990831801
ls1_11to0 533 0 0.12519638816636n
rl1_12to0 240 534 119.492361132
ls1_12to0 534 0 0.12639292874386n
rl1_13to0 241 535 120.68814817841
ls1_13to0 535 0 0.13063771935565n
rl1_14to0 242 536 118.83782517391
ls1_14to0 536 0 0.12356576613396n
rl1_15to0 243 537 119.3871170943
ls1_15to0 537 0 0.12829271603443n
rl1_16to0 244 538 114.98644001556
ls1_16to0 538 0 0.12089686999882n
rl1_17to0 245 539 88.927886198789
ls1_17to0 539 0 0.053627064989602n
rl1_18to0 246 540 114.93720533743
ls1_18to0 540 0 0.12182205394054n
rl1_19to0 247 541 120.20101107939
ls1_19to0 541 0 0.12945085231735n
rl1_20to0 248 542 122.27785722655
ls1_20to0 542 0 0.14396200494478n
rl1_21to0 249 543 119.76911294946
ls1_21to0 543 0 0.12672409536333n
rl1_22to0 250 544 118.97916628268
ls1_22to0 544 0 0.12341384276195n
rl1_23to0 251 545 118.93694666975
ls1_23to0 545 0 0.12604523085331n
rl1_24to0 252 546 118.67544172726
ls1_24to0 546 0 0.12861667252027n
rl1_25to0 253 547 88.858568999943
ls1_25to0 547 0 0.055145413794501n
rl1_26to0 254 548 118.92282090963
ls1_26to0 548 0 0.13216547042228n
rl1_27to0 255 549 119.94526396104
ls1_27to0 549 0 0.12659964030924n
rl1_28to0 256 550 120.14065674023
ls1_28to0 550 0 0.12758447488816n
rl1_29to0 257 551 120.05058356148
ls1_29to0 551 0 0.13124446303421n
rl1_30to0 258 552 119.2684633506
ls1_30to0 552 0 0.11864590507933n
rl1_31to0 259 553 119.10515062712
ls1_31to0 553 0 0.13130906790983n
rl1_32to0 260 554 115.988007689
ls1_32to0 554 0 0.1208891272233n
.ends m16lines_port_lfws

