* begin ansoft header
* node 1 Diff1
* node 2 Comm1
* node 3 Diff2
* node 4 Comm2
* node 5 Diff3
* node 6 Comm3
* node 7 Diff4
* node 8 Comm4
* node 9 Diff5
* node 10 Comm5
* node 11 Diff6
* node 12 Comm6
* node 13 Diff7
* node 14 Comm7
* node 15 Diff8
* node 16 Comm8
* node 17 Diff9
* node 18 Comm9
* node 19 Diff10
* node 20 Comm10
* node 21 Diff11
* node 22 Comm11
* node 23 Diff12
* node 24 Comm12
* node 25 Diff13
* node 26 Comm13
* node 27 Diff14
* node 28 Comm14
* node 29 Diff15
* node 30 Comm15
* node 31 Diff16
* node 32 Comm16
* 
* created by ElectronicsDesktop
* end ansoft header

.subckt m16lines_HFSS_lfws 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 
rc1_2to1 2 33 1e-05
cs1_2to1 33 1 0.43205595593445p
rp_2to1 2 1 41635.171640727
rc1_2to3 2 34 1e-05
cs1_2to3 34 3 10.704112145101p
rp_2to3 2 3 985.10353990483
rc1_2to4 2 35 1e-05
cs1_2to4 35 4 97.11498735042p
rp_2to4 2 4 75.337710312183
rc1_2to5 2 36 1e-05
cs1_2to5 36 5 451.43885895712p
rp_2to5 2 5 13.425283416368
rc1_2to6 2 37 1e-05
cs1_2to6 37 6 2114.1579943766p
rp_2to6 2 6 1.6459888812735
rc1_2to7 2 38 1e-05
cs1_2to7 38 7 3454.5752894831p
rp_2to7 2 7 0.018861888842586
rl1_2to8 2 39 0.0029467681990766
ls1_2to8 39 8 0.0033975959512862n
rl1_2to9 2 40 0.0015455624637297
ls1_2to9 40 9 0.0067181541742473n
rc1_2to10 2 41 1e-05
cs1_2to10 41 10 3.436066138431p
rp_2to10 2 10 3790.8259417284
rc1_2to11 2 42 1e-05
cs1_2to11 42 11 45.396448298919p
rp_2to11 2 11 180.84986383776
rc1_2to12 2 43 1e-05
cs1_2to12 43 12 255.7000845964p
rp_2to12 2 12 24.62697279905
rc1_2to13 2 44 1e-05
cs1_2to13 44 13 1082.3791022065p
rp_2to13 2 13 4.3238576049882
rc1_2to14 2 45 1e-05
cs1_2to14 45 14 2288.5607468065p
rp_2to14 2 14 0.027929654751166
rl1_2to15 2 46 0.0038450109211658
ls1_2to15 46 15 0.00040269732022433n
rl1_2to16 2 47 0.0020330397534818
ls1_2to16 47 16 0.0059102036121897n
rc1_2to17 2 48 1e-05
cs1_2to17 48 17 21657.828522239p
rp_2to17 2 17 0.0018217288489344
rc1_2to18 2 49 1e-05
cs1_2to18 49 18 0.42752753571161p
rp_2to18 2 18 42643.658669234
rc1_2to19 2 50 1e-05
cs1_2to19 50 19 10.418878844298p
rp_2to19 2 19 1034.8070104834
rc1_2to20 2 51 1e-05
cs1_2to20 51 20 91.843058569027p
rp_2to20 2 20 83.508342516317
rc1_2to21 2 52 1e-05
cs1_2to21 52 21 414.8280961928p
rp_2to21 2 21 15.892566089028
rc1_2to22 2 53 1e-05
cs1_2to22 53 22 1797.1835491418p
rp_2to22 2 22 2.358651424328
rc1_2to23 2 54 1e-05
cs1_2to23 54 23 3449.8837413119p
rp_2to23 2 23 0.018844421968121
rl1_2to24 2 55 0.002933380221788
ls1_2to24 55 24 0.0030005155927925n
rl1_2to25 2 56 0.0015424514975678
ls1_2to25 56 25 0.0065702167821572n
rc1_2to26 2 57 1e-05
cs1_2to26 57 26 3.37407002087p
rp_2to26 2 26 3926.2308197522
rc1_2to27 2 58 1e-05
cs1_2to27 58 27 43.449204025868p
rp_2to27 2 27 196.2034390224
rc1_2to28 2 59 1e-05
cs1_2to28 59 28 237.96065043112p
rp_2to28 2 28 28.164031140873
rc1_2to29 2 60 1e-05
cs1_2to29 60 29 965.99542256993p
rp_2to29 2 29 5.459459799163
rc1_2to30 2 61 1e-05
cs1_2to30 61 30 8363.2089527947p
rp_2to30 2 30 0.10092067307685
rc1_2to31 2 62 1e-05
cs1_2to31 62 31 6452.8902911876p
rp_2to31 2 31 0.010426873686674
rl1_2to32 2 63 0.0020277307099189
ls1_2to32 63 32 0.0056833811554996n
rc1_3to1 3 64 1e-05
cs1_3to1 64 1 0.40626200861044p
rp_3to1 3 1 42788.726091277
rc1_3to4 3 65 1e-05
cs1_3to4 65 4 9.7165824665553p
rp_3to4 3 4 1047.4937478884
rc1_3to5 3 66 1e-05
cs1_3to5 66 5 84.972145850244p
rp_3to5 3 5 83.389800863712
rc1_3to6 3 67 1e-05
cs1_3to6 67 6 391.54039811379p
rp_3to6 3 6 14.722348019942
rc1_3to7 3 68 1e-05
cs1_3to7 68 7 1955.0469028997p
rp_3to7 3 7 1.5528118963162
rc1_3to8 3 69 1e-05
cs1_3to8 69 8 2907.2231021231p
rp_3to8 3 8 0.022922802827525
rl1_3to9 3 70 0.0036422489927194
ls1_3to9 70 9 0.0049556755629048n
rc1_3to10 3 71 1e-05
cs1_3to10 71 10 1.6466303231992p
rp_3to10 3 10 8426.1950378722
rc1_3to11 3 72 1e-05
cs1_3to11 72 11 3.1668489949587p
rp_3to11 3 11 3961.2471300691
rc1_3to12 3 73 1e-05
cs1_3to12 73 12 40.244460103914p
rp_3to12 3 12 197.79538634935
rc1_3to13 3 74 1e-05
cs1_3to13 74 13 221.37720420217p
rp_3to13 3 13 28.124551649337
rc1_3to14 3 75 1e-05
cs1_3to14 75 14 957.70502816412p
rp_3to14 3 14 4.5798927732915
rc1_3to15 3 76 1e-05
cs1_3to15 76 15 1926.2533976979p
rp_3to15 3 15 0.033939272903525
rl1_3to16 3 77 0.004747608988421
ls1_3to16 77 16 0.0015380722916525n
rl1_3to17 3 78 6.2403854797824
ls1_3to17 78 17 0.15899288028969n
rc1_3to18 3 79 1e-05
cs1_3to18 79 18 10.392755320568p
rp_3to18 3 18 1039.8200608731
rc1_3to19 3 80 1e-05
cs1_3to19 80 19 0.40187521374663p
rp_3to19 3 19 43823.053153259
rc1_3to20 3 81 1e-05
cs1_3to20 81 20 9.4466847126922p
rp_3to20 3 20 1101.9805751639
rc1_3to21 3 82 1e-05
cs1_3to21 82 21 80.212141039128p
rp_3to21 3 21 92.685590683915
rc1_3to22 3 83 1e-05
cs1_3to22 83 22 358.44500916496p
rp_3to22 3 22 17.554021908527
rc1_3to23 3 84 1e-05
cs1_3to23 84 23 1621.7665337684p
rp_3to23 3 23 2.375106240214
rc1_3to24 3 85 1e-05
cs1_3to24 85 24 2903.0095920882p
rp_3to24 3 24 0.022900415374612
rl1_3to25 3 86 0.0036079318818942
ls1_3to25 86 25 0.0044429638554738n
rc1_3to26 3 87 1e-05
cs1_3to26 87 26 1.6207845225582p
rp_3to26 3 26 8668.9748014713
rc1_3to27 3 88 1e-05
cs1_3to27 88 27 3.1072556606469p
rp_3to27 3 27 4106.2084529174
rc1_3to28 3 89 1e-05
cs1_3to28 89 28 38.455758990668p
rp_3to28 3 28 215.11939297182
rc1_3to29 3 90 1e-05
cs1_3to29 90 29 205.51262965597p
rp_3to29 3 29 32.396125490162
rc1_3to30 3 91 1e-05
cs1_3to30 91 30 846.73343411801p
rp_3to30 3 30 5.9212970043915
rc1_3to31 3 92 1e-05
cs1_3to31 92 31 1923.6300760046p
rp_3to31 3 31 0.033904845986179
rl1_3to32 3 93 0.0047027197919298
ls1_3to32 93 32 0.00080436935216836n
rc1_4to1 4 94 1e-05
cs1_4to1 94 1 0.40573780066987p
rp_4to1 4 1 42859.340391007
rc1_4to5 4 95 1e-05
cs1_4to5 95 5 9.6995375455962p
rp_4to5 4 5 1048.7492892978
rc1_4to6 4 96 1e-05
cs1_4to6 96 6 84.813098986161p
rp_4to6 4 6 83.373624193408
rc1_4to7 4 97 1e-05
cs1_4to7 97 7 390.71670551564p
rp_4to7 4 7 14.724250421605
rc1_4to8 4 98 1e-05
cs1_4to8 98 8 1955.4919953838p
rp_4to8 4 8 1.5430062672214
rc1_4to9 4 99 1e-05
cs1_4to9 99 9 2842.1614736203p
rp_4to9 4 9 0.0234273267254
rc1_4to10 4 100 1e-05
cs1_4to10 100 10 25.739138398345p
rp_4to10 4 10 332.69220739141
rc1_4to11 4 101 1e-05
cs1_4to11 101 11 1.6401486963428p
rp_4to11 4 11 8439.9264168274
rc1_4to12 4 102 1e-05
cs1_4to12 102 12 3.1626992318096p
rp_4to12 4 12 3964.2882428467
rc1_4to13 4 103 1e-05
cs1_4to13 103 13 40.183998451163p
rp_4to13 4 13 197.79304832058
rc1_4to14 4 104 1e-05
cs1_4to14 104 14 221.01800934964p
rp_4to14 4 14 28.152523220485
rc1_4to15 4 105 1e-05
cs1_4to15 105 15 956.57879813147p
rp_4to15 4 15 4.5677937630222
rc1_4to16 4 106 1e-05
cs1_4to16 106 16 1907.8997544069p
rp_4to16 4 16 0.034288455496019
rl1_4to17 4 107 0.79720246589297
ls1_4to17 107 17 0.07599622173417n
rc1_4to18 4 108 1e-05
cs1_4to18 108 18 91.134400010341p
rp_4to18 4 18 84.741361914476
rc1_4to19 4 109 1e-05
cs1_4to19 109 19 9.4464968075332p
rp_4to19 4 19 1101.9618297453
rc1_4to20 4 110 1e-05
cs1_4to20 110 20 0.40135872772945p
rp_4to20 4 20 43892.285737762
rc1_4to21 4 111 1e-05
cs1_4to21 111 21 9.4300883443396p
rp_4to21 4 21 1103.2080175141
rc1_4to22 4 112 1e-05
cs1_4to22 112 22 80.06150511997p
rp_4to22 4 22 92.634870897934
rc1_4to23 4 113 1e-05
cs1_4to23 113 23 357.76352846624p
rp_4to23 4 23 17.521198723898
rc1_4to24 4 114 1e-05
cs1_4to24 114 24 1622.5494491963p
rp_4to24 4 24 2.3508720440316
rc1_4to25 4 115 1e-05
cs1_4to25 115 25 2838.2697223067p
rp_4to25 4 25 0.023405481219501
rc1_4to26 4 116 1e-05
cs1_4to26 116 26 24.731996020343p
rp_4to26 4 26 357.0319864697
rc1_4to27 4 117 1e-05
cs1_4to27 117 27 1.6143828418828p
rp_4to27 4 27 8682.3991068815
rc1_4to28 4 118 1e-05
cs1_4to28 118 28 3.1031492523155p
rp_4to28 4 28 4109.1663161836
rc1_4to29 4 119 1e-05
cs1_4to29 119 29 38.397424269601p
rp_4to29 4 29 215.06378253037
rc1_4to30 4 120 1e-05
cs1_4to30 120 30 205.16679306571p
rp_4to30 4 30 32.497242092935
rc1_4to31 4 121 1e-05
cs1_4to31 121 31 845.95647981157p
rp_4to31 4 31 5.8892372523815
rc1_4to32 4 122 1e-05
cs1_4to32 122 32 1905.3604530749p
rp_4to32 4 32 0.034256949545561
rc1_5to1 5 123 1e-05
cs1_5to1 123 1 0.40583130126867p
rp_5to1 5 1 42835.618308236
rc1_5to6 5 124 1e-05
cs1_5to6 124 6 9.711774124449p
rp_5to6 5 6 1046.4560755824
rc1_5to7 5 125 1e-05
cs1_5to7 125 7 84.842847703765p
rp_5to7 5 7 83.364201905084
rc1_5to8 5 126 1e-05
cs1_5to8 126 8 390.12516627558p
rp_5to8 5 8 14.776985124348
rc1_5to9 5 127 1e-05
cs1_5to9 127 9 1863.414571598p
rp_5to9 5 9 1.6968067071792
rc1_5to10 5 128 1e-05
cs1_5to10 128 10 163.09688918896p
rp_5to10 5 10 39.673477585148
rc1_5to11 5 129 1e-05
cs1_5to11 129 11 25.56599023728p
rp_5to11 5 11 333.53351721979
rc1_5to12 5 130 1e-05
cs1_5to12 130 12 1.6405649561555p
rp_5to12 5 12 8436.2259322449
rc1_5to13 5 131 1e-05
cs1_5to13 131 13 3.1669579983978p
rp_5to13 5 13 3954.7333742574
rc1_5to14 5 132 1e-05
cs1_5to14 132 14 40.228916104078p
rp_5to14 5 14 197.51488594115
rc1_5to15 5 133 1e-05
cs1_5to15 133 15 220.88868384126p
rp_5to15 5 15 28.154730970825
rc1_5to16 5 134 1e-05
cs1_5to16 134 16 944.89306077379p
rp_5to16 5 16 4.67407866527
rl1_5to17 5 135 -0.0061322999835198
ls1_5to17 135 17 -0.000440431014487n
rc1_5to18 5 136 1e-05
cs1_5to18 136 18 409.16144454524p
rp_5to18 5 18 16.352832408718
rc1_5to19 5 137 1e-05
cs1_5to19 137 19 80.208378927998p
rp_5to19 5 19 92.679777604764
rc1_5to20 5 138 1e-05
cs1_5to20 138 20 9.4300773242707p
rp_5to20 5 20 1103.2191683186
rc1_5to21 5 139 1e-05
cs1_5to21 139 21 0.40144924729133p
rp_5to21 5 21 43869.938980465
rc1_5to22 5 140 1e-05
cs1_5to22 140 22 9.4416406912977p
rp_5to22 5 22 1100.9514700177
rc1_5to23 5 141 1e-05
cs1_5to23 141 23 80.08816018328p
rp_5to23 5 23 92.63746295524
rc1_5to24 5 142 1e-05
cs1_5to24 142 24 357.20376204571p
rp_5to24 5 24 17.620351977085
rc1_5to25 5 143 1e-05
cs1_5to25 143 25 1558.3376611267p
rp_5to25 5 25 2.5343983782507
rc1_5to26 5 144 1e-05
cs1_5to26 144 26 152.1094119881p
rp_5to26 5 26 45.088390673496
rc1_5to27 5 145 1e-05
cs1_5to27 145 27 24.567983187666p
rp_5to27 5 27 357.84664813765
rc1_5to28 5 146 1e-05
cs1_5to28 146 28 1.6147970916736p
rp_5to28 5 28 8678.1391009698
rc1_5to29 5 147 1e-05
cs1_5to29 147 29 3.1072615905695p
rp_5to29 5 29 4099.9281812322
rc1_5to30 5 148 1e-05
cs1_5to30 148 30 38.438338570442p
rp_5to30 5 30 214.76456738468
rc1_5to31 5 149 1e-05
cs1_5to31 149 31 205.04999884796p
rp_5to31 5 31 32.402919225425
rc1_5to32 5 150 1e-05
cs1_5to32 150 32 836.36669235715p
rp_5to32 5 32 6.0140862301377
rc1_6to1 6 151 1e-05
cs1_6to1 151 1 0.40600532741774p
rp_6to1 6 1 42803.139741081
rc1_6to7 6 152 1e-05
cs1_6to7 152 7 9.7128034628209p
rp_6to7 6 7 1046.5189226564
rc1_6to8 6 153 1e-05
cs1_6to8 153 8 84.80940284473p
rp_6to8 6 8 83.511702822299
rc1_6to9 6 154 1e-05
cs1_6to9 154 9 381.6810636966p
rp_6to9 6 9 15.068358009142
rc1_6to10 6 155 1e-05
cs1_6to10 155 10 698.16383546957p
rp_6to10 6 10 7.1759536891439
rc1_6to11 6 156 1e-05
cs1_6to11 156 11 161.66963928979p
rp_6to11 6 11 39.798328323699
rc1_6to12 6 157 1e-05
cs1_6to12 157 12 25.597955213121p
rp_6to12 6 12 332.86926647655
rc1_6to13 6 158 1e-05
cs1_6to13 158 13 1.6400247164688p
rp_6to13 6 13 8440.0020268762
rc1_6to14 6 159 1e-05
cs1_6to14 159 14 3.1682316612317p
rp_6to14 6 14 3953.2600011963
rc1_6to15 6 160 1e-05
cs1_6to15 160 15 40.196106658385p
rp_6to15 6 15 197.88943546491
rc1_6to16 6 161 1e-05
cs1_6to16 161 16 219.61921763974p
rp_6to16 6 16 27.851030339379
rl1_6to17 6 162 -0.0015999304287326
ls1_6to17 162 17 -5.9902295046993e-05n
rc1_6to18 6 163 1e-05
cs1_6to18 163 18 1744.1818554784p
rp_6to18 6 18 2.5269164613694
rc1_6to19 6 164 1e-05
cs1_6to19 164 19 358.40077234109p
rp_6to19 6 19 17.547779833536
rc1_6to20 6 165 1e-05
cs1_6to20 165 20 80.057941465185p
rp_6to20 6 20 92.663433080163
rc1_6to21 6 166 1e-05
cs1_6to21 166 21 9.441596046784p
rp_6to21 6 21 1100.9651513898
rc1_6to22 6 167 1e-05
cs1_6to22 167 22 0.40161994633705p
rp_6to22 6 22 43836.501671041
rc1_6to23 6 168 1e-05
cs1_6to23 168 23 9.442726004011p
rp_6to23 6 23 1100.9223810914
rc1_6to24 6 169 1e-05
cs1_6to24 169 24 80.054736822881p
rp_6to24 6 24 92.813681984384
rc1_6to25 6 170 1e-05
cs1_6to25 170 25 349.83954918354p
rp_6to25 6 25 18.015921063857
rc1_6to26 6 171 1e-05
cs1_6to26 171 26 626.17648357788p
rp_6to26 6 26 8.9513928448468
rc1_6to27 6 172 1e-05
cs1_6to27 172 27 150.81212439755p
rp_6to27 6 27 45.215679518399
rc1_6to28 6 173 1e-05
cs1_6to28 173 28 24.597572927145p
rp_6to28 6 28 357.18754399852
rc1_6to29 6 174 1e-05
cs1_6to29 174 29 1.6142609855823p
rp_6to29 6 29 8682.3523317272
rc1_6to30 6 175 1e-05
cs1_6to30 175 30 3.1085015461342p
rp_6to30 6 30 4098.4354233996
rc1_6to31 6 176 1e-05
cs1_6to31 176 31 38.407527390131p
rp_6to31 6 31 215.17791849147
rc1_6to32 6 177 1e-05
cs1_6to32 177 32 203.8944678765p
rp_6to32 6 32 32.01538626177
rc1_7to1 7 178 1e-05
cs1_7to1 178 1 0.40583794000295p
rp_7to1 7 1 42851.596433086
rc1_7to8 7 179 1e-05
cs1_7to8 179 8 9.701698621956p
rp_7to8 7 8 1048.2753077003
rc1_7to9 7 180 1e-05
cs1_7to9 180 9 83.355597022358p
rp_7to9 7 9 85.142083312703
rc1_7to10 7 181 1e-05
cs1_7to10 181 10 5967.8282254613p
rp_7to10 7 10 0.11966308567281
rc1_7to11 7 182 1e-05
cs1_7to11 182 11 694.5321436218p
rp_7to11 7 11 7.1206559237182
rc1_7to12 7 183 1e-05
cs1_7to12 183 12 161.74811198846p
rp_7to12 7 12 39.7486122354
rc1_7to13 7 184 1e-05
cs1_7to13 184 13 25.582665101762p
rp_7to13 7 13 333.14802111994
rc1_7to14 7 185 1e-05
cs1_7to14 185 14 1.6398503238652p
rp_7to14 7 14 8439.5362421019
rc1_7to15 7 186 1e-05
cs1_7to15 186 15 3.1608837684056p
rp_7to15 7 15 3967.3686553408
rc1_7to16 7 187 1e-05
cs1_7to16 187 16 40.036943092265p
rp_7to16 7 16 198.55871343349
rc1_7to17 7 188 1e-05
cs1_7to17 188 17 3269269.5913312p
rp_7to17 7 17 100000
rc1_7to18 7 189 1e-05
cs1_7to18 189 18 3448.7300499146p
rp_7to18 7 18 0.018925023171117
rc1_7to19 7 190 1e-05
cs1_7to19 190 19 1622.4409944559p
rp_7to19 7 19 2.3685625777489
rc1_7to20 7 191 1e-05
cs1_7to20 191 20 357.73909877484p
rp_7to20 7 20 17.535023914429
rc1_7to21 7 192 1e-05
cs1_7to21 192 21 80.087377375074p
rp_7to21 7 21 92.629305322202
rc1_7to22 7 193 1e-05
cs1_7to22 193 22 9.4427503943079p
rp_7to22 7 22 1100.9083020056
rc1_7to23 7 194 1e-05
cs1_7to23 194 23 0.40145708609785p
rp_7to23 7 23 43886.300602739
rc1_7to24 7 195 1e-05
cs1_7to24 195 24 9.4319988571024p
rp_7to24 7 24 1102.8609302053
rc1_7to25 7 196 1e-05
cs1_7to25 196 25 78.697463433819p
rp_7to25 7 25 94.526075262209
rc1_7to26 7 197 1e-05
cs1_7to26 197 26 4049.595210578p
rp_7to26 7 26 0.46185187377003
rc1_7to27 7 198 1e-05
cs1_7to27 198 27 623.08965165691p
rp_7to27 7 27 8.8689876914712
rc1_7to28 7 199 1e-05
cs1_7to28 199 28 150.89619095984p
rp_7to28 7 28 45.144871640653
rc1_7to29 7 200 1e-05
cs1_7to29 200 29 24.583833567574p
rp_7to29 7 29 357.41446002895
rc1_7to30 7 201 1e-05
cs1_7to30 201 30 1.6140990143405p
rp_7to30 7 30 8681.2220851641
rc1_7to31 7 202 1e-05
cs1_7to31 202 31 3.1013663057303p
rp_7to31 7 31 4112.4363275106
rc1_7to32 7 203 1e-05
cs1_7to32 203 32 38.255611069629p
rp_7to32 7 32 215.86112591294
rc1_8to1 8 204 1e-05
cs1_8to1 204 1 0.40561162028453p
rp_8to1 8 1 42861.855355587
rc1_8to9 8 205 1e-05
cs1_8to9 205 9 9.6155987226392p
rp_8to9 8 9 1055.7354524038
rc1_8to10 8 206 1e-05
cs1_8to10 206 10 4431.7790821574p
rp_8to10 8 10 0.015358598778474
rc1_8to11 8 207 1e-05
cs1_8to11 207 11 5931.4272753237p
rp_8to11 8 11 0.094643579145449
rc1_8to12 8 208 1e-05
cs1_8to12 208 12 693.6940518357p
rp_8to12 8 12 7.1385981848571
rc1_8to13 8 209 1e-05
cs1_8to13 209 13 161.49570959353p
rp_8to13 8 13 39.868483654363
rc1_8to14 8 210 1e-05
cs1_8to14 210 14 25.562069577568p
rp_8to14 8 14 333.56072941881
rc1_8to15 8 211 1e-05
cs1_8to15 211 15 1.6427857888779p
rp_8to15 8 15 8420.1521585334
rc1_8to16 8 212 1e-05
cs1_8to16 212 16 3.1613946518646p
rp_8to16 8 16 3963.0760493396
rl1_8to17 8 213 -0.00084147399420337
ls1_8to17 213 17 -0.00032002197557139n
rl1_8to18 8 214 0.002905321958686
ls1_8to18 214 18 0.0028540975217764n
rc1_8to19 8 215 1e-05
cs1_8to19 215 19 2902.9157848262p
rp_8to19 8 19 0.022666646630452
rc1_8to20 8 216 1e-05
cs1_8to20 216 20 1621.5417163216p
rp_8to20 8 20 2.3583940596954
rc1_8to21 8 217 1e-05
cs1_8to21 217 21 357.16713962125p
rp_8to21 8 21 17.621829808842
rc1_8to22 8 218 1e-05
cs1_8to22 218 22 80.055677026034p
rp_8to22 8 22 92.812147652312
rc1_8to23 8 219 1e-05
cs1_8to23 219 23 9.4319801796449p
rp_8to23 8 23 1102.8653684653
rc1_8to24 8 220 1e-05
cs1_8to24 220 24 0.40123161763682p
rp_8to24 8 24 43893.895514121
rc1_8to25 8 221 1e-05
cs1_8to25 221 25 9.3470387406011p
rp_8to25 8 25 1110.5113823033
rc1_8to26 8 222 1e-05
cs1_8to26 222 26 4425.0504609505p
rp_8to26 8 26 0.015341141437028
rc1_8to27 8 223 1e-05
cs1_8to27 223 27 4205.5260743125p
rp_8to27 8 27 0.4067303171706
rc1_8to28 8 224 1e-05
cs1_8to28 224 28 622.33129217298p
rp_8to28 8 28 8.8960380875909
rc1_8to29 8 225 1e-05
cs1_8to29 225 29 150.66567571827p
rp_8to29 8 29 45.28020048717
rc1_8to30 8 226 1e-05
cs1_8to30 226 30 24.563895617107p
rp_8to30 8 30 357.89629292023
rc1_8to31 8 227 1e-05
cs1_8to31 227 31 1.6169539503781p
rp_8to31 8 31 8662.6921206785
rc1_8to32 8 228 1e-05
cs1_8to32 228 32 3.1017193721174p
rp_8to32 8 32 4107.9423979003
rc1_9to1 9 229 1e-05
cs1_9to1 229 1 0.40382021005576p
rp_9to1 9 1 42943.828160249
rl1_9to10 9 230 0.0026850496054009
ls1_9to10 230 10 0.006932350365818n
rc1_9to11 9 231 1e-05
cs1_9to11 231 11 4287.5353265642p
rp_9to11 9 11 0.015925656591591
rc1_9to12 9 232 1e-05
cs1_9to12 232 12 5750.7971534006p
rp_9to12 9 12 0.13042053633246
rc1_9to13 9 233 1e-05
cs1_9to13 233 13 673.8682659522p
rp_9to13 9 13 7.6257792931041
rc1_9to14 9 234 1e-05
cs1_9to14 234 14 158.47215877371p
rp_9to14 9 14 40.939739082727
rc1_9to15 9 235 1e-05
cs1_9to15 235 15 25.301912831441p
rp_9to15 9 15 336.85547225712
rc1_9to16 9 236 1e-05
cs1_9to16 236 16 1.6299223642184p
rp_9to16 9 16 8469.8681473436
rc1_9to17 9 237 1e-05
cs1_9to17 237 17 18108227.331404p
rp_9to17 9 17 100000
rl1_9to18 9 238 0.0015587098151223
ls1_9to18 238 18 0.0064579400829072n
rl1_9to19 9 239 0.003615742664456
ls1_9to19 239 19 0.004433931369869n
rc1_9to20 9 240 1e-05
cs1_9to20 240 20 2838.267936495p
rp_9to20 9 20 0.023397774705907
rc1_9to21 9 241 1e-05
cs1_9to21 241 21 1555.7488157209p
rp_9to21 9 21 2.5412588777892
rc1_9to22 9 242 1e-05
cs1_9to22 242 22 349.77333719853p
rp_9to22 9 22 18.016880421941
rc1_9to23 9 243 1e-05
cs1_9to23 243 23 78.691629514145p
rp_9to23 9 23 94.534493052011
rc1_9to24 9 244 1e-05
cs1_9to24 244 24 9.3469715434746p
rp_9to24 9 24 1110.4981671739
rc1_9to25 9 245 1e-05
cs1_9to25 245 25 0.39943950901649p
rp_9to25 9 25 43974.344679034
rl1_9to26 9 246 0.0026731194591077
ls1_9to26 246 26 0.0065522875843943n
rc1_9to27 9 247 1e-05
cs1_9to27 247 27 4281.1577838526p
rp_9to27 9 27 0.015912945689185
rc1_9to28 9 248 1e-05
cs1_9to28 248 28 3899.8969626337p
rp_9to28 9 28 0.48529484290298
rc1_9to29 9 249 1e-05
cs1_9to29 249 29 605.58343097377p
rp_9to29 9 29 9.4757904140238
rc1_9to30 9 250 1e-05
cs1_9to30 250 30 147.88387029941p
rp_9to30 9 30 46.436905975363
rc1_9to31 9 251 1e-05
cs1_9to31 251 31 24.310317803266p
rp_9to31 9 31 361.37522214039
rc1_9to32 9 252 1e-05
cs1_9to32 252 32 1.6041631597542p
rp_9to32 9 32 8713.0718214109
rc1_10to1 10 253 1e-05
cs1_10to1 253 1 0.40636350388921p
rp_10to1 10 1 42897.437550603
rc1_10to11 10 254 1e-05
cs1_10to11 254 11 9.7534415289756p
rp_10to11 10 11 1046.6648534744
rc1_10to12 10 255 1e-05
cs1_10to12 255 12 85.513355124921p
rp_10to12 10 12 83.211014812159
rc1_10to13 10 256 1e-05
cs1_10to13 256 13 393.70921043916p
rp_10to13 10 13 14.766425448409
rc1_10to14 10 257 1e-05
cs1_10to14 257 14 1943.2012129304p
rp_10to14 10 14 1.6002712212527
rc1_10to15 10 258 1e-05
cs1_10to15 258 15 2939.9832022806p
rp_10to15 10 15 0.022612629642644
rl1_10to16 10 259 0.0035526857876504
ls1_10to16 259 16 0.0048444994739226n
rc1_10to17 10 260 1e-05
cs1_10to17 260 17 35885.17206559p
rp_10to17 10 17 100000
rc1_10to18 10 261 1e-05
cs1_10to18 261 18 3.3703726472357p
rp_10to18 10 18 3935.1177286154
rc1_10to19 10 262 1e-05
cs1_10to19 262 19 1.6208390348434p
rp_10to19 10 19 8668.3734289474
rc1_10to20 10 263 1e-05
cs1_10to20 263 20 24.7387562641p
rp_10to20 10 20 356.86694857703
rc1_10to21 10 264 1e-05
cs1_10to21 264 21 152.22085292265p
rp_10to21 10 21 45.021500739638
rc1_10to22 10 265 1e-05
cs1_10to22 265 22 627.32235227554p
rp_10to22 10 22 8.9125581959742
rc1_10to23 10 266 1e-05
cs1_10to23 266 23 4084.7808183994p
rp_10to23 10 23 0.45075916415057
rc1_10to24 10 267 1e-05
cs1_10to24 267 24 4425.5685475435p
rp_10to24 10 24 0.015372519766107
rl1_10to25 10 268 0.0026575330206623
ls1_10to25 268 25 0.0066010625242719n
rc1_10to26 10 269 1e-05
cs1_10to26 269 26 0.40198870333404p
rp_10to26 10 26 43932.429832926
rc1_10to27 10 270 1e-05
cs1_10to27 270 27 9.4835635734014p
rp_10to27 10 27 1100.8882411551
rc1_10to28 10 271 1e-05
cs1_10to28 271 28 80.746149979743p
rp_10to28 10 28 92.429317124211
rc1_10to29 10 272 1e-05
cs1_10to29 272 29 360.77901226245p
rp_10to29 10 29 17.569635950273
rc1_10to30 10 273 1e-05
cs1_10to30 273 30 1621.4491369896p
rp_10to30 10 30 2.4060254426134
rc1_10to31 10 274 1e-05
cs1_10to31 274 31 2935.8742229572p
rp_10to31 10 31 0.022589584017435
rl1_10to32 10 275 0.0035295613646958
ls1_10to32 275 32 0.0043566918654198n
rc1_11to1 11 276 1e-05
cs1_11to1 276 1 0.40576593477687p
rp_11to1 11 1 42863.055081532
rc1_11to12 11 277 1e-05
cs1_11to12 277 12 9.7015863390109p
rp_11to12 11 12 1048.4228335704
rc1_11to13 11 278 1e-05
cs1_11to13 278 13 84.807776297973p
rp_11to13 11 13 83.407298179659
rc1_11to14 11 279 1e-05
cs1_11to14 279 14 390.99093972337p
rp_11to14 11 14 14.7129926232
rc1_11to15 11 280 1e-05
cs1_11to15 280 15 1960.9896883342p
rp_11to15 11 15 1.5340768034505
rc1_11to16 11 281 1e-05
cs1_11to16 281 16 2881.8339772447p
rp_11to16 11 16 0.02312766686465
rc1_11to17 11 282 1e-05
cs1_11to17 282 17 116097.14514493p
rp_11to17 11 17 100000
rc1_11to18 11 283 1e-05
cs1_11to18 283 18 43.211981684193p
rp_11to18 11 18 198.28052055293
rc1_11to19 11 284 1e-05
cs1_11to19 284 19 3.1072297223142p
rp_11to19 11 19 4106.1941326705
rc1_11to20 11 285 1e-05
cs1_11to20 285 20 1.6143837021878p
rp_11to20 11 20 8682.3706612232
rc1_11to21 11 286 1e-05
cs1_11to21 286 21 24.568157597748p
rp_11to21 11 21 357.82503351449
rc1_11to22 11 287 1e-05
cs1_11to22 287 22 150.82602616511p
rp_11to22 11 22 45.194765902662
rc1_11to23 11 288 1e-05
cs1_11to23 288 23 623.16866381565p
rp_11to23 11 23 8.8624257726193
rc1_11to24 11 289 1e-05
cs1_11to24 289 24 4212.9197336488p
rp_11to24 11 24 0.40343286395758
rc1_11to25 11 290 1e-05
cs1_11to25 290 25 4281.2575105763p
rp_11to25 11 25 0.015833537447251
rc1_11to26 11 291 1e-05
cs1_11to26 291 26 9.4821953641238p
rp_11to26 11 26 1101.1698910978
rc1_11to27 11 292 1e-05
cs1_11to27 292 27 0.4013871616437p
rp_11to27 11 27 43897.357756381
rc1_11to28 11 293 1e-05
cs1_11to28 293 28 9.4319728266126p
rp_11to28 11 28 1102.9379465719
rc1_11to29 11 294 1e-05
cs1_11to29 294 29 80.057268422579p
rp_11to29 11 29 92.676487059669
rc1_11to30 11 295 1e-05
cs1_11to30 295 30 357.98274226349p
rp_11to30 11 30 17.502917516041
rc1_11to31 11 296 1e-05
cs1_11to31 296 31 1626.0356351512p
rp_11to31 11 31 2.3414400322683
rc1_11to32 11 297 1e-05
cs1_11to32 297 32 2877.7848039898p
rp_11to32 11 32 0.023106941937176
rc1_12to1 12 298 1e-05
cs1_12to1 298 1 0.40593361090161p
rp_12to1 12 1 42816.88333976
rc1_12to13 12 299 1e-05
cs1_12to13 299 13 9.7146778270048p
rp_12to13 12 13 1046.0253744493
rc1_12to14 12 300 1e-05
cs1_12to14 300 14 84.91713667402p
rp_12to14 12 14 83.221230108118
rc1_12to15 12 301 1e-05
cs1_12to15 301 15 390.85483901588p
rp_12to15 12 15 14.720739503755
rc1_12to16 12 302 1e-05
cs1_12to16 302 16 1927.7907804827p
rp_12to16 12 16 1.5906581273764
rc1_12to17 12 303 1e-05
cs1_12to17 303 17 339668.02413863p
rp_12to17 12 17 100000
rc1_12to18 12 304 1e-05
cs1_12to18 304 18 235.31520518942p
rp_12to18 12 18 28.796761181298
rc1_12to19 12 305 1e-05
cs1_12to19 305 19 38.4535062151p
rp_12to19 12 19 215.13084524273
rc1_12to20 12 306 1e-05
cs1_12to20 306 20 3.1031433448361p
rp_12to20 12 20 4109.2463607485
rc1_12to21 12 307 1e-05
cs1_12to21 307 21 1.6147956113083p
rp_12to21 12 21 8678.173535196
rc1_12to22 12 308 1e-05
cs1_12to22 308 22 24.597541128933p
rp_12to22 12 22 357.18612109718
rc1_12to23 12 309 1e-05
cs1_12to23 309 23 150.88784134738p
rp_12to23 12 23 45.154571809079
rc1_12to24 12 310 1e-05
cs1_12to24 310 24 622.26411098323p
rp_12to24 12 24 8.8987899615666
rc1_12to25 12 311 1e-05
cs1_12to25 311 25 3911.1575201822p
rp_12to25 12 25 0.48250531266968
rc1_12to26 12 312 1e-05
cs1_12to26 312 26 80.700563982526p
rp_12to26 12 26 92.537042491415
rc1_12to27 12 313 1e-05
cs1_12to27 313 27 9.4318993001427p
rp_12to27 12 27 1102.9994612529
rc1_12to28 12 314 1e-05
cs1_12to28 314 28 0.40154940339553p
rp_12to28 12 28 43849.832474915
rc1_12to29 12 315 1e-05
cs1_12to29 315 29 9.4444490760561p
rp_12to29 12 29 1100.463347048
rc1_12to30 12 316 1e-05
cs1_12to30 316 30 80.152562653249p
rp_12to30 12 30 92.492197401394
rc1_12to31 12 317 1e-05
cs1_12to31 317 31 357.79243601747p
rp_12to31 12 31 17.534239385876
rc1_12to32 12 318 1e-05
cs1_12to32 318 32 1601.6442149206p
rp_12to32 12 32 2.4163036689279
rc1_13to1 13 319 1e-05
cs1_13to1 319 1 0.40596030448156p
rp_13to1 13 1 42819.270556697
rc1_13to14 13 320 1e-05
cs1_13to14 320 14 9.7119539125129p
rp_13to14 13 14 1046.5684431132
rc1_13to15 13 321 1e-05
cs1_13to15 321 15 84.790570368422p
rp_13to15 13 15 83.507396790488
rc1_13to16 13 322 1e-05
cs1_13to16 322 16 387.35295412852p
rp_13to16 13 16 15.067403905632
rl1_13to17 13 323 -0.0019157788746038
ls1_13to17 323 17 -4.1288460601954e-05n
rc1_13to18 13 324 1e-05
cs1_13to18 324 18 946.84066062168p
rp_13to18 13 18 5.6990917624822
rc1_13to19 13 325 1e-05
cs1_13to19 325 19 205.49837714865p
rp_13to19 13 19 32.390991789611
rc1_13to20 13 326 1e-05
cs1_13to20 326 20 38.396928558854p
rp_13to20 13 20 215.09029160223
rc1_13to21 13 327 1e-05
cs1_13to21 327 21 3.1072592177309p
rp_13to21 13 21 4099.9543354474
rc1_13to22 13 328 1e-05
cs1_13to22 328 22 1.6142614294654p
rp_13to22 13 22 8682.3718684422
rc1_13to23 13 329 1e-05
cs1_13to23 329 23 24.583763049487p
rp_13to23 13 23 357.423328584
rc1_13to24 13 330 1e-05
cs1_13to24 330 24 150.66700837684p
rp_13to24 13 24 45.279936597947
rc1_13to25 13 331 1e-05
cs1_13to25 331 25 605.86494542509p
rp_13to25 13 25 9.4841775400526
rc1_13to26 13 332 1e-05
cs1_13to26 332 26 360.34342860089p
rp_13to26 13 26 17.622219767278
rc1_13to27 13 333 1e-05
cs1_13to27 333 27 80.054420664563p
rp_13to27 13 27 92.700553463004
rc1_13to28 13 334 1e-05
cs1_13to28 334 28 9.4444779718259p
rp_13to28 13 28 1100.457701788
rc1_13to29 13 335 1e-05
cs1_13to29 335 29 0.40157684446716p
rp_13to29 13 29 43852.550791082
rc1_13to30 13 336 1e-05
cs1_13to30 336 30 9.4418477578572p
rp_13to30 13 30 1101.04289794
rc1_13to31 13 337 1e-05
cs1_13to31 337 31 80.039180338628p
rp_13to31 13 31 92.798785637949
rc1_13to32 13 338 1e-05
cs1_13to32 338 32 354.77538575213p
rp_13to32 13 32 17.936115684071
rc1_14to1 14 339 1e-05
cs1_14to1 339 1 0.40592490236081p
rp_14to1 14 1 42817.176665294
rc1_14to15 14 340 1e-05
cs1_14to15 340 15 9.6951620186188p
rp_14to15 14 15 1049.1228050183
rc1_14to16 14 341 1e-05
cs1_14to16 341 16 84.417838851598p
rp_14to16 14 16 84.021815797529
rl1_14to17 14 342 -0.0015376011305242
ls1_14to17 342 17 -2.2123627673632e-05n
rc1_14to18 14 343 1e-05
cs1_14to18 343 18 7635.8182810117p
rp_14to18 14 18 0.14764147392388
rc1_14to19 14 344 1e-05
cs1_14to19 344 19 846.88809419401p
rp_14to19 14 19 5.9107902285661
rc1_14to20 14 345 1e-05
cs1_14to20 345 20 205.1607459868p
rp_14to20 14 20 32.506139934823
rc1_14to21 14 346 1e-05
cs1_14to21 346 21 38.438244410548p
rp_14to21 14 21 214.75675238359
rc1_14to22 14 347 1e-05
cs1_14to22 347 22 3.1085052850192p
rp_14to22 14 22 4098.3858668782
rc1_14to23 14 348 1e-05
cs1_14to23 348 23 1.6140992879236p
rp_14to23 14 23 8681.1654206662
rc1_14to24 14 349 1e-05
cs1_14to24 349 24 24.564039760145p
rp_14to24 14 24 357.87806223896
rc1_14to25 14 350 1e-05
cs1_14to25 350 25 147.90478081113p
rp_14to25 14 25 46.4344325209
rc1_14to26 14 351 1e-05
cs1_14to26 351 26 1616.1831587718p
rp_14to26 14 26 2.4238052103942
rc1_14to27 14 352 1e-05
cs1_14to27 352 27 357.96138566719p
rp_14to27 14 27 17.506153732872
rc1_14to28 14 353 1e-05
cs1_14to28 353 28 80.155372343449p
rp_14to28 14 28 92.476720897356
rc1_14to29 14 354 1e-05
cs1_14to29 354 29 9.4418681807587p
rp_14to29 14 29 1101.0230593759
rc1_14to30 14 355 1e-05
cs1_14to30 355 30 0.40154025402077p
rp_14to30 14 30 43852.016211628
rc1_14to31 14 356 1e-05
cs1_14to31 356 31 9.4257808544023p
rp_14to31 14 31 1103.5769097689
rc1_14to32 14 357 1e-05
cs1_14to32 357 32 79.690211019667p
rp_14to32 14 32 93.333514996139
rc1_15to1 15 358 1e-05
cs1_15to1 358 1 0.40611709010247p
rp_15to1 15 1 42778.231243437
rc1_15to16 15 359 1e-05
cs1_15to16 359 16 9.7046430253688p
rp_15to16 15 16 1046.977474235
rl1_15to17 15 360 -0.0015962388438325
ls1_15to17 360 17 -0.00029631991092396n
rc1_15to18 15 361 1e-05
cs1_15to18 361 18 6450.2640933358p
rp_15to18 15 18 0.010457909252505
rc1_15to19 15 362 1e-05
cs1_15to19 362 19 1923.5373528311p
rp_15to19 15 19 0.033814488562545
rc1_15to20 15 363 1e-05
cs1_15to20 363 20 845.62500499493p
rp_15to20 15 20 5.8992910529199
rc1_15to21 15 364 1e-05
cs1_15to21 364 21 205.03384981556p
rp_15to21 15 21 32.409074881686
rc1_15to22 15 365 1e-05
cs1_15to22 365 22 38.407634344382p
rp_15to22 15 22 215.16838442024
rc1_15to23 15 366 1e-05
cs1_15to23 366 23 3.1013640471335p
rp_15to23 15 23 4112.4349342132
rc1_15to24 15 367 1e-05
cs1_15to24 367 24 1.6169540000411p
rp_15to24 15 24 8662.7036514111
rc1_15to25 15 368 1e-05
cs1_15to25 368 25 24.310725072133p
rp_15to25 15 25 361.37159584574
rc1_15to26 15 369 1e-05
cs1_15to26 369 26 2935.5864667831p
rp_15to26 15 26 0.022680491541016
rc1_15to27 15 370 1e-05
cs1_15to27 370 27 1624.7087887794p
rp_15to27 15 27 2.3488467433714
rc1_15to28 15 371 1e-05
cs1_15to28 371 28 357.80271289486p
rp_15to28 15 28 17.534854200563
rc1_15to29 15 372 1e-05
cs1_15to29 372 29 80.03827701963p
rp_15to29 15 29 92.799569527043
rc1_15to30 15 373 1e-05
cs1_15to30 373 30 9.4257545739553p
rp_15to30 15 30 1103.6054582704
rc1_15to31 15 374 1e-05
cs1_15to31 374 31 0.40172903228212p
rp_15to31 15 31 43809.894960861
rc1_15to32 15 375 1e-05
cs1_15to32 375 32 9.4341473905223p
rp_15to32 15 32 1101.4910677676
rc1_16to1 16 376 1e-05
cs1_16to1 376 1 0.40563866637065p
rp_16to1 16 1 42837.890626691
rl1_16to17 16 377 -0.00053796298241023
ls1_16to17 377 17 -0.00021119767950794n
rl1_16to18 16 378 0.0020043498887601
ls1_16to18 378 18 0.0055761848797159n
rl1_16to19 16 379 0.00470007444172
ls1_16to19 379 19 0.00081858479228345n
rc1_16to20 16 380 1e-05
cs1_16to20 380 20 1905.3449670611p
rp_16to20 16 20 0.034247194659992
rc1_16to21 16 381 1e-05
cs1_16to21 381 21 836.26881369959p
rp_16to21 16 21 6.0150585845314
rc1_16to22 16 382 1e-05
cs1_16to22 382 22 203.90692624029p
rp_16to22 16 22 32.025833166338
rc1_16to23 16 383 1e-05
cs1_16to23 383 23 38.255544958162p
rp_16to23 16 23 215.8621252811
rc1_16to24 16 384 1e-05
cs1_16to24 384 24 3.1017215455118p
rp_16to24 16 24 4107.9281976881
rc1_16to25 16 385 1e-05
cs1_16to25 385 25 1.6041656742642p
rp_16to25 16 25 8713.0534000004
rl1_16to26 16 386 0.0035323269327029
ls1_16to26 386 26 0.0043289727902135n
rc1_16to27 16 387 1e-05
cs1_16to27 387 27 2877.6540350893p
rp_16to27 16 27 0.023178898088768
rc1_16to28 16 388 1e-05
cs1_16to28 388 28 1602.5066478999p
rp_16to28 16 28 2.4123470094235
rc1_16to29 16 389 1e-05
cs1_16to29 389 29 354.78481853476p
rp_16to29 16 29 17.92998372001
rc1_16to30 16 390 1e-05
cs1_16to30 390 30 79.68971685294p
rp_16to30 16 30 93.336982339848
rc1_16to31 16 391 1e-05
cs1_16to31 391 31 9.4341687854027p
rp_16to31 16 31 1101.4865168827
rc1_16to32 16 392 1e-05
cs1_16to32 392 32 0.40125218508848p
rp_16to32 16 32 43871.706163175
rl1_17to1 17 393 4069.5196953433
ls1_17to1 393 1 234.46944364689n
rs2_17to1 17 394 0.045024888478556
ls2_17to1 394 1 2.1262758616504n
rl1_17to18 17 395 0.010902906193865
ls1_17to18 395 18 0.64512361477305n
rl1_17to19 17 396 0.00059154914502269
ls1_17to19 396 19 0.080482571253722n
rl1_17to20 17 397 -29.465530221036
ls1_17to20 397 20 -4.2722513768733n
rs2_17to20 17 398 0.000307588357465
ls2_17to20 398 20 0.020980359053249n
rl1_17to21 17 399 0.0002679739381116
ls1_17to21 399 21 0.0072244368508427n
rl1_17to22 17 400 0.00015294413746195
ls1_17to22 400 22 0.0028148792604339n
rl1_17to23 17 401 8.8136680126018e-05
ls1_17to23 401 23 0.0011520912324482n
rl1_17to24 17 402 5.2520660824885e-05
ls1_17to24 402 24 0.00045344656055357n
rl1_17to25 17 403 3.1086546130782e-05
ls1_17to25 403 25 0.0001570727763413n
rl1_17to26 17 404 0.0018602140372799
ls1_17to26 404 26 0.16167464768478n
rl1_17to27 17 405 10.426550229406
ls1_17to27 405 27 5.1639584439222n
rs2_17to27 17 406 0.00031079307925277
ls2_17to27 406 27 0.033686206246325n
rl1_17to28 17 407 0.00027607092320056
ls1_17to28 407 28 0.010724038799013n
rl1_17to29 17 408 0.00019291388607519
ls1_17to29 408 29 0.0040419667392133n
rl1_17to30 17 409 0.00011801347262176
ls1_17to30 409 30 0.0016343874582087n
rl1_17to31 17 410 6.7635822381382e-05
ls1_17to31 410 31 0.00065398039718159n
rl1_17to32 17 411 3.9686571015755e-05
ls1_17to32 411 32 0.00024949696706294n
rc1_18to1 18 412 1e-05
cs1_18to1 412 1 0.43298616961017p
rp_18to1 18 1 41491.488920972
rc1_18to19 18 413 1e-05
cs1_18to19 413 19 10.772703044598p
rp_18to19 18 19 974.91443599522
rc1_18to20 18 414 1e-05
cs1_18to20 414 20 98.701675890599p
rp_18to20 18 20 73.103128075548
rc1_18to21 18 415 1e-05
cs1_18to21 415 21 465.84580630041p
rp_18to21 18 21 12.521374837882
rc1_18to22 18 416 1e-05
cs1_18to22 416 22 2297.198909076p
rp_18to22 18 22 1.3375598739112
rc1_18to23 18 417 1e-05
cs1_18to23 417 23 3457.9624206628p
rp_18to23 18 23 0.018875996177116
rl1_18to24 18 418 0.0030093279271015
ls1_18to24 418 24 0.0037025455955647n
rl1_18to25 18 419 0.0015944124650371
ls1_18to25 419 25 0.0068854301459153n
rc1_18to26 18 420 1e-05
cs1_18to26 420 26 3.45031361314p
rp_18to26 18 26 3765.8396742715
rc1_18to27 18 421 1e-05
cs1_18to27 421 27 45.929104391786p
rp_18to27 18 27 177.16571702539
rc1_18to28 18 422 1e-05
cs1_18to28 422 28 261.9445609924p
rp_18to28 18 28 23.458514065156
rc1_18to29 18 423 1e-05
cs1_18to29 423 29 1138.5155061859p
rp_18to29 18 29 3.8494809313927
rc1_18to30 18 424 1e-05
cs1_18to30 424 30 2290.4260504326p
rp_18to30 18 30 0.027947122379457
rl1_18to31 18 425 0.003923412106832
ls1_18to31 425 31 0.00079664187600247n
rl1_18to32 18 426 0.0020889530043902
ls1_18to32 426 32 0.0061182835736309n
rc1_19to1 19 427 1e-05
cs1_19to1 427 1 0.40627723351314p
rp_19to1 19 1 42786.053763237
rc1_19to20 19 428 1e-05
cs1_19to20 428 20 9.720345549135p
rp_19to20 19 20 1046.361759538
rc1_19to21 19 429 1e-05
cs1_19to21 429 21 85.172332566295p
rp_19to21 19 21 82.867614552953
rc1_19to22 19 430 1e-05
cs1_19to22 430 22 394.7080106099p
rp_19to22 19 22 14.400731936724
rc1_19to23 19 431 1e-05
cs1_19to23 431 23 2024.3723243656p
rp_19to23 19 23 1.4084632572182
rc1_19to24 19 432 1e-05
cs1_19to24 432 24 2908.5643487458p
rp_19to24 19 24 0.022932112209635
rl1_19to25 19 433 0.0036976849655179
ls1_19to25 433 25 0.005178288951651n
rc1_19to26 19 434 1e-05
cs1_19to26 434 26 1.6470307441643p
rp_19to26 19 26 8422.8201658281
rc1_19to27 19 435 1e-05
cs1_19to27 435 27 3.1673416375692p
rp_19to27 19 27 3959.5503942303
rc1_19to28 19 436 1e-05
cs1_19to28 436 28 40.295058985114p
rp_19to28 19 28 197.1742090784
rc1_19to29 19 437 1e-05
cs1_19to29 437 29 222.54369580354p
rp_19to29 19 29 27.672833051519
rc1_19to30 19 438 1e-05
cs1_19to30 438 30 974.67949271402p
rp_19to30 19 30 4.3642634847173
rc1_19to31 19 439 1e-05
cs1_19to31 439 31 1926.9533015115p
rp_19to31 19 31 0.033950358973915
rl1_19to32 19 440 0.0048072192233508
ls1_19to32 440 32 0.0017946222277593n
rc1_20to1 20 441 1e-05
cs1_20to1 441 1 0.40574437658665p
rp_20to1 20 1 42856.846043001
rc1_20to21 20 442 1e-05
cs1_20to21 442 21 9.7022827227051p
rp_20to21 20 21 1047.7037525656
rc1_20to22 20 443 1e-05
cs1_20to22 443 22 84.99368606703p
rp_20to22 20 22 82.849423685231
rc1_20to23 20 444 1e-05
cs1_20to23 444 23 393.9341324034p
rp_20to23 20 23 14.369811842738
rc1_20to24 20 445 1e-05
cs1_20to24 445 24 2026.4848521994p
rp_20to24 20 24 1.3918247248737
rc1_20to25 20 446 1e-05
cs1_20to25 446 25 2843.6327957763p
rp_20to25 20 25 0.023439001141783
rc1_20to26 20 447 1e-05
cs1_20to26 447 26 25.775617009965p
rp_20to26 20 26 331.59603542355
rc1_20to27 20 448 1e-05
cs1_20to27 448 27 1.6402389391099p
rp_20to27 20 27 8437.9751831806
rc1_20to28 20 449 1e-05
cs1_20to28 449 28 3.163007660765p
rp_20to28 20 28 3962.2691439446
rc1_20to29 20 450 1e-05
cs1_20to29 450 29 40.227949041049p
rp_20to29 20 29 197.16405397547
rc1_20to30 20 451 1e-05
cs1_20to30 451 30 222.12021832437p
rp_20to30 20 30 27.804138286745
rc1_20to31 20 452 1e-05
cs1_20to31 452 31 973.59056953418p
rp_20to31 20 31 4.3426649186041
rc1_20to32 20 453 1e-05
cs1_20to32 453 32 1908.6407554896p
rp_20to32 20 32 0.034301813124795
rc1_21to1 21 454 1e-05
cs1_21to1 454 1 0.40583755590414p
rp_21to1 21 1 42833.576765623
rc1_21to22 21 455 1e-05
cs1_21to22 455 22 9.714415242436p
rp_21to22 21 22 1045.4893272849
rc1_21to23 21 456 1e-05
cs1_21to23 456 23 85.022190742332p
rp_21to23 21 23 82.845411602183
rc1_21to24 21 457 1e-05
cs1_21to24 457 24 393.18358276695p
rp_21to24 21 24 14.471141266411
rc1_21to25 21 458 1e-05
cs1_21to25 458 25 1928.3892634494p
rp_21to25 21 25 1.5381729208358
rc1_21to26 21 459 1e-05
cs1_21to26 459 26 163.95240845262p
rp_21to26 21 26 39.154704977015
rc1_21to27 21 460 1e-05
cs1_21to27 460 27 25.584483000632p
rp_21to27 21 27 332.75724821681
rc1_21to28 21 461 1e-05
cs1_21to28 461 28 1.6406425807123p
rp_21to28 21 28 8434.4449339482
rc1_21to29 21 462 1e-05
cs1_21to29 462 29 3.1672576394348p
rp_21to29 21 29 3953.6188774808
rc1_21to30 21 463 1e-05
cs1_21to30 463 30 40.27198858387p
rp_21to30 21 30 196.82415799154
rc1_21to31 21 464 1e-05
cs1_21to31 464 31 221.95622220934p
rp_21to31 21 31 27.683076585254
rc1_21to32 21 465 1e-05
cs1_21to32 465 32 961.18749264044p
rp_21to32 21 32 4.4513821309469
rc1_22to1 22 466 1e-05
cs1_22to1 466 1 0.40601177759407p
rp_22to1 22 1 42801.180056543
rc1_22to23 22 467 1e-05
cs1_22to23 467 23 9.7154884058189p
rp_22to23 22 23 1045.5649157072
rc1_22to24 22 468 1e-05
cs1_22to24 468 24 84.985730181275p
rp_22to24 22 24 83.002546641782
rc1_22to25 22 469 1e-05
cs1_22to25 469 25 384.70524647243p
rp_22to25 22 25 14.946754438802
rc1_22to26 22 470 1e-05
cs1_22to26 470 26 709.00730575701p
rp_22to26 22 26 6.8849625162435
rc1_22to27 22 471 1e-05
cs1_22to27 471 27 162.27796449355p
rp_22to27 22 27 39.362995029
rc1_22to28 22 472 1e-05
cs1_22to28 472 28 25.6154056625p
rp_22to28 22 28 332.15334667908
rc1_22to29 22 473 1e-05
cs1_22to29 473 29 1.6401012316401p
rp_22to29 22 29 8438.2766059586
rc1_22to30 22 474 1e-05
cs1_22to30 474 30 3.1685346726089p
rp_22to30 22 30 3952.1078850743
rc1_22to31 22 475 1e-05
cs1_22to31 475 31 40.238276416453p
rp_22to31 22 31 197.24288425028
rc1_22to32 22 476 1e-05
cs1_22to32 476 32 220.67641656785p
rp_22to32 22 32 27.50709152786
rc1_23to1 23 477 1e-05
cs1_23to1 477 1 0.40584432438078p
rp_23to1 23 1 42849.503236943
rc1_23to24 23 478 1e-05
cs1_23to24 478 24 9.7043773717418p
rp_23to24 23 24 1047.2900714811
rc1_23to25 23 479 1e-05
cs1_23to25 479 25 83.53545364612p
rp_23to25 23 25 84.604147508999
rc1_23to26 23 480 1e-05
cs1_23to26 480 26 5749.6253429538p
rp_23to26 23 26 0.080552547482226
rc1_23to27 23 481 1e-05
cs1_23to27 481 27 703.87926076626p
rp_23to27 23 27 6.8459737966681
rc1_23to28 23 482 1e-05
cs1_23to28 482 28 162.35039350367p
rp_23to28 23 28 39.330321663809
rc1_23to29 23 483 1e-05
cs1_23to29 483 29 25.600572044361p
rp_23to29 23 29 332.41842421687
rc1_23to30 23 484 1e-05
cs1_23to30 484 30 1.6399294576581p
rp_23to30 23 30 8437.7128793376
rc1_23to31 23 485 1e-05
cs1_23to31 485 31 3.1611768950567p
rp_23to31 23 31 3965.4691965646
rc1_23to32 23 486 1e-05
cs1_23to32 486 32 40.080031082405p
rp_23to32 23 32 197.91476882081
rc1_24to1 24 487 1e-05
cs1_24to1 487 1 0.40561749459376p
rp_24to1 24 1 42859.643144341
rc1_24to25 24 488 1e-05
cs1_24to25 488 25 9.6183084803188p
rp_24to25 24 25 1054.7304198344
rc1_24to26 24 489 1e-05
cs1_24to26 489 26 4434.8194278094p
rp_24to26 24 26 0.015366170038386
rc1_24to27 24 490 1e-05
cs1_24to27 490 27 1543.4346161513p
rp_24to27 24 27 0.042308679857434
rc1_24to28 24 491 1e-05
cs1_24to28 491 28 702.61676020236p
rp_24to28 24 28 6.8837366125805
rc1_24to29 24 492 1e-05
cs1_24to29 492 29 162.09502007432p
rp_24to29 24 29 39.451039441062
rc1_24to30 24 493 1e-05
cs1_24to30 493 30 25.579908935857p
rp_24to30 24 30 332.83194308333
rc1_24to31 24 494 1e-05
cs1_24to31 494 31 1.6428697019955p
rp_24to31 24 31 8418.6122282375
rc1_24to32 24 495 1e-05
cs1_24to32 495 32 3.1616960678635p
rp_24to32 24 32 3961.4261437739
rc1_25to1 25 496 1e-05
cs1_25to1 496 1 0.40382701505571p
rp_25to1 25 1 42941.656563542
rl1_25to26 25 497 0.0027405021527526
ls1_25to26 497 26 0.0071413866864488n
rc1_25to27 25 498 1e-05
cs1_25to27 498 27 4290.3753370065p
rp_25to27 25 27 0.015936054287024
rc1_25to28 25 499 1e-05
cs1_25to28 499 28 5702.7187306267p
rp_25to28 25 28 0.090531720800414
rc1_25to29 25 500 1e-05
cs1_25to29 500 29 682.66265130296p
rp_25to29 25 29 7.3329589187613
rc1_25to30 25 501 1e-05
cs1_25to30 501 30 159.07744476134p
rp_25to30 25 30 40.487365619484
rc1_25to31 25 502 1e-05
cs1_25to31 502 31 25.3199644328p
rp_25to31 25 31 336.09818151614
rc1_25to32 25 503 1e-05
cs1_25to32 503 32 1.6300037566837p
rp_25to32 25 32 8468.2947192628
rc1_26to1 26 504 1e-05
cs1_26to1 504 1 0.40641199337029p
rp_26to1 26 1 42889.687594037
rc1_26to27 26 505 1e-05
cs1_26to27 505 27 9.7604981798369p
rp_26to27 26 27 1044.9918318926
rc1_26to28 26 506 1e-05
cs1_26to28 506 28 85.793745439329p
rp_26to28 26 28 82.550655439247
rc1_26to29 26 507 1e-05
cs1_26to29 507 29 397.65433681609p
rp_26to29 26 29 14.393872957867
rc1_26to30 26 508 1e-05
cs1_26to30 508 30 2021.6422777511p
rp_26to30 26 30 1.4323877955469
rc1_26to31 26 509 1e-05
cs1_26to31 509 31 2941.5672697043p
rp_26to31 26 31 0.022622945099888
rl1_26to32 26 510 0.0036137883603056
ls1_26to32 510 32 0.0050851925181991n
rc1_27to1 27 511 1e-05
cs1_27to1 511 1 0.40577345456889p
rp_27to1 27 1 42860.710301192
rc1_27to28 27 512 1e-05
cs1_27to28 512 28 9.7044142956059p
rp_27to28 27 28 1047.3655060332
rc1_27to29 27 513 1e-05
cs1_27to29 513 29 84.991520451766p
rp_27to29 27 29 82.884458644134
rc1_27to30 27 514 1e-05
cs1_27to30 514 30 394.19928893047p
rp_27to30 27 30 14.338884813469
rc1_27to31 27 515 1e-05
cs1_27to31 515 31 2031.1314766688p
rp_27to31 27 31 1.3843849942608
rc1_27to32 27 516 1e-05
cs1_27to32 516 32 2883.2678873169p
rp_27to32 27 32 0.023139639541654
rc1_28to1 28 517 1e-05
cs1_28to1 517 1 0.40593970621883p
rp_28to1 28 1 42814.681134363
rc1_28to29 28 518 1e-05
cs1_28to29 518 29 9.7173540330142p
rp_28to29 28 29 1045.0424188131
rc1_28to30 28 519 1e-05
cs1_28to30 519 30 85.09612908955p
rp_28to30 28 30 82.697931710588
rc1_28to31 28 520 1e-05
cs1_28to31 520 31 393.9114969778p
rp_28to31 28 31 14.383725875485
rc1_28to32 28 521 1e-05
cs1_28to32 521 32 1994.5859811683p
rp_28to32 28 32 1.4415927311594
rc1_29to1 29 522 1e-05
cs1_29to1 522 1 0.40596684747184p
rp_29to1 29 1 42817.339892573
rc1_29to30 29 523 1e-05
cs1_29to30 523 30 9.7146548903963p
rp_29to30 29 30 1045.5779984786
rc1_29to31 29 524 1e-05
cs1_29to31 524 31 84.968077870741p
rp_29to31 29 31 82.9954849553
rc1_29to32 29 525 1e-05
cs1_29to32 525 32 390.4465296422p
rp_29to32 29 32 14.695696616178
rc1_30to1 30 526 1e-05
cs1_30to1 526 1 0.40593119183859p
rp_30to1 30 1 42815.037442806
rc1_30to31 30 527 1e-05
cs1_30to31 527 31 9.6978215832833p
rp_30to31 30 31 1048.1257934703
rc1_30to32 30 528 1e-05
cs1_30to32 528 32 84.597699361319p
rp_30to32 30 32 83.4832478845
rc1_31to1 31 529 1e-05
cs1_31to1 529 1 0.40612358448068p
rp_31to1 31 1 42776.508660012
rc1_31to32 31 530 1e-05
cs1_31to32 530 32 9.7073846050711p
rp_31to32 31 32 1045.9834142785
rc1_32to1 32 531 1e-05
cs1_32to1 531 1 0.40564496675129p
rp_32to1 32 1 42835.838103073
rc1_1to0 1 532 1e-05
cs1_1to0 532 0 0.15828045803983p
rp_1to0 1 0 103163.59176811
rc1_2to0 2 533 1e-05
cs1_2to0 533 0 0.13711365766277p
rp_2to0 2 0 110587.50142019
rc1_3to0 3 534 1e-05
cs1_3to0 534 0 0.1351691049655p
rp_3to0 3 0 111514.60521895
rc1_4to0 4 535 1e-05
cs1_4to0 535 0 0.13454022112813p
rp_4to0 4 0 111191.86506292
rc1_5to0 5 536 1e-05
cs1_5to0 536 0 0.13449856329044p
rp_5to0 5 0 110478.85971134
rc1_6to0 6 537 1e-05
cs1_6to0 537 0 0.13460860187787p
rp_6to0 6 0 116435.06310034
rc1_7to0 7 538 1e-05
cs1_7to0 538 0 0.13466315806189p
rp_7to0 7 0 110880.46960973
rc1_8to0 8 539 1e-05
cs1_8to0 539 0 0.13537892665714p
rp_8to0 8 0 113054.6210311
rc1_9to0 9 540 1e-05
cs1_9to0 540 0 0.15818911632458p
rp_9to0 9 0 103899.14607306
rc1_10to0 10 541 1e-05
cs1_10to0 541 0 0.13535046246074p
rp_10to0 10 0 113438.10763738
rc1_11to0 11 542 1e-05
cs1_11to0 542 0 0.13466426202679p
rp_11to0 11 0 111539.84924008
rc1_12to0 12 543 1e-05
cs1_12to0 543 0 0.1346058899936p
rp_12to0 12 0 112230.98080211
rc1_13to0 13 544 1e-05
cs1_13to0 544 0 0.13457832857187p
rp_13to0 13 0 109661.66660797
rc1_14to0 14 545 1e-05
cs1_14to0 545 0 0.13462750898413p
rp_14to0 14 0 111798.40059284
rc1_15to0 15 546 1e-05
cs1_15to0 546 0 0.13512212113875p
rp_15to0 15 0 110382.75704512
rc1_16to0 16 547 1e-05
cs1_16to0 547 0 0.13718366364731p
rp_16to0 16 0 111554.57055898
rc1_17to0 17 548 1e-05
cs1_17to0 548 0 0.15735245320767p
rp_17to0 17 0 102621.03549512
rc1_18to0 18 549 1e-05
cs1_18to0 549 0 0.13632625172402p
rp_18to0 18 0 115661.47270854
rc1_19to0 19 550 1e-05
cs1_19to0 550 0 0.13422659347244p
rp_19to0 19 0 114514.16924424
rc1_20to0 20 551 1e-05
cs1_20to0 551 0 0.13361185371055p
rp_20to0 20 0 115385.56069783
rc1_21to0 21 552 1e-05
cs1_21to0 552 0 0.13357409345759p
rp_21to0 21 0 116027.81736224
rc1_22to0 22 553 1e-05
cs1_22to0 553 0 0.13364769225729p
rp_22to0 22 0 109915.57995897
rc1_23to0 23 554 1e-05
cs1_23to0 554 0 0.13373273500924p
rp_23to0 23 0 115813.34636057
rc1_24to0 24 555 1e-05
cs1_24to0 555 0 0.13456981787534p
rp_24to0 24 0 113573.1532417
rc1_25to0 25 556 1e-05
cs1_25to0 556 0 0.15719934371391p
rp_25to0 25 0 102182.75257135
rc1_26to0 26 557 1e-05
cs1_26to0 557 0 0.13454326011948p
rp_26to0 26 0 113269.52864015
rc1_27to0 27 558 1e-05
cs1_27to0 558 0 0.13375816833412p
rp_27to0 27 0 115051.05790188
rc1_28to0 28 559 1e-05
cs1_28to0 559 0 0.1335864557518p
rp_28to0 28 0 114021.40058994
rc1_29to0 29 560 1e-05
cs1_29to0 560 0 0.13356634739669p
rp_29to0 29 0 116871.72877678
rc1_30to0 30 561 1e-05
cs1_30to0 561 0 0.13370630968212p
rp_30to0 30 0 114459.73750749
rc1_31to0 31 562 1e-05
cs1_31to0 562 0 0.13421266863567p
rp_31to0 31 0 115804.98407774
rc1_32to0 32 563 1e-05
cs1_32to0 563 0 0.1364335128246p
rp_32to0 32 0 114423.3610862
.ends m16lines_HFSS_lfws

