* BEGIN ANSOFT HEADER
* node 1    trace_p_0_T1
* node 2    trace_n_0_T1
* node 3    trace_p_1_T1
* node 4    trace_n_1_T1
* node 5    trace_p_2_T1
* node 6    trace_n_2_T1
* node 7    trace_p_3_T1
* node 8    trace_n_3_T1
* node 9    trace_p_4_T1
* node 10   trace_n_4_T1
* node 11   trace_p_5_T1
* node 12   trace_n_5_T1
* node 13   trace_p_6_T1
* node 14   trace_n_6_T1
* node 15   trace_p_7_T1
* node 16   trace_n_7_T1
* node 17   trace_p_0_T2
* node 18   trace_n_0_T2
* node 19   trace_p_1_T2
* node 20   trace_n_1_T2
* node 21   trace_p_2_T2
* node 22   trace_n_2_T2
* node 23   trace_p_3_T2
* node 24   trace_n_3_T2
* node 25   trace_p_4_T2
* node 26   trace_n_4_T2
* node 27   trace_p_5_T2
* node 28   trace_n_5_T2
* node 29   trace_p_6_T2
* node 30   trace_n_6_T2
* node 31   trace_p_7_T2
* node 32   trace_n_7_T2
*   Format: HSPICE
*   Topckt: m16lines_port_fws
*     Date: Sat Jun 06 11:16:33 2020
*    Notes: Frequency range: 1e+08 to 7e+10 Hz, 700 points
*         : Maximum number of poles: 10000
*         : S-Matrix fitting error tolerance: 0.001
*         : Causality check tolerance: auto
*         : Passivity enforcement: on (by iterated fitting)
*         : Causality enforcement: off
*         : Fitting method: FastFit
*         : Matrix fitting: By entire matrix (required by FastFit)
*         : Ensure Z-parameter accuracy: on
*         : Relative error control: off
*         : Common ground option: on
*         : Final fitting error: 0.0148652
*         : Final model order: 256
* END ANSOFT HEADER

.subckt m16lines_port_fws 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21
+ 22 23 24 25 26 27 28 29 30 31 32
Vam1 1 n2 dc 0
Rport1 n2 0 50 noise=0
Vam2 2 n4 dc 0
Rport2 n4 0 50 noise=0
Vam3 3 n6 dc 0
Rport3 n6 0 50 noise=0
Vam4 4 n8 dc 0
Rport4 n8 0 50 noise=0
Vam5 5 n10 dc 0
Rport5 n10 0 50 noise=0
Vam6 6 n12 dc 0
Rport6 n12 0 50 noise=0
Vam7 7 n14 dc 0
Rport7 n14 0 50 noise=0
Vam8 8 n16 dc 0
Rport8 n16 0 50 noise=0
Vam9 9 n18 dc 0
Rport9 n18 0 50 noise=0
Vam10 10 n20 dc 0
Rport10 n20 0 50 noise=0
Vam11 11 n22 dc 0
Rport11 n22 0 50 noise=0
Vam12 12 n24 dc 0
Rport12 n24 0 50 noise=0
Vam13 13 n26 dc 0
Rport13 n26 0 50 noise=0
Vam14 14 n28 dc 0
Rport14 n28 0 50 noise=0
Vam15 15 n30 dc 0
Rport15 n30 0 50 noise=0
Vam16 16 n32 dc 0
Rport16 n32 0 50 noise=0
Vam17 17 n34 dc 0
Rport17 n34 0 50 noise=0
Vam18 18 n36 dc 0
Rport18 n36 0 50 noise=0
Vam19 19 n38 dc 0
Rport19 n38 0 50 noise=0
Vam20 20 n40 dc 0
Rport20 n40 0 50 noise=0
Vam21 21 n42 dc 0
Rport21 n42 0 50 noise=0
Vam22 22 n44 dc 0
Rport22 n44 0 50 noise=0
Vam23 23 n46 dc 0
Rport23 n46 0 50 noise=0
Vam24 24 n48 dc 0
Rport24 n48 0 50 noise=0
Vam25 25 n50 dc 0
Rport25 n50 0 50 noise=0
Vam26 26 n52 dc 0
Rport26 n52 0 50 noise=0
Vam27 27 n54 dc 0
Rport27 n54 0 50 noise=0
Vam28 28 n56 dc 0
Rport28 n56 0 50 noise=0
Vam29 29 n58 dc 0
Rport29 n58 0 50 noise=0
Vam30 30 n60 dc 0
Rport30 n60 0 50 noise=0
Vam31 31 n62 dc 0
Rport31 n62 0 50 noise=0
Vam32 32 n64 dc 0
Rport32 n64 0 50 noise=0

Fi1 0 ni1 Vam1 50
Gi1 0 ni1 1 0 1
Rt1 ni1 0 1 noise=0
Fi2 0 ni2 Vam2 50
Gi2 0 ni2 2 0 1
Rt2 ni2 0 1 noise=0
Fi3 0 ni3 Vam3 50
Gi3 0 ni3 3 0 1
Rt3 ni3 0 1 noise=0
Fi4 0 ni4 Vam4 50
Gi4 0 ni4 4 0 1
Rt4 ni4 0 1 noise=0
Fi5 0 ni5 Vam5 50
Gi5 0 ni5 5 0 1
Rt5 ni5 0 1 noise=0
Fi6 0 ni6 Vam6 50
Gi6 0 ni6 6 0 1
Rt6 ni6 0 1 noise=0
Fi7 0 ni7 Vam7 50
Gi7 0 ni7 7 0 1
Rt7 ni7 0 1 noise=0
Fi8 0 ni8 Vam8 50
Gi8 0 ni8 8 0 1
Rt8 ni8 0 1 noise=0
Fi9 0 ni9 Vam9 50
Gi9 0 ni9 9 0 1
Rt9 ni9 0 1 noise=0
Fi10 0 ni10 Vam10 50
Gi10 0 ni10 10 0 1
Rt10 ni10 0 1 noise=0
Fi11 0 ni11 Vam11 50
Gi11 0 ni11 11 0 1
Rt11 ni11 0 1 noise=0
Fi12 0 ni12 Vam12 50
Gi12 0 ni12 12 0 1
Rt12 ni12 0 1 noise=0
Fi13 0 ni13 Vam13 50
Gi13 0 ni13 13 0 1
Rt13 ni13 0 1 noise=0
Fi14 0 ni14 Vam14 50
Gi14 0 ni14 14 0 1
Rt14 ni14 0 1 noise=0
Fi15 0 ni15 Vam15 50
Gi15 0 ni15 15 0 1
Rt15 ni15 0 1 noise=0
Fi16 0 ni16 Vam16 50
Gi16 0 ni16 16 0 1
Rt16 ni16 0 1 noise=0
Fi17 0 ni17 Vam17 50
Gi17 0 ni17 17 0 1
Rt17 ni17 0 1 noise=0
Fi18 0 ni18 Vam18 50
Gi18 0 ni18 18 0 1
Rt18 ni18 0 1 noise=0
Fi19 0 ni19 Vam19 50
Gi19 0 ni19 19 0 1
Rt19 ni19 0 1 noise=0
Fi20 0 ni20 Vam20 50
Gi20 0 ni20 20 0 1
Rt20 ni20 0 1 noise=0
Fi21 0 ni21 Vam21 50
Gi21 0 ni21 21 0 1
Rt21 ni21 0 1 noise=0
Fi22 0 ni22 Vam22 50
Gi22 0 ni22 22 0 1
Rt22 ni22 0 1 noise=0
Fi23 0 ni23 Vam23 50
Gi23 0 ni23 23 0 1
Rt23 ni23 0 1 noise=0
Fi24 0 ni24 Vam24 50
Gi24 0 ni24 24 0 1
Rt24 ni24 0 1 noise=0
Fi25 0 ni25 Vam25 50
Gi25 0 ni25 25 0 1
Rt25 ni25 0 1 noise=0
Fi26 0 ni26 Vam26 50
Gi26 0 ni26 26 0 1
Rt26 ni26 0 1 noise=0
Fi27 0 ni27 Vam27 50
Gi27 0 ni27 27 0 1
Rt27 ni27 0 1 noise=0
Fi28 0 ni28 Vam28 50
Gi28 0 ni28 28 0 1
Rt28 ni28 0 1 noise=0
Fi29 0 ni29 Vam29 50
Gi29 0 ni29 29 0 1
Rt29 ni29 0 1 noise=0
Fi30 0 ni30 Vam30 50
Gi30 0 ni30 30 0 1
Rt30 ni30 0 1 noise=0
Fi31 0 ni31 Vam31 50
Gi31 0 ni31 31 0 1
Rt31 ni31 0 1 noise=0
Fi32 0 ni32 Vam32 50
Gi32 0 ni32 32 0 1
Rt32 ni32 0 1 noise=0

Ca1 ns1 0 1e-12
Ra1 ns1 0 0.246835352493 noise=0
Ca2 ns2 0 1e-12
Ca3 ns3 0 1e-12
Ra2 ns2 0 5.85392236353 noise=0
Ra3 ns3 0 5.85392236353 noise=0
Ga2 ns2 0 ns3 0 -1.24965224039
Ga3 ns3 0 ns2 0 1.24965224039
Ca4 ns4 0 1e-12
Ca5 ns5 0 1e-12
Ra4 ns4 0 3.75353660859 noise=0
Ra5 ns5 0 3.75353660859 noise=0
Ga4 ns4 0 ns5 0 -0.431489095244
Ga5 ns5 0 ns4 0 0.431489095244
Ca6 ns6 0 1e-12
Ra6 ns6 0 12.1731904857 noise=0
Ca7 ns7 0 1e-12
Ra7 ns7 0 531.342615159 noise=0
Ca8 ns8 0 1e-12
Ra8 ns8 0 4008.18525934 noise=0
Ca9 ns9 0 1e-12
Ra9 ns9 0 0.246835352493 noise=0
Ca10 ns10 0 1e-12
Ca11 ns11 0 1e-12
Ra10 ns10 0 5.85392236353 noise=0
Ra11 ns11 0 5.85392236353 noise=0
Ga10 ns10 0 ns11 0 -1.24965224039
Ga11 ns11 0 ns10 0 1.24965224039
Ca12 ns12 0 1e-12
Ca13 ns13 0 1e-12
Ra12 ns12 0 3.75353660859 noise=0
Ra13 ns13 0 3.75353660859 noise=0
Ga12 ns12 0 ns13 0 -0.431489095244
Ga13 ns13 0 ns12 0 0.431489095244
Ca14 ns14 0 1e-12
Ra14 ns14 0 12.1731904857 noise=0
Ca15 ns15 0 1e-12
Ra15 ns15 0 531.342615159 noise=0
Ca16 ns16 0 1e-12
Ra16 ns16 0 4008.18525934 noise=0
Ca17 ns17 0 1e-12
Ra17 ns17 0 0.246835352493 noise=0
Ca18 ns18 0 1e-12
Ca19 ns19 0 1e-12
Ra18 ns18 0 5.85392236353 noise=0
Ra19 ns19 0 5.85392236353 noise=0
Ga18 ns18 0 ns19 0 -1.24965224039
Ga19 ns19 0 ns18 0 1.24965224039
Ca20 ns20 0 1e-12
Ca21 ns21 0 1e-12
Ra20 ns20 0 3.75353660859 noise=0
Ra21 ns21 0 3.75353660859 noise=0
Ga20 ns20 0 ns21 0 -0.431489095244
Ga21 ns21 0 ns20 0 0.431489095244
Ca22 ns22 0 1e-12
Ra22 ns22 0 12.1731904857 noise=0
Ca23 ns23 0 1e-12
Ra23 ns23 0 531.342615159 noise=0
Ca24 ns24 0 1e-12
Ra24 ns24 0 4008.18525934 noise=0
Ca25 ns25 0 1e-12
Ra25 ns25 0 0.246835352493 noise=0
Ca26 ns26 0 1e-12
Ca27 ns27 0 1e-12
Ra26 ns26 0 5.85392236353 noise=0
Ra27 ns27 0 5.85392236353 noise=0
Ga26 ns26 0 ns27 0 -1.24965224039
Ga27 ns27 0 ns26 0 1.24965224039
Ca28 ns28 0 1e-12
Ca29 ns29 0 1e-12
Ra28 ns28 0 3.75353660859 noise=0
Ra29 ns29 0 3.75353660859 noise=0
Ga28 ns28 0 ns29 0 -0.431489095244
Ga29 ns29 0 ns28 0 0.431489095244
Ca30 ns30 0 1e-12
Ra30 ns30 0 12.1731904857 noise=0
Ca31 ns31 0 1e-12
Ra31 ns31 0 531.342615159 noise=0
Ca32 ns32 0 1e-12
Ra32 ns32 0 4008.18525934 noise=0
Ca33 ns33 0 1e-12
Ra33 ns33 0 0.246835352493 noise=0
Ca34 ns34 0 1e-12
Ca35 ns35 0 1e-12
Ra34 ns34 0 5.85392236353 noise=0
Ra35 ns35 0 5.85392236353 noise=0
Ga34 ns34 0 ns35 0 -1.24965224039
Ga35 ns35 0 ns34 0 1.24965224039
Ca36 ns36 0 1e-12
Ca37 ns37 0 1e-12
Ra36 ns36 0 3.75353660859 noise=0
Ra37 ns37 0 3.75353660859 noise=0
Ga36 ns36 0 ns37 0 -0.431489095244
Ga37 ns37 0 ns36 0 0.431489095244
Ca38 ns38 0 1e-12
Ra38 ns38 0 12.1731904857 noise=0
Ca39 ns39 0 1e-12
Ra39 ns39 0 531.342615159 noise=0
Ca40 ns40 0 1e-12
Ra40 ns40 0 4008.18525934 noise=0
Ca41 ns41 0 1e-12
Ra41 ns41 0 0.246835352493 noise=0
Ca42 ns42 0 1e-12
Ca43 ns43 0 1e-12
Ra42 ns42 0 5.85392236353 noise=0
Ra43 ns43 0 5.85392236353 noise=0
Ga42 ns42 0 ns43 0 -1.24965224039
Ga43 ns43 0 ns42 0 1.24965224039
Ca44 ns44 0 1e-12
Ca45 ns45 0 1e-12
Ra44 ns44 0 3.75353660859 noise=0
Ra45 ns45 0 3.75353660859 noise=0
Ga44 ns44 0 ns45 0 -0.431489095244
Ga45 ns45 0 ns44 0 0.431489095244
Ca46 ns46 0 1e-12
Ra46 ns46 0 12.1731904857 noise=0
Ca47 ns47 0 1e-12
Ra47 ns47 0 531.342615159 noise=0
Ca48 ns48 0 1e-12
Ra48 ns48 0 4008.18525934 noise=0
Ca49 ns49 0 1e-12
Ra49 ns49 0 0.246835352493 noise=0
Ca50 ns50 0 1e-12
Ca51 ns51 0 1e-12
Ra50 ns50 0 5.85392236353 noise=0
Ra51 ns51 0 5.85392236353 noise=0
Ga50 ns50 0 ns51 0 -1.24965224039
Ga51 ns51 0 ns50 0 1.24965224039
Ca52 ns52 0 1e-12
Ca53 ns53 0 1e-12
Ra52 ns52 0 3.75353660859 noise=0
Ra53 ns53 0 3.75353660859 noise=0
Ga52 ns52 0 ns53 0 -0.431489095244
Ga53 ns53 0 ns52 0 0.431489095244
Ca54 ns54 0 1e-12
Ra54 ns54 0 12.1731904857 noise=0
Ca55 ns55 0 1e-12
Ra55 ns55 0 531.342615159 noise=0
Ca56 ns56 0 1e-12
Ra56 ns56 0 4008.18525934 noise=0
Ca57 ns57 0 1e-12
Ra57 ns57 0 0.246835352493 noise=0
Ca58 ns58 0 1e-12
Ca59 ns59 0 1e-12
Ra58 ns58 0 5.85392236353 noise=0
Ra59 ns59 0 5.85392236353 noise=0
Ga58 ns58 0 ns59 0 -1.24965224039
Ga59 ns59 0 ns58 0 1.24965224039
Ca60 ns60 0 1e-12
Ca61 ns61 0 1e-12
Ra60 ns60 0 3.75353660859 noise=0
Ra61 ns61 0 3.75353660859 noise=0
Ga60 ns60 0 ns61 0 -0.431489095244
Ga61 ns61 0 ns60 0 0.431489095244
Ca62 ns62 0 1e-12
Ra62 ns62 0 12.1731904857 noise=0
Ca63 ns63 0 1e-12
Ra63 ns63 0 531.342615159 noise=0
Ca64 ns64 0 1e-12
Ra64 ns64 0 4008.18525934 noise=0
Ca65 ns65 0 1e-12
Ra65 ns65 0 0.246835352493 noise=0
Ca66 ns66 0 1e-12
Ca67 ns67 0 1e-12
Ra66 ns66 0 5.85392236353 noise=0
Ra67 ns67 0 5.85392236353 noise=0
Ga66 ns66 0 ns67 0 -1.24965224039
Ga67 ns67 0 ns66 0 1.24965224039
Ca68 ns68 0 1e-12
Ca69 ns69 0 1e-12
Ra68 ns68 0 3.75353660859 noise=0
Ra69 ns69 0 3.75353660859 noise=0
Ga68 ns68 0 ns69 0 -0.431489095244
Ga69 ns69 0 ns68 0 0.431489095244
Ca70 ns70 0 1e-12
Ra70 ns70 0 12.1731904857 noise=0
Ca71 ns71 0 1e-12
Ra71 ns71 0 531.342615159 noise=0
Ca72 ns72 0 1e-12
Ra72 ns72 0 4008.18525934 noise=0
Ca73 ns73 0 1e-12
Ra73 ns73 0 0.246835352493 noise=0
Ca74 ns74 0 1e-12
Ca75 ns75 0 1e-12
Ra74 ns74 0 5.85392236353 noise=0
Ra75 ns75 0 5.85392236353 noise=0
Ga74 ns74 0 ns75 0 -1.24965224039
Ga75 ns75 0 ns74 0 1.24965224039
Ca76 ns76 0 1e-12
Ca77 ns77 0 1e-12
Ra76 ns76 0 3.75353660859 noise=0
Ra77 ns77 0 3.75353660859 noise=0
Ga76 ns76 0 ns77 0 -0.431489095244
Ga77 ns77 0 ns76 0 0.431489095244
Ca78 ns78 0 1e-12
Ra78 ns78 0 12.1731904857 noise=0
Ca79 ns79 0 1e-12
Ra79 ns79 0 531.342615159 noise=0
Ca80 ns80 0 1e-12
Ra80 ns80 0 4008.18525934 noise=0
Ca81 ns81 0 1e-12
Ra81 ns81 0 0.246835352493 noise=0
Ca82 ns82 0 1e-12
Ca83 ns83 0 1e-12
Ra82 ns82 0 5.85392236353 noise=0
Ra83 ns83 0 5.85392236353 noise=0
Ga82 ns82 0 ns83 0 -1.24965224039
Ga83 ns83 0 ns82 0 1.24965224039
Ca84 ns84 0 1e-12
Ca85 ns85 0 1e-12
Ra84 ns84 0 3.75353660859 noise=0
Ra85 ns85 0 3.75353660859 noise=0
Ga84 ns84 0 ns85 0 -0.431489095244
Ga85 ns85 0 ns84 0 0.431489095244
Ca86 ns86 0 1e-12
Ra86 ns86 0 12.1731904857 noise=0
Ca87 ns87 0 1e-12
Ra87 ns87 0 531.342615159 noise=0
Ca88 ns88 0 1e-12
Ra88 ns88 0 4008.18525934 noise=0
Ca89 ns89 0 1e-12
Ra89 ns89 0 0.246835352493 noise=0
Ca90 ns90 0 1e-12
Ca91 ns91 0 1e-12
Ra90 ns90 0 5.85392236353 noise=0
Ra91 ns91 0 5.85392236353 noise=0
Ga90 ns90 0 ns91 0 -1.24965224039
Ga91 ns91 0 ns90 0 1.24965224039
Ca92 ns92 0 1e-12
Ca93 ns93 0 1e-12
Ra92 ns92 0 3.75353660859 noise=0
Ra93 ns93 0 3.75353660859 noise=0
Ga92 ns92 0 ns93 0 -0.431489095244
Ga93 ns93 0 ns92 0 0.431489095244
Ca94 ns94 0 1e-12
Ra94 ns94 0 12.1731904857 noise=0
Ca95 ns95 0 1e-12
Ra95 ns95 0 531.342615159 noise=0
Ca96 ns96 0 1e-12
Ra96 ns96 0 4008.18525934 noise=0
Ca97 ns97 0 1e-12
Ra97 ns97 0 0.246835352493 noise=0
Ca98 ns98 0 1e-12
Ca99 ns99 0 1e-12
Ra98 ns98 0 5.85392236353 noise=0
Ra99 ns99 0 5.85392236353 noise=0
Ga98 ns98 0 ns99 0 -1.24965224039
Ga99 ns99 0 ns98 0 1.24965224039
Ca100 ns100 0 1e-12
Ca101 ns101 0 1e-12
Ra100 ns100 0 3.75353660859 noise=0
Ra101 ns101 0 3.75353660859 noise=0
Ga100 ns100 0 ns101 0 -0.431489095244
Ga101 ns101 0 ns100 0 0.431489095244
Ca102 ns102 0 1e-12
Ra102 ns102 0 12.1731904857 noise=0
Ca103 ns103 0 1e-12
Ra103 ns103 0 531.342615159 noise=0
Ca104 ns104 0 1e-12
Ra104 ns104 0 4008.18525934 noise=0
Ca105 ns105 0 1e-12
Ra105 ns105 0 0.246835352493 noise=0
Ca106 ns106 0 1e-12
Ca107 ns107 0 1e-12
Ra106 ns106 0 5.85392236353 noise=0
Ra107 ns107 0 5.85392236353 noise=0
Ga106 ns106 0 ns107 0 -1.24965224039
Ga107 ns107 0 ns106 0 1.24965224039
Ca108 ns108 0 1e-12
Ca109 ns109 0 1e-12
Ra108 ns108 0 3.75353660859 noise=0
Ra109 ns109 0 3.75353660859 noise=0
Ga108 ns108 0 ns109 0 -0.431489095244
Ga109 ns109 0 ns108 0 0.431489095244
Ca110 ns110 0 1e-12
Ra110 ns110 0 12.1731904857 noise=0
Ca111 ns111 0 1e-12
Ra111 ns111 0 531.342615159 noise=0
Ca112 ns112 0 1e-12
Ra112 ns112 0 4008.18525934 noise=0
Ca113 ns113 0 1e-12
Ra113 ns113 0 0.246835352493 noise=0
Ca114 ns114 0 1e-12
Ca115 ns115 0 1e-12
Ra114 ns114 0 5.85392236353 noise=0
Ra115 ns115 0 5.85392236353 noise=0
Ga114 ns114 0 ns115 0 -1.24965224039
Ga115 ns115 0 ns114 0 1.24965224039
Ca116 ns116 0 1e-12
Ca117 ns117 0 1e-12
Ra116 ns116 0 3.75353660859 noise=0
Ra117 ns117 0 3.75353660859 noise=0
Ga116 ns116 0 ns117 0 -0.431489095244
Ga117 ns117 0 ns116 0 0.431489095244
Ca118 ns118 0 1e-12
Ra118 ns118 0 12.1731904857 noise=0
Ca119 ns119 0 1e-12
Ra119 ns119 0 531.342615159 noise=0
Ca120 ns120 0 1e-12
Ra120 ns120 0 4008.18525934 noise=0
Ca121 ns121 0 1e-12
Ra121 ns121 0 0.246835352493 noise=0
Ca122 ns122 0 1e-12
Ca123 ns123 0 1e-12
Ra122 ns122 0 5.85392236353 noise=0
Ra123 ns123 0 5.85392236353 noise=0
Ga122 ns122 0 ns123 0 -1.24965224039
Ga123 ns123 0 ns122 0 1.24965224039
Ca124 ns124 0 1e-12
Ca125 ns125 0 1e-12
Ra124 ns124 0 3.75353660859 noise=0
Ra125 ns125 0 3.75353660859 noise=0
Ga124 ns124 0 ns125 0 -0.431489095244
Ga125 ns125 0 ns124 0 0.431489095244
Ca126 ns126 0 1e-12
Ra126 ns126 0 12.1731904857 noise=0
Ca127 ns127 0 1e-12
Ra127 ns127 0 531.342615159 noise=0
Ca128 ns128 0 1e-12
Ra128 ns128 0 4008.18525934 noise=0
Ca129 ns129 0 1e-12
Ra129 ns129 0 0.246835352493 noise=0
Ca130 ns130 0 1e-12
Ca131 ns131 0 1e-12
Ra130 ns130 0 5.85392236353 noise=0
Ra131 ns131 0 5.85392236353 noise=0
Ga130 ns130 0 ns131 0 -1.24965224039
Ga131 ns131 0 ns130 0 1.24965224039
Ca132 ns132 0 1e-12
Ca133 ns133 0 1e-12
Ra132 ns132 0 3.75353660859 noise=0
Ra133 ns133 0 3.75353660859 noise=0
Ga132 ns132 0 ns133 0 -0.431489095244
Ga133 ns133 0 ns132 0 0.431489095244
Ca134 ns134 0 1e-12
Ra134 ns134 0 12.1731904857 noise=0
Ca135 ns135 0 1e-12
Ra135 ns135 0 531.342615159 noise=0
Ca136 ns136 0 1e-12
Ra136 ns136 0 4008.18525934 noise=0
Ca137 ns137 0 1e-12
Ra137 ns137 0 0.246835352493 noise=0
Ca138 ns138 0 1e-12
Ca139 ns139 0 1e-12
Ra138 ns138 0 5.85392236353 noise=0
Ra139 ns139 0 5.85392236353 noise=0
Ga138 ns138 0 ns139 0 -1.24965224039
Ga139 ns139 0 ns138 0 1.24965224039
Ca140 ns140 0 1e-12
Ca141 ns141 0 1e-12
Ra140 ns140 0 3.75353660859 noise=0
Ra141 ns141 0 3.75353660859 noise=0
Ga140 ns140 0 ns141 0 -0.431489095244
Ga141 ns141 0 ns140 0 0.431489095244
Ca142 ns142 0 1e-12
Ra142 ns142 0 12.1731904857 noise=0
Ca143 ns143 0 1e-12
Ra143 ns143 0 531.342615159 noise=0
Ca144 ns144 0 1e-12
Ra144 ns144 0 4008.18525934 noise=0
Ca145 ns145 0 1e-12
Ra145 ns145 0 0.246835352493 noise=0
Ca146 ns146 0 1e-12
Ca147 ns147 0 1e-12
Ra146 ns146 0 5.85392236353 noise=0
Ra147 ns147 0 5.85392236353 noise=0
Ga146 ns146 0 ns147 0 -1.24965224039
Ga147 ns147 0 ns146 0 1.24965224039
Ca148 ns148 0 1e-12
Ca149 ns149 0 1e-12
Ra148 ns148 0 3.75353660859 noise=0
Ra149 ns149 0 3.75353660859 noise=0
Ga148 ns148 0 ns149 0 -0.431489095244
Ga149 ns149 0 ns148 0 0.431489095244
Ca150 ns150 0 1e-12
Ra150 ns150 0 12.1731904857 noise=0
Ca151 ns151 0 1e-12
Ra151 ns151 0 531.342615159 noise=0
Ca152 ns152 0 1e-12
Ra152 ns152 0 4008.18525934 noise=0
Ca153 ns153 0 1e-12
Ra153 ns153 0 0.246835352493 noise=0
Ca154 ns154 0 1e-12
Ca155 ns155 0 1e-12
Ra154 ns154 0 5.85392236353 noise=0
Ra155 ns155 0 5.85392236353 noise=0
Ga154 ns154 0 ns155 0 -1.24965224039
Ga155 ns155 0 ns154 0 1.24965224039
Ca156 ns156 0 1e-12
Ca157 ns157 0 1e-12
Ra156 ns156 0 3.75353660859 noise=0
Ra157 ns157 0 3.75353660859 noise=0
Ga156 ns156 0 ns157 0 -0.431489095244
Ga157 ns157 0 ns156 0 0.431489095244
Ca158 ns158 0 1e-12
Ra158 ns158 0 12.1731904857 noise=0
Ca159 ns159 0 1e-12
Ra159 ns159 0 531.342615159 noise=0
Ca160 ns160 0 1e-12
Ra160 ns160 0 4008.18525934 noise=0
Ca161 ns161 0 1e-12
Ra161 ns161 0 0.246835352493 noise=0
Ca162 ns162 0 1e-12
Ca163 ns163 0 1e-12
Ra162 ns162 0 5.85392236353 noise=0
Ra163 ns163 0 5.85392236353 noise=0
Ga162 ns162 0 ns163 0 -1.24965224039
Ga163 ns163 0 ns162 0 1.24965224039
Ca164 ns164 0 1e-12
Ca165 ns165 0 1e-12
Ra164 ns164 0 3.75353660859 noise=0
Ra165 ns165 0 3.75353660859 noise=0
Ga164 ns164 0 ns165 0 -0.431489095244
Ga165 ns165 0 ns164 0 0.431489095244
Ca166 ns166 0 1e-12
Ra166 ns166 0 12.1731904857 noise=0
Ca167 ns167 0 1e-12
Ra167 ns167 0 531.342615159 noise=0
Ca168 ns168 0 1e-12
Ra168 ns168 0 4008.18525934 noise=0
Ca169 ns169 0 1e-12
Ra169 ns169 0 0.246835352493 noise=0
Ca170 ns170 0 1e-12
Ca171 ns171 0 1e-12
Ra170 ns170 0 5.85392236353 noise=0
Ra171 ns171 0 5.85392236353 noise=0
Ga170 ns170 0 ns171 0 -1.24965224039
Ga171 ns171 0 ns170 0 1.24965224039
Ca172 ns172 0 1e-12
Ca173 ns173 0 1e-12
Ra172 ns172 0 3.75353660859 noise=0
Ra173 ns173 0 3.75353660859 noise=0
Ga172 ns172 0 ns173 0 -0.431489095244
Ga173 ns173 0 ns172 0 0.431489095244
Ca174 ns174 0 1e-12
Ra174 ns174 0 12.1731904857 noise=0
Ca175 ns175 0 1e-12
Ra175 ns175 0 531.342615159 noise=0
Ca176 ns176 0 1e-12
Ra176 ns176 0 4008.18525934 noise=0
Ca177 ns177 0 1e-12
Ra177 ns177 0 0.246835352493 noise=0
Ca178 ns178 0 1e-12
Ca179 ns179 0 1e-12
Ra178 ns178 0 5.85392236353 noise=0
Ra179 ns179 0 5.85392236353 noise=0
Ga178 ns178 0 ns179 0 -1.24965224039
Ga179 ns179 0 ns178 0 1.24965224039
Ca180 ns180 0 1e-12
Ca181 ns181 0 1e-12
Ra180 ns180 0 3.75353660859 noise=0
Ra181 ns181 0 3.75353660859 noise=0
Ga180 ns180 0 ns181 0 -0.431489095244
Ga181 ns181 0 ns180 0 0.431489095244
Ca182 ns182 0 1e-12
Ra182 ns182 0 12.1731904857 noise=0
Ca183 ns183 0 1e-12
Ra183 ns183 0 531.342615159 noise=0
Ca184 ns184 0 1e-12
Ra184 ns184 0 4008.18525934 noise=0
Ca185 ns185 0 1e-12
Ra185 ns185 0 0.246835352493 noise=0
Ca186 ns186 0 1e-12
Ca187 ns187 0 1e-12
Ra186 ns186 0 5.85392236353 noise=0
Ra187 ns187 0 5.85392236353 noise=0
Ga186 ns186 0 ns187 0 -1.24965224039
Ga187 ns187 0 ns186 0 1.24965224039
Ca188 ns188 0 1e-12
Ca189 ns189 0 1e-12
Ra188 ns188 0 3.75353660859 noise=0
Ra189 ns189 0 3.75353660859 noise=0
Ga188 ns188 0 ns189 0 -0.431489095244
Ga189 ns189 0 ns188 0 0.431489095244
Ca190 ns190 0 1e-12
Ra190 ns190 0 12.1731904857 noise=0
Ca191 ns191 0 1e-12
Ra191 ns191 0 531.342615159 noise=0
Ca192 ns192 0 1e-12
Ra192 ns192 0 4008.18525934 noise=0
Ca193 ns193 0 1e-12
Ra193 ns193 0 0.246835352493 noise=0
Ca194 ns194 0 1e-12
Ca195 ns195 0 1e-12
Ra194 ns194 0 5.85392236353 noise=0
Ra195 ns195 0 5.85392236353 noise=0
Ga194 ns194 0 ns195 0 -1.24965224039
Ga195 ns195 0 ns194 0 1.24965224039
Ca196 ns196 0 1e-12
Ca197 ns197 0 1e-12
Ra196 ns196 0 3.75353660859 noise=0
Ra197 ns197 0 3.75353660859 noise=0
Ga196 ns196 0 ns197 0 -0.431489095244
Ga197 ns197 0 ns196 0 0.431489095244
Ca198 ns198 0 1e-12
Ra198 ns198 0 12.1731904857 noise=0
Ca199 ns199 0 1e-12
Ra199 ns199 0 531.342615159 noise=0
Ca200 ns200 0 1e-12
Ra200 ns200 0 4008.18525934 noise=0
Ca201 ns201 0 1e-12
Ra201 ns201 0 0.246835352493 noise=0
Ca202 ns202 0 1e-12
Ca203 ns203 0 1e-12
Ra202 ns202 0 5.85392236353 noise=0
Ra203 ns203 0 5.85392236353 noise=0
Ga202 ns202 0 ns203 0 -1.24965224039
Ga203 ns203 0 ns202 0 1.24965224039
Ca204 ns204 0 1e-12
Ca205 ns205 0 1e-12
Ra204 ns204 0 3.75353660859 noise=0
Ra205 ns205 0 3.75353660859 noise=0
Ga204 ns204 0 ns205 0 -0.431489095244
Ga205 ns205 0 ns204 0 0.431489095244
Ca206 ns206 0 1e-12
Ra206 ns206 0 12.1731904857 noise=0
Ca207 ns207 0 1e-12
Ra207 ns207 0 531.342615159 noise=0
Ca208 ns208 0 1e-12
Ra208 ns208 0 4008.18525934 noise=0
Ca209 ns209 0 1e-12
Ra209 ns209 0 0.246835352493 noise=0
Ca210 ns210 0 1e-12
Ca211 ns211 0 1e-12
Ra210 ns210 0 5.85392236353 noise=0
Ra211 ns211 0 5.85392236353 noise=0
Ga210 ns210 0 ns211 0 -1.24965224039
Ga211 ns211 0 ns210 0 1.24965224039
Ca212 ns212 0 1e-12
Ca213 ns213 0 1e-12
Ra212 ns212 0 3.75353660859 noise=0
Ra213 ns213 0 3.75353660859 noise=0
Ga212 ns212 0 ns213 0 -0.431489095244
Ga213 ns213 0 ns212 0 0.431489095244
Ca214 ns214 0 1e-12
Ra214 ns214 0 12.1731904857 noise=0
Ca215 ns215 0 1e-12
Ra215 ns215 0 531.342615159 noise=0
Ca216 ns216 0 1e-12
Ra216 ns216 0 4008.18525934 noise=0
Ca217 ns217 0 1e-12
Ra217 ns217 0 0.246835352493 noise=0
Ca218 ns218 0 1e-12
Ca219 ns219 0 1e-12
Ra218 ns218 0 5.85392236353 noise=0
Ra219 ns219 0 5.85392236353 noise=0
Ga218 ns218 0 ns219 0 -1.24965224039
Ga219 ns219 0 ns218 0 1.24965224039
Ca220 ns220 0 1e-12
Ca221 ns221 0 1e-12
Ra220 ns220 0 3.75353660859 noise=0
Ra221 ns221 0 3.75353660859 noise=0
Ga220 ns220 0 ns221 0 -0.431489095244
Ga221 ns221 0 ns220 0 0.431489095244
Ca222 ns222 0 1e-12
Ra222 ns222 0 12.1731904857 noise=0
Ca223 ns223 0 1e-12
Ra223 ns223 0 531.342615159 noise=0
Ca224 ns224 0 1e-12
Ra224 ns224 0 4008.18525934 noise=0
Ca225 ns225 0 1e-12
Ra225 ns225 0 0.246835352493 noise=0
Ca226 ns226 0 1e-12
Ca227 ns227 0 1e-12
Ra226 ns226 0 5.85392236353 noise=0
Ra227 ns227 0 5.85392236353 noise=0
Ga226 ns226 0 ns227 0 -1.24965224039
Ga227 ns227 0 ns226 0 1.24965224039
Ca228 ns228 0 1e-12
Ca229 ns229 0 1e-12
Ra228 ns228 0 3.75353660859 noise=0
Ra229 ns229 0 3.75353660859 noise=0
Ga228 ns228 0 ns229 0 -0.431489095244
Ga229 ns229 0 ns228 0 0.431489095244
Ca230 ns230 0 1e-12
Ra230 ns230 0 12.1731904857 noise=0
Ca231 ns231 0 1e-12
Ra231 ns231 0 531.342615159 noise=0
Ca232 ns232 0 1e-12
Ra232 ns232 0 4008.18525934 noise=0
Ca233 ns233 0 1e-12
Ra233 ns233 0 0.246835352493 noise=0
Ca234 ns234 0 1e-12
Ca235 ns235 0 1e-12
Ra234 ns234 0 5.85392236353 noise=0
Ra235 ns235 0 5.85392236353 noise=0
Ga234 ns234 0 ns235 0 -1.24965224039
Ga235 ns235 0 ns234 0 1.24965224039
Ca236 ns236 0 1e-12
Ca237 ns237 0 1e-12
Ra236 ns236 0 3.75353660859 noise=0
Ra237 ns237 0 3.75353660859 noise=0
Ga236 ns236 0 ns237 0 -0.431489095244
Ga237 ns237 0 ns236 0 0.431489095244
Ca238 ns238 0 1e-12
Ra238 ns238 0 12.1731904857 noise=0
Ca239 ns239 0 1e-12
Ra239 ns239 0 531.342615159 noise=0
Ca240 ns240 0 1e-12
Ra240 ns240 0 4008.18525934 noise=0
Ca241 ns241 0 1e-12
Ra241 ns241 0 0.246835352493 noise=0
Ca242 ns242 0 1e-12
Ca243 ns243 0 1e-12
Ra242 ns242 0 5.85392236353 noise=0
Ra243 ns243 0 5.85392236353 noise=0
Ga242 ns242 0 ns243 0 -1.24965224039
Ga243 ns243 0 ns242 0 1.24965224039
Ca244 ns244 0 1e-12
Ca245 ns245 0 1e-12
Ra244 ns244 0 3.75353660859 noise=0
Ra245 ns245 0 3.75353660859 noise=0
Ga244 ns244 0 ns245 0 -0.431489095244
Ga245 ns245 0 ns244 0 0.431489095244
Ca246 ns246 0 1e-12
Ra246 ns246 0 12.1731904857 noise=0
Ca247 ns247 0 1e-12
Ra247 ns247 0 531.342615159 noise=0
Ca248 ns248 0 1e-12
Ra248 ns248 0 4008.18525934 noise=0
Ca249 ns249 0 1e-12
Ra249 ns249 0 0.246835352493 noise=0
Ca250 ns250 0 1e-12
Ca251 ns251 0 1e-12
Ra250 ns250 0 5.85392236353 noise=0
Ra251 ns251 0 5.85392236353 noise=0
Ga250 ns250 0 ns251 0 -1.24965224039
Ga251 ns251 0 ns250 0 1.24965224039
Ca252 ns252 0 1e-12
Ca253 ns253 0 1e-12
Ra252 ns252 0 3.75353660859 noise=0
Ra253 ns253 0 3.75353660859 noise=0
Ga252 ns252 0 ns253 0 -0.431489095244
Ga253 ns253 0 ns252 0 0.431489095244
Ca254 ns254 0 1e-12
Ra254 ns254 0 12.1731904857 noise=0
Ca255 ns255 0 1e-12
Ra255 ns255 0 531.342615159 noise=0
Ca256 ns256 0 1e-12
Ra256 ns256 0 4008.18525934 noise=0

Gb1_1 ns1 0 ni1 0 -4.05128353739
Gb2_1 ns2 0 ni1 0 1.17655154414
Gb3_1 ns3 0 ni1 0 0.705584069575
Gb4_1 ns4 0 ni1 0 -0.436081647803
Gb5_1 ns5 0 ni1 0 0.258977266879
Gb6_1 ns6 0 ni1 0 -0.0821477328543
Gb7_1 ns7 0 ni1 0 0.00188202483947
Gb8_1 ns8 0 ni1 0 -0.000249489466004
Gb9_2 ns9 0 ni2 0 -4.05128353739
Gb10_2 ns10 0 ni2 0 1.17655154414
Gb11_2 ns11 0 ni2 0 0.705584069575
Gb12_2 ns12 0 ni2 0 -0.436081647803
Gb13_2 ns13 0 ni2 0 0.258977266879
Gb14_2 ns14 0 ni2 0 -0.0821477328543
Gb15_2 ns15 0 ni2 0 0.00188202483947
Gb16_2 ns16 0 ni2 0 -0.000249489466004
Gb17_3 ns17 0 ni3 0 -4.05128353739
Gb18_3 ns18 0 ni3 0 1.17655154414
Gb19_3 ns19 0 ni3 0 0.705584069575
Gb20_3 ns20 0 ni3 0 -0.436081647803
Gb21_3 ns21 0 ni3 0 0.258977266879
Gb22_3 ns22 0 ni3 0 -0.0821477328543
Gb23_3 ns23 0 ni3 0 0.00188202483947
Gb24_3 ns24 0 ni3 0 -0.000249489466004
Gb25_4 ns25 0 ni4 0 -4.05128353739
Gb26_4 ns26 0 ni4 0 1.17655154414
Gb27_4 ns27 0 ni4 0 0.705584069575
Gb28_4 ns28 0 ni4 0 -0.436081647803
Gb29_4 ns29 0 ni4 0 0.258977266879
Gb30_4 ns30 0 ni4 0 -0.0821477328543
Gb31_4 ns31 0 ni4 0 0.00188202483947
Gb32_4 ns32 0 ni4 0 -0.000249489466004
Gb33_5 ns33 0 ni5 0 -4.05128353739
Gb34_5 ns34 0 ni5 0 1.17655154414
Gb35_5 ns35 0 ni5 0 0.705584069575
Gb36_5 ns36 0 ni5 0 -0.436081647803
Gb37_5 ns37 0 ni5 0 0.258977266879
Gb38_5 ns38 0 ni5 0 -0.0821477328543
Gb39_5 ns39 0 ni5 0 0.00188202483947
Gb40_5 ns40 0 ni5 0 -0.000249489466004
Gb41_6 ns41 0 ni6 0 -4.05128353739
Gb42_6 ns42 0 ni6 0 1.17655154414
Gb43_6 ns43 0 ni6 0 0.705584069575
Gb44_6 ns44 0 ni6 0 -0.436081647803
Gb45_6 ns45 0 ni6 0 0.258977266879
Gb46_6 ns46 0 ni6 0 -0.0821477328543
Gb47_6 ns47 0 ni6 0 0.00188202483947
Gb48_6 ns48 0 ni6 0 -0.000249489466004
Gb49_7 ns49 0 ni7 0 -4.05128353739
Gb50_7 ns50 0 ni7 0 1.17655154414
Gb51_7 ns51 0 ni7 0 0.705584069575
Gb52_7 ns52 0 ni7 0 -0.436081647803
Gb53_7 ns53 0 ni7 0 0.258977266879
Gb54_7 ns54 0 ni7 0 -0.0821477328543
Gb55_7 ns55 0 ni7 0 0.00188202483947
Gb56_7 ns56 0 ni7 0 -0.000249489466004
Gb57_8 ns57 0 ni8 0 -4.05128353739
Gb58_8 ns58 0 ni8 0 1.17655154414
Gb59_8 ns59 0 ni8 0 0.705584069575
Gb60_8 ns60 0 ni8 0 -0.436081647803
Gb61_8 ns61 0 ni8 0 0.258977266879
Gb62_8 ns62 0 ni8 0 -0.0821477328543
Gb63_8 ns63 0 ni8 0 0.00188202483947
Gb64_8 ns64 0 ni8 0 -0.000249489466004
Gb65_9 ns65 0 ni9 0 -4.05128353739
Gb66_9 ns66 0 ni9 0 1.17655154414
Gb67_9 ns67 0 ni9 0 0.705584069575
Gb68_9 ns68 0 ni9 0 -0.436081647803
Gb69_9 ns69 0 ni9 0 0.258977266879
Gb70_9 ns70 0 ni9 0 -0.0821477328543
Gb71_9 ns71 0 ni9 0 0.00188202483947
Gb72_9 ns72 0 ni9 0 -0.000249489466004
Gb73_10 ns73 0 ni10 0 -4.05128353739
Gb74_10 ns74 0 ni10 0 1.17655154414
Gb75_10 ns75 0 ni10 0 0.705584069575
Gb76_10 ns76 0 ni10 0 -0.436081647803
Gb77_10 ns77 0 ni10 0 0.258977266879
Gb78_10 ns78 0 ni10 0 -0.0821477328543
Gb79_10 ns79 0 ni10 0 0.00188202483947
Gb80_10 ns80 0 ni10 0 -0.000249489466004
Gb81_11 ns81 0 ni11 0 -4.05128353739
Gb82_11 ns82 0 ni11 0 1.17655154414
Gb83_11 ns83 0 ni11 0 0.705584069575
Gb84_11 ns84 0 ni11 0 -0.436081647803
Gb85_11 ns85 0 ni11 0 0.258977266879
Gb86_11 ns86 0 ni11 0 -0.0821477328543
Gb87_11 ns87 0 ni11 0 0.00188202483947
Gb88_11 ns88 0 ni11 0 -0.000249489466004
Gb89_12 ns89 0 ni12 0 -4.05128353739
Gb90_12 ns90 0 ni12 0 1.17655154414
Gb91_12 ns91 0 ni12 0 0.705584069575
Gb92_12 ns92 0 ni12 0 -0.436081647803
Gb93_12 ns93 0 ni12 0 0.258977266879
Gb94_12 ns94 0 ni12 0 -0.0821477328543
Gb95_12 ns95 0 ni12 0 0.00188202483947
Gb96_12 ns96 0 ni12 0 -0.000249489466004
Gb97_13 ns97 0 ni13 0 -4.05128353739
Gb98_13 ns98 0 ni13 0 1.17655154414
Gb99_13 ns99 0 ni13 0 0.705584069575
Gb100_13 ns100 0 ni13 0 -0.436081647803
Gb101_13 ns101 0 ni13 0 0.258977266879
Gb102_13 ns102 0 ni13 0 -0.0821477328543
Gb103_13 ns103 0 ni13 0 0.00188202483947
Gb104_13 ns104 0 ni13 0 -0.000249489466004
Gb105_14 ns105 0 ni14 0 -4.05128353739
Gb106_14 ns106 0 ni14 0 1.17655154414
Gb107_14 ns107 0 ni14 0 0.705584069575
Gb108_14 ns108 0 ni14 0 -0.436081647803
Gb109_14 ns109 0 ni14 0 0.258977266879
Gb110_14 ns110 0 ni14 0 -0.0821477328543
Gb111_14 ns111 0 ni14 0 0.00188202483947
Gb112_14 ns112 0 ni14 0 -0.000249489466004
Gb113_15 ns113 0 ni15 0 -4.05128353739
Gb114_15 ns114 0 ni15 0 1.17655154414
Gb115_15 ns115 0 ni15 0 0.705584069575
Gb116_15 ns116 0 ni15 0 -0.436081647803
Gb117_15 ns117 0 ni15 0 0.258977266879
Gb118_15 ns118 0 ni15 0 -0.0821477328543
Gb119_15 ns119 0 ni15 0 0.00188202483947
Gb120_15 ns120 0 ni15 0 -0.000249489466004
Gb121_16 ns121 0 ni16 0 -4.05128353739
Gb122_16 ns122 0 ni16 0 1.17655154414
Gb123_16 ns123 0 ni16 0 0.705584069575
Gb124_16 ns124 0 ni16 0 -0.436081647803
Gb125_16 ns125 0 ni16 0 0.258977266879
Gb126_16 ns126 0 ni16 0 -0.0821477328543
Gb127_16 ns127 0 ni16 0 0.00188202483947
Gb128_16 ns128 0 ni16 0 -0.000249489466004
Gb129_17 ns129 0 ni17 0 -4.05128353739
Gb130_17 ns130 0 ni17 0 1.17655154414
Gb131_17 ns131 0 ni17 0 0.705584069575
Gb132_17 ns132 0 ni17 0 -0.436081647803
Gb133_17 ns133 0 ni17 0 0.258977266879
Gb134_17 ns134 0 ni17 0 -0.0821477328543
Gb135_17 ns135 0 ni17 0 0.00188202483947
Gb136_17 ns136 0 ni17 0 -0.000249489466004
Gb137_18 ns137 0 ni18 0 -4.05128353739
Gb138_18 ns138 0 ni18 0 1.17655154414
Gb139_18 ns139 0 ni18 0 0.705584069575
Gb140_18 ns140 0 ni18 0 -0.436081647803
Gb141_18 ns141 0 ni18 0 0.258977266879
Gb142_18 ns142 0 ni18 0 -0.0821477328543
Gb143_18 ns143 0 ni18 0 0.00188202483947
Gb144_18 ns144 0 ni18 0 -0.000249489466004
Gb145_19 ns145 0 ni19 0 -4.05128353739
Gb146_19 ns146 0 ni19 0 1.17655154414
Gb147_19 ns147 0 ni19 0 0.705584069575
Gb148_19 ns148 0 ni19 0 -0.436081647803
Gb149_19 ns149 0 ni19 0 0.258977266879
Gb150_19 ns150 0 ni19 0 -0.0821477328543
Gb151_19 ns151 0 ni19 0 0.00188202483947
Gb152_19 ns152 0 ni19 0 -0.000249489466004
Gb153_20 ns153 0 ni20 0 -4.05128353739
Gb154_20 ns154 0 ni20 0 1.17655154414
Gb155_20 ns155 0 ni20 0 0.705584069575
Gb156_20 ns156 0 ni20 0 -0.436081647803
Gb157_20 ns157 0 ni20 0 0.258977266879
Gb158_20 ns158 0 ni20 0 -0.0821477328543
Gb159_20 ns159 0 ni20 0 0.00188202483947
Gb160_20 ns160 0 ni20 0 -0.000249489466004
Gb161_21 ns161 0 ni21 0 -4.05128353739
Gb162_21 ns162 0 ni21 0 1.17655154414
Gb163_21 ns163 0 ni21 0 0.705584069575
Gb164_21 ns164 0 ni21 0 -0.436081647803
Gb165_21 ns165 0 ni21 0 0.258977266879
Gb166_21 ns166 0 ni21 0 -0.0821477328543
Gb167_21 ns167 0 ni21 0 0.00188202483947
Gb168_21 ns168 0 ni21 0 -0.000249489466004
Gb169_22 ns169 0 ni22 0 -4.05128353739
Gb170_22 ns170 0 ni22 0 1.17655154414
Gb171_22 ns171 0 ni22 0 0.705584069575
Gb172_22 ns172 0 ni22 0 -0.436081647803
Gb173_22 ns173 0 ni22 0 0.258977266879
Gb174_22 ns174 0 ni22 0 -0.0821477328543
Gb175_22 ns175 0 ni22 0 0.00188202483947
Gb176_22 ns176 0 ni22 0 -0.000249489466004
Gb177_23 ns177 0 ni23 0 -4.05128353739
Gb178_23 ns178 0 ni23 0 1.17655154414
Gb179_23 ns179 0 ni23 0 0.705584069575
Gb180_23 ns180 0 ni23 0 -0.436081647803
Gb181_23 ns181 0 ni23 0 0.258977266879
Gb182_23 ns182 0 ni23 0 -0.0821477328543
Gb183_23 ns183 0 ni23 0 0.00188202483947
Gb184_23 ns184 0 ni23 0 -0.000249489466004
Gb185_24 ns185 0 ni24 0 -4.05128353739
Gb186_24 ns186 0 ni24 0 1.17655154414
Gb187_24 ns187 0 ni24 0 0.705584069575
Gb188_24 ns188 0 ni24 0 -0.436081647803
Gb189_24 ns189 0 ni24 0 0.258977266879
Gb190_24 ns190 0 ni24 0 -0.0821477328543
Gb191_24 ns191 0 ni24 0 0.00188202483947
Gb192_24 ns192 0 ni24 0 -0.000249489466004
Gb193_25 ns193 0 ni25 0 -4.05128353739
Gb194_25 ns194 0 ni25 0 1.17655154414
Gb195_25 ns195 0 ni25 0 0.705584069575
Gb196_25 ns196 0 ni25 0 -0.436081647803
Gb197_25 ns197 0 ni25 0 0.258977266879
Gb198_25 ns198 0 ni25 0 -0.0821477328543
Gb199_25 ns199 0 ni25 0 0.00188202483947
Gb200_25 ns200 0 ni25 0 -0.000249489466004
Gb201_26 ns201 0 ni26 0 -4.05128353739
Gb202_26 ns202 0 ni26 0 1.17655154414
Gb203_26 ns203 0 ni26 0 0.705584069575
Gb204_26 ns204 0 ni26 0 -0.436081647803
Gb205_26 ns205 0 ni26 0 0.258977266879
Gb206_26 ns206 0 ni26 0 -0.0821477328543
Gb207_26 ns207 0 ni26 0 0.00188202483947
Gb208_26 ns208 0 ni26 0 -0.000249489466004
Gb209_27 ns209 0 ni27 0 -4.05128353739
Gb210_27 ns210 0 ni27 0 1.17655154414
Gb211_27 ns211 0 ni27 0 0.705584069575
Gb212_27 ns212 0 ni27 0 -0.436081647803
Gb213_27 ns213 0 ni27 0 0.258977266879
Gb214_27 ns214 0 ni27 0 -0.0821477328543
Gb215_27 ns215 0 ni27 0 0.00188202483947
Gb216_27 ns216 0 ni27 0 -0.000249489466004
Gb217_28 ns217 0 ni28 0 -4.05128353739
Gb218_28 ns218 0 ni28 0 1.17655154414
Gb219_28 ns219 0 ni28 0 0.705584069575
Gb220_28 ns220 0 ni28 0 -0.436081647803
Gb221_28 ns221 0 ni28 0 0.258977266879
Gb222_28 ns222 0 ni28 0 -0.0821477328543
Gb223_28 ns223 0 ni28 0 0.00188202483947
Gb224_28 ns224 0 ni28 0 -0.000249489466004
Gb225_29 ns225 0 ni29 0 -4.05128353739
Gb226_29 ns226 0 ni29 0 1.17655154414
Gb227_29 ns227 0 ni29 0 0.705584069575
Gb228_29 ns228 0 ni29 0 -0.436081647803
Gb229_29 ns229 0 ni29 0 0.258977266879
Gb230_29 ns230 0 ni29 0 -0.0821477328543
Gb231_29 ns231 0 ni29 0 0.00188202483947
Gb232_29 ns232 0 ni29 0 -0.000249489466004
Gb233_30 ns233 0 ni30 0 -4.05128353739
Gb234_30 ns234 0 ni30 0 1.17655154414
Gb235_30 ns235 0 ni30 0 0.705584069575
Gb236_30 ns236 0 ni30 0 -0.436081647803
Gb237_30 ns237 0 ni30 0 0.258977266879
Gb238_30 ns238 0 ni30 0 -0.0821477328543
Gb239_30 ns239 0 ni30 0 0.00188202483947
Gb240_30 ns240 0 ni30 0 -0.000249489466004
Gb241_31 ns241 0 ni31 0 -4.05128353739
Gb242_31 ns242 0 ni31 0 1.17655154414
Gb243_31 ns243 0 ni31 0 0.705584069575
Gb244_31 ns244 0 ni31 0 -0.436081647803
Gb245_31 ns245 0 ni31 0 0.258977266879
Gb246_31 ns246 0 ni31 0 -0.0821477328543
Gb247_31 ns247 0 ni31 0 0.00188202483947
Gb248_31 ns248 0 ni31 0 -0.000249489466004
Gb249_32 ns249 0 ni32 0 -4.05128353739
Gb250_32 ns250 0 ni32 0 1.17655154414
Gb251_32 ns251 0 ni32 0 0.705584069575
Gb252_32 ns252 0 ni32 0 -0.436081647803
Gb253_32 ns253 0 ni32 0 0.258977266879
Gb254_32 ns254 0 ni32 0 -0.0821477328543
Gb255_32 ns255 0 ni32 0 0.00188202483947
Gb256_32 ns256 0 ni32 0 -0.000249489466004

Gc1_1 0 n2 ns1 0 0.00507615873051
Gc1_2 0 n2 ns2 0 -0.000100404574865
Gc1_3 0 n2 ns3 0 0.000615793769192
Gc1_4 0 n2 ns4 0 0.00100079419327
Gc1_5 0 n2 ns5 0 0.000370180865665
Gc1_6 0 n2 ns6 0 -7.10856477935e-05
Gc1_7 0 n2 ns7 0 1.66435089871e-05
Gc1_8 0 n2 ns8 0 0.000582222339371
Gc1_9 0 n2 ns9 0 0.00170344945102
Gc1_10 0 n2 ns10 0 -2.7551388872e-05
Gc1_11 0 n2 ns11 0 -4.37654841207e-06
Gc1_12 0 n2 ns12 0 0.000271099227809
Gc1_13 0 n2 ns13 0 -1.63421590458e-05
Gc1_14 0 n2 ns14 0 -0.000120082274237
Gc1_15 0 n2 ns15 0 9.55288533273e-05
Gc1_16 0 n2 ns16 0 -8.89608401891e-05
Gc1_17 0 n2 ns17 0 -0.00059012372801
Gc1_18 0 n2 ns18 0 1.25618860156e-05
Gc1_19 0 n2 ns19 0 -8.71731718617e-05
Gc1_20 0 n2 ns20 0 -0.000146208400641
Gc1_21 0 n2 ns21 0 -0.000127315799585
Gc1_22 0 n2 ns22 0 -4.84194511262e-05
Gc1_23 0 n2 ns23 0 -1.67327972321e-05
Gc1_24 0 n2 ns24 0 -5.48870170322e-05
Gc1_25 0 n2 ns25 0 6.19520587657e-06
Gc1_26 0 n2 ns26 0 2.3784522811e-07
Gc1_27 0 n2 ns27 0 4.43393574485e-07
Gc1_28 0 n2 ns28 0 -5.71073410869e-06
Gc1_29 0 n2 ns29 0 -7.17293235846e-06
Gc1_30 0 n2 ns30 0 8.20625932242e-06
Gc1_31 0 n2 ns31 0 -1.44159389408e-07
Gc1_32 0 n2 ns32 0 -8.97282516464e-07
Gc1_33 0 n2 ns33 0 1.20370228915e-05
Gc1_34 0 n2 ns34 0 -1.22155562566e-07
Gc1_35 0 n2 ns35 0 1.70327311833e-06
Gc1_36 0 n2 ns36 0 -1.59210198577e-06
Gc1_37 0 n2 ns37 0 -2.74622201324e-06
Gc1_38 0 n2 ns38 0 3.41159763809e-06
Gc1_39 0 n2 ns39 0 1.06493496518e-07
Gc1_40 0 n2 ns40 0 6.31246642884e-07
Gc1_41 0 n2 ns41 0 -2.45215524068e-05
Gc1_42 0 n2 ns42 0 5.30778522145e-07
Gc1_43 0 n2 ns43 0 -3.08396167442e-06
Gc1_44 0 n2 ns44 0 -7.06056896579e-06
Gc1_45 0 n2 ns45 0 -8.13413540933e-06
Gc1_46 0 n2 ns46 0 -1.08609338201e-06
Gc1_47 0 n2 ns47 0 -1.11224817746e-06
Gc1_48 0 n2 ns48 0 -1.866996702e-06
Gc1_49 0 n2 ns49 0 -1.32249483454e-05
Gc1_50 0 n2 ns50 0 2.83410547229e-07
Gc1_51 0 n2 ns51 0 -1.61625567114e-06
Gc1_52 0 n2 ns52 0 -2.84037829234e-06
Gc1_53 0 n2 ns53 0 -4.75881817387e-06
Gc1_54 0 n2 ns54 0 -1.80587315176e-07
Gc1_55 0 n2 ns55 0 -7.15829998279e-07
Gc1_56 0 n2 ns56 0 -1.02093447752e-06
Gc1_57 0 n2 ns57 0 -3.79933865695e-06
Gc1_58 0 n2 ns58 0 9.26575079366e-08
Gc1_59 0 n2 ns59 0 -4.6585241826e-07
Gc1_60 0 n2 ns60 0 -6.70550860828e-07
Gc1_61 0 n2 ns61 0 -1.59604541563e-06
Gc1_62 0 n2 ns62 0 4.38427267323e-07
Gc1_63 0 n2 ns63 0 -2.49472249676e-07
Gc1_64 0 n2 ns64 0 -3.31086261474e-07
Gc1_65 0 n2 ns65 0 5.10187713518e-07
Gc1_66 0 n2 ns66 0 5.26057012904e-09
Gc1_67 0 n2 ns67 0 6.29743488325e-08
Gc1_68 0 n2 ns68 0 -2.93206361134e-07
Gc1_69 0 n2 ns69 0 -2.77246705676e-07
Gc1_70 0 n2 ns70 0 5.26181318434e-07
Gc1_71 0 n2 ns71 0 -4.56625062905e-09
Gc1_72 0 n2 ns72 0 -1.91908117475e-09
Gc1_73 0 n2 ns73 0 0.000255627852429
Gc1_74 0 n2 ns74 0 -6.42873416842e-06
Gc1_75 0 n2 ns75 0 1.23217762639e-05
Gc1_76 0 n2 ns76 0 2.02328290635e-06
Gc1_77 0 n2 ns77 0 -0.000111142392723
Gc1_78 0 n2 ns78 0 -8.6404752839e-05
Gc1_79 0 n2 ns79 0 3.3281281639e-06
Gc1_80 0 n2 ns80 0 3.28649442325e-07
Gc1_81 0 n2 ns81 0 -0.000193365998062
Gc1_82 0 n2 ns82 0 4.30579104473e-06
Gc1_83 0 n2 ns83 0 -2.71300115619e-05
Gc1_84 0 n2 ns84 0 -5.13233030284e-05
Gc1_85 0 n2 ns85 0 -5.19808613777e-05
Gc1_86 0 n2 ns86 0 -1.02447817267e-05
Gc1_87 0 n2 ns87 0 -7.07990052351e-06
Gc1_88 0 n2 ns88 0 -1.68316835908e-05
Gc1_89 0 n2 ns89 0 7.63131403312e-05
Gc1_90 0 n2 ns90 0 -1.40056905352e-06
Gc1_91 0 n2 ns91 0 1.0545317299e-05
Gc1_92 0 n2 ns92 0 6.49273343603e-06
Gc1_93 0 n2 ns93 0 4.21332579687e-06
Gc1_94 0 n2 ns94 0 7.20418779089e-06
Gc1_95 0 n2 ns95 0 2.02985677331e-06
Gc1_96 0 n2 ns96 0 5.6811216195e-06
Gc1_97 0 n2 ns97 0 -3.20265433397e-06
Gc1_98 0 n2 ns98 0 1.01729570115e-07
Gc1_99 0 n2 ns99 0 -1.13660528189e-07
Gc1_100 0 n2 ns100 0 -5.15790751499e-06
Gc1_101 0 n2 ns101 0 -6.28834330417e-06
Gc1_102 0 n2 ns102 0 -1.50893624818e-07
Gc1_103 0 n2 ns103 0 -4.67872151664e-07
Gc1_104 0 n2 ns104 0 -1.57725381117e-07
Gc1_105 0 n2 ns105 0 -1.61502683143e-05
Gc1_106 0 n2 ns106 0 3.42125010003e-07
Gc1_107 0 n2 ns107 0 -1.95785849689e-06
Gc1_108 0 n2 ns108 0 -4.58958248434e-06
Gc1_109 0 n2 ns109 0 -6.11549326171e-06
Gc1_110 0 n2 ns110 0 -7.62966198547e-07
Gc1_111 0 n2 ns111 0 -8.29055558816e-07
Gc1_112 0 n2 ns112 0 -1.19183030654e-06
Gc1_113 0 n2 ns113 0 -3.87286364384e-06
Gc1_114 0 n2 ns114 0 8.98701049763e-08
Gc1_115 0 n2 ns115 0 -4.3163990464e-07
Gc1_116 0 n2 ns116 0 -1.50958242733e-06
Gc1_117 0 n2 ns117 0 -2.20913932122e-06
Gc1_118 0 n2 ns118 0 8.02495980396e-08
Gc1_119 0 n2 ns119 0 -2.61380148037e-07
Gc1_120 0 n2 ns120 0 -2.92972664086e-07
Gc1_121 0 n2 ns121 0 -4.57363747614e-07
Gc1_122 0 n2 ns122 0 2.31169762556e-08
Gc1_123 0 n2 ns123 0 -4.45258905153e-08
Gc1_124 0 n2 ns124 0 -3.66780861288e-07
Gc1_125 0 n2 ns125 0 -6.7277140007e-07
Gc1_126 0 n2 ns126 0 4.58997778174e-07
Gc1_127 0 n2 ns127 0 -7.27149246216e-08
Gc1_128 0 n2 ns128 0 -6.5843443029e-08
Gd1_1 0 n2 ni1 0 -0.00381103241716
Gd1_2 0 n2 ni2 0 0.00221362745707
Gd1_3 0 n2 ni3 0 0.000757511167204
Gd1_4 0 n2 ni4 0 1.04371483175e-05
Gd1_5 0 n2 ni5 0 -8.10531801031e-06
Gd1_6 0 n2 ni6 0 2.51435809681e-05
Gd1_7 0 n2 ni7 0 1.25802383049e-05
Gd1_8 0 n2 ni8 0 3.78622145149e-06
Gd1_9 0 n2 ni9 0 7.03349055232e-08
Gd1_10 0 n2 ni10 0 0.000191911773795
Gd1_11 0 n2 ni11 0 0.00023448060264
Gd1_12 0 n2 ni12 0 -7.20545335786e-05
Gd1_13 0 n2 ni13 0 3.92471066114e-06
Gd1_14 0 n2 ni14 0 1.57662550726e-05
Gd1_15 0 n2 ni15 0 3.85756382057e-06
Gd1_16 0 n2 ni16 0 7.68098493696e-07
Gc2_1 0 n4 ns1 0 0.00170344945102
Gc2_2 0 n4 ns2 0 -2.7551388872e-05
Gc2_3 0 n4 ns3 0 -4.37654841208e-06
Gc2_4 0 n4 ns4 0 0.000271099227809
Gc2_5 0 n4 ns5 0 -1.63421590459e-05
Gc2_6 0 n4 ns6 0 -0.000120082274237
Gc2_7 0 n4 ns7 0 9.55288533273e-05
Gc2_8 0 n4 ns8 0 -8.89608401891e-05
Gc2_9 0 n4 ns9 0 0.00260069059754
Gc2_10 0 n4 ns10 0 -4.47030416596e-05
Gc2_11 0 n4 ns11 0 0.000269322332498
Gc2_12 0 n4 ns12 0 0.000579768132752
Gc2_13 0 n4 ns13 0 0.000141976282936
Gc2_14 0 n4 ns14 0 -8.62561773966e-05
Gc2_15 0 n4 ns15 0 -5.24522154865e-05
Gc2_16 0 n4 ns16 0 0.000385843976967
Gc2_17 0 n4 ns17 0 0.000122412402595
Gc2_18 0 n4 ns18 0 -2.95107049888e-06
Gc2_19 0 n4 ns19 0 -6.57063608794e-06
Gc2_20 0 n4 ns20 0 -1.32783068216e-05
Gc2_21 0 n4 ns21 0 -8.66364038405e-05
Gc2_22 0 n4 ns22 0 -6.44744477251e-05
Gc2_23 0 n4 ns23 0 3.70709367749e-06
Gc2_24 0 n4 ns24 0 -1.30379249287e-05
Gc2_25 0 n4 ns25 0 -0.0001769890814
Gc2_26 0 n4 ns26 0 3.86264013441e-06
Gc2_27 0 n4 ns27 0 -2.48379927636e-05
Gc2_28 0 n4 ns28 0 -4.88702866317e-05
Gc2_29 0 n4 ns29 0 -4.94357623498e-05
Gc2_30 0 n4 ns30 0 -1.30485639412e-05
Gc2_31 0 n4 ns31 0 -6.63418616448e-06
Gc2_32 0 n4 ns32 0 -1.48935406905e-05
Gc2_33 0 n4 ns33 0 3.99528001588e-05
Gc2_34 0 n4 ns34 0 -6.26679121221e-07
Gc2_35 0 n4 ns35 0 5.33199386441e-06
Gc2_36 0 n4 ns36 0 3.11141579631e-06
Gc2_37 0 n4 ns37 0 1.98244796347e-06
Gc2_38 0 n4 ns38 0 6.546770846e-06
Gc2_39 0 n4 ns39 0 1.02194771538e-06
Gc2_40 0 n4 ns40 0 2.66323791257e-06
Gc2_41 0 n4 ns41 0 -5.87851167022e-06
Gc2_42 0 n4 ns42 0 1.66872821775e-07
Gc2_43 0 n4 ns43 0 -6.18210754769e-07
Gc2_44 0 n4 ns44 0 -4.87381382673e-06
Gc2_45 0 n4 ns45 0 -4.97813371834e-06
Gc2_46 0 n4 ns46 0 -8.00957143498e-09
Gc2_47 0 n4 ns47 0 -4.23845974177e-07
Gc2_48 0 n4 ns48 0 -4.02718130643e-07
Gc2_49 0 n4 ns49 0 -1.43956027769e-05
Gc2_50 0 n4 ns50 0 3.07874694091e-07
Gc2_51 0 n4 ns51 0 -1.77502818613e-06
Gc2_52 0 n4 ns52 0 -4.1324000856e-06
Gc2_53 0 n4 ns53 0 -5.13919841725e-06
Gc2_54 0 n4 ns54 0 -6.7150129803e-07
Gc2_55 0 n4 ns55 0 -7.04269457944e-07
Gc2_56 0 n4 ns56 0 -1.06363861359e-06
Gc2_57 0 n4 ns57 0 -5.92132847777e-06
Gc2_58 0 n4 ns58 0 1.33479806124e-07
Gc2_59 0 n4 ns59 0 -7.19054638995e-07
Gc2_60 0 n4 ns60 0 -1.18706051592e-06
Gc2_61 0 n4 ns61 0 -2.33458023821e-06
Gc2_62 0 n4 ns62 0 2.06921765449e-07
Gc2_63 0 n4 ns63 0 -3.57348366654e-07
Gc2_64 0 n4 ns64 0 -4.71494958902e-07
Gc2_65 0 n4 ns65 0 -1.69854637436e-06
Gc2_66 0 n4 ns66 0 4.8167449143e-08
Gc2_67 0 n4 ns67 0 -1.92968863617e-07
Gc2_68 0 n4 ns68 0 -2.43468214806e-07
Gc2_69 0 n4 ns69 0 -1.05675369117e-06
Gc2_70 0 n4 ns70 0 5.24336706599e-07
Gc2_71 0 n4 ns71 0 -1.60597604508e-07
Gc2_72 0 n4 ns72 0 -1.67112279397e-07
Gc2_73 0 n4 ns73 0 0.00200724653791
Gc2_74 0 n4 ns74 0 -3.91419194742e-05
Gc2_75 0 n4 ns75 0 0.000172003051018
Gc2_76 0 n4 ns76 0 0.000506691300361
Gc2_77 0 n4 ns77 0 2.3999336226e-05
Gc2_78 0 n4 ns78 0 -1.98679104574e-05
Gc2_79 0 n4 ns79 0 3.49336170623e-05
Gc2_80 0 n4 ns80 0 9.69560154653e-05
Gc2_81 0 n4 ns81 0 -0.000252088360404
Gc2_82 0 n4 ns82 0 4.93715114592e-06
Gc2_83 0 n4 ns83 0 -3.70945505007e-05
Gc2_84 0 n4 ns84 0 -7.48361684392e-05
Gc2_85 0 n4 ns85 0 -9.53200089991e-05
Gc2_86 0 n4 ns86 0 -4.33828894287e-05
Gc2_87 0 n4 ns87 0 -1.10705058984e-05
Gc2_88 0 n4 ns88 0 -2.13691782657e-05
Gc2_89 0 n4 ns89 0 3.93712811119e-05
Gc2_90 0 n4 ns90 0 -6.35542271504e-07
Gc2_91 0 n4 ns91 0 5.44236055417e-06
Gc2_92 0 n4 ns92 0 -5.25514533149e-06
Gc2_93 0 n4 ns93 0 -5.4450295489e-06
Gc2_94 0 n4 ns94 0 2.39747494239e-06
Gc2_95 0 n4 ns95 0 7.29437069202e-07
Gc2_96 0 n4 ns96 0 3.03402833101e-06
Gc2_97 0 n4 ns97 0 3.07376504922e-05
Gc2_98 0 n4 ns98 0 -5.61900590216e-07
Gc2_99 0 n4 ns99 0 4.42595244919e-06
Gc2_100 0 n4 ns100 0 4.81790138288e-07
Gc2_101 0 n4 ns101 0 -8.57540513525e-07
Gc2_102 0 n4 ns102 0 2.45427058053e-06
Gc2_103 0 n4 ns103 0 6.28826906924e-07
Gc2_104 0 n4 ns104 0 2.46635985147e-06
Gc2_105 0 n4 ns105 0 -1.19920105989e-05
Gc2_106 0 n4 ns106 0 2.61321680393e-07
Gc2_107 0 n4 ns107 0 -1.41279687907e-06
Gc2_108 0 n4 ns108 0 -5.16645518409e-06
Gc2_109 0 n4 ns109 0 -5.55650341292e-06
Gc2_110 0 n4 ns110 0 -9.49498283206e-07
Gc2_111 0 n4 ns111 0 -6.23081541388e-07
Gc2_112 0 n4 ns112 0 -8.14458859871e-07
Gc2_113 0 n4 ns113 0 -6.19618196583e-06
Gc2_114 0 n4 ns114 0 1.34841100182e-07
Gc2_115 0 n4 ns115 0 -7.18391090887e-07
Gc2_116 0 n4 ns116 0 -2.45395147122e-06
Gc2_117 0 n4 ns117 0 -2.96452147234e-06
Gc2_118 0 n4 ns118 0 -3.22964885518e-07
Gc2_119 0 n4 ns119 0 -3.47571912745e-07
Gc2_120 0 n4 ns120 0 -4.3294432116e-07
Gc2_121 0 n4 ns121 0 -2.51080993226e-06
Gc2_122 0 n4 ns122 0 6.2873687703e-08
Gc2_123 0 n4 ns123 0 -2.83810068169e-07
Gc2_124 0 n4 ns124 0 -4.83521858314e-07
Gc2_125 0 n4 ns125 0 -1.4035843426e-06
Gc2_126 0 n4 ns126 0 3.89496879272e-07
Gc2_127 0 n4 ns127 0 -2.07335119414e-07
Gc2_128 0 n4 ns128 0 -2.12477278762e-07
Gd2_1 0 n4 ni1 0 0.00221362745707
Gd2_2 0 n4 ni2 0 -0.00118212441964
Gd2_3 0 n4 ni3 0 0.000315917309198
Gd2_4 0 n4 ni4 0 0.000216076688167
Gd2_5 0 n4 ni5 0 -3.37144605455e-05
Gd2_6 0 n4 ni6 0 7.60703473324e-06
Gd2_7 0 n4 ni7 0 1.43812698675e-05
Gd2_8 0 n4 ni8 0 5.68761425467e-06
Gd2_9 0 n4 ni9 0 1.67449036216e-06
Gd2_10 0 n4 ni10 0 -0.000349284122458
Gd2_11 0 n4 ni11 0 0.000347779628347
Gd2_12 0 n4 ni12 0 -2.82324269034e-05
Gd2_13 0 n4 ni13 0 -2.93691804214e-05
Gd2_14 0 n4 ni14 0 1.24984800771e-05
Gd2_15 0 n4 ni15 0 6.23069991758e-06
Gd2_16 0 n4 ni16 0 2.35642833709e-06
Gc3_1 0 n6 ns1 0 -0.00059012372801
Gc3_2 0 n6 ns2 0 1.25618860156e-05
Gc3_3 0 n6 ns3 0 -8.71731718617e-05
Gc3_4 0 n6 ns4 0 -0.000146208400641
Gc3_5 0 n6 ns5 0 -0.000127315799585
Gc3_6 0 n6 ns6 0 -4.84194511262e-05
Gc3_7 0 n6 ns7 0 -1.67327972321e-05
Gc3_8 0 n6 ns8 0 -5.48870170322e-05
Gc3_9 0 n6 ns9 0 0.000122412402595
Gc3_10 0 n6 ns10 0 -2.95107049888e-06
Gc3_11 0 n6 ns11 0 -6.57063608794e-06
Gc3_12 0 n6 ns12 0 -1.32783068216e-05
Gc3_13 0 n6 ns13 0 -8.66364038405e-05
Gc3_14 0 n6 ns14 0 -6.44744477251e-05
Gc3_15 0 n6 ns15 0 3.70709367749e-06
Gc3_16 0 n6 ns16 0 -1.30379249287e-05
Gc3_17 0 n6 ns17 0 0.00251905080759
Gc3_18 0 n6 ns18 0 -4.30604082668e-05
Gc3_19 0 n6 ns19 0 0.000271677910728
Gc3_20 0 n6 ns20 0 0.000594928207119
Gc3_21 0 n6 ns21 0 0.00014707668778
Gc3_22 0 n6 ns22 0 -6.92591515693e-05
Gc3_23 0 n6 ns23 0 -6.34976044128e-05
Gc3_24 0 n6 ns24 0 0.000399939082929
Gc3_25 0 n6 ns25 0 0.000279634092761
Gc3_26 0 n6 ns26 0 -6.48976219973e-06
Gc3_27 0 n6 ns27 0 1.56566215486e-05
Gc3_28 0 n6 ns28 0 1.532421475e-05
Gc3_29 0 n6 ns29 0 -7.12432987436e-05
Gc3_30 0 n6 ns30 0 -6.47325068318e-05
Gc3_31 0 n6 ns31 0 7.25159927378e-06
Gc3_32 0 n6 ns32 0 1.3190210159e-06
Gc3_33 0 n6 ns33 0 -0.000243981691387
Gc3_34 0 n6 ns34 0 5.45955876037e-06
Gc3_35 0 n6 ns35 0 -3.46841541441e-05
Gc3_36 0 n6 ns36 0 -5.60766663964e-05
Gc3_37 0 n6 ns37 0 -4.87489289226e-05
Gc3_38 0 n6 ns38 0 -9.12308526774e-06
Gc3_39 0 n6 ns39 0 -7.86672946601e-06
Gc3_40 0 n6 ns40 0 -2.10525569138e-05
Gc3_41 0 n6 ns41 0 4.96728515638e-05
Gc3_42 0 n6 ns42 0 -8.24559214036e-07
Gc3_43 0 n6 ns43 0 6.51862176208e-06
Gc3_44 0 n6 ns44 0 2.67618678468e-06
Gc3_45 0 n6 ns45 0 4.92694351455e-06
Gc3_46 0 n6 ns46 0 6.1317161694e-06
Gc3_47 0 n6 ns47 0 1.637804931e-06
Gc3_48 0 n6 ns48 0 3.5120663778e-06
Gc3_49 0 n6 ns49 0 4.59036299543e-07
Gc3_50 0 n6 ns50 0 4.08272732409e-08
Gc3_51 0 n6 ns51 0 1.15919400617e-07
Gc3_52 0 n6 ns52 0 -5.11515573862e-06
Gc3_53 0 n6 ns53 0 -2.70796449419e-06
Gc3_54 0 n6 ns54 0 -1.89877957179e-07
Gc3_55 0 n6 ns55 0 3.38233236775e-08
Gc3_56 0 n6 ns56 0 9.13761507797e-08
Gc3_57 0 n6 ns57 0 -1.19625816287e-05
Gc3_58 0 n6 ns58 0 2.62646452171e-07
Gc3_59 0 n6 ns59 0 -1.52906907275e-06
Gc3_60 0 n6 ns60 0 -4.34176643557e-06
Gc3_61 0 n6 ns61 0 -3.90455962093e-06
Gc3_62 0 n6 ns62 0 -7.43265055281e-07
Gc3_63 0 n6 ns63 0 -4.77460262438e-07
Gc3_64 0 n6 ns64 0 -8.86443564675e-07
Gc3_65 0 n6 ns65 0 -5.38569718614e-06
Gc3_66 0 n6 ns66 0 1.20928343182e-07
Gc3_67 0 n6 ns67 0 -6.19617568441e-07
Gc3_68 0 n6 ns68 0 -1.42170536585e-06
Gc3_69 0 n6 ns69 0 -2.61192606132e-06
Gc3_70 0 n6 ns70 0 1.45873987595e-07
Gc3_71 0 n6 ns71 0 -3.55447237246e-07
Gc3_72 0 n6 ns72 0 -4.19395235924e-07
Gc3_73 0 n6 ns73 0 0.00146919185322
Gc3_74 0 n6 ns74 0 -2.12857910264e-05
Gc3_75 0 n6 ns75 0 -4.2977754716e-05
Gc3_76 0 n6 ns76 0 0.000246698064878
Gc3_77 0 n6 ns77 0 1.24625551942e-06
Gc3_78 0 n6 ns78 0 -9.54218550464e-05
Gc3_79 0 n6 ns79 0 9.24107291793e-05
Gc3_80 0 n6 ns80 0 -0.000112217613401
Gc3_81 0 n6 ns81 0 0.0017314763145
Gc3_82 0 n6 ns82 0 -3.29028759871e-05
Gc3_83 0 n6 ns83 0 0.00012794972743
Gc3_84 0 n6 ns84 0 0.000424052302862
Gc3_85 0 n6 ns85 0 1.94550881083e-05
Gc3_86 0 n6 ns86 0 -2.65260469772e-05
Gc3_87 0 n6 ns87 0 3.83172714771e-05
Gc3_88 0 n6 ns88 0 6.11434746033e-05
Gc3_89 0 n6 ns89 0 -0.000190010036797
Gc3_90 0 n6 ns90 0 3.49364153638e-06
Gc3_91 0 n6 ns91 0 -2.83968096019e-05
Gc3_92 0 n6 ns92 0 -6.85762365233e-05
Gc3_93 0 n6 ns93 0 -8.98826290617e-05
Gc3_94 0 n6 ns94 0 -4.70144525347e-05
Gc3_95 0 n6 ns95 0 -9.36190505878e-06
Gc3_96 0 n6 ns96 0 -1.54310405027e-05
Gc3_97 0 n6 ns97 0 2.82408980511e-05
Gc3_98 0 n6 ns98 0 -3.7441614715e-07
Gc3_99 0 n6 ns99 0 3.67738043991e-06
Gc3_100 0 n6 ns100 0 -6.85504679692e-06
Gc3_101 0 n6 ns101 0 -4.24614979483e-06
Gc3_102 0 n6 ns102 0 2.56667383025e-06
Gc3_103 0 n6 ns103 0 6.93161381618e-07
Gc3_104 0 n6 ns104 0 1.99197980264e-06
Gc3_105 0 n6 ns105 0 2.80279685742e-05
Gc3_106 0 n6 ns106 0 -4.93144821695e-07
Gc3_107 0 n6 ns107 0 3.83671043534e-06
Gc3_108 0 n6 ns108 0 -1.36289478433e-06
Gc3_109 0 n6 ns109 0 9.09554492912e-07
Gc3_110 0 n6 ns110 0 1.84427314005e-06
Gc3_111 0 n6 ns111 0 8.92518168504e-07
Gc3_112 0 n6 ns112 0 2.23198932125e-06
Gc3_113 0 n6 ns113 0 -6.24111369122e-06
Gc3_114 0 n6 ns114 0 1.4587871265e-07
Gc3_115 0 n6 ns115 0 -7.41931778459e-07
Gc3_116 0 n6 ns116 0 -5.71700638605e-06
Gc3_117 0 n6 ns117 0 -3.55787956916e-06
Gc3_118 0 n6 ns118 0 -1.26140224618e-06
Gc3_119 0 n6 ns119 0 -1.92929668152e-07
Gc3_120 0 n6 ns120 0 -3.46911814172e-07
Gc3_121 0 n6 ns121 0 -6.61507577058e-06
Gc3_122 0 n6 ns122 0 1.44858704987e-07
Gc3_123 0 n6 ns123 0 -7.81728229064e-07
Gc3_124 0 n6 ns124 0 -2.43268002078e-06
Gc3_125 0 n6 ns125 0 -2.96651042326e-06
Gc3_126 0 n6 ns126 0 -2.80914841197e-07
Gc3_127 0 n6 ns127 0 -3.61299282375e-07
Gc3_128 0 n6 ns128 0 -4.72741089205e-07
Gd3_1 0 n6 ni1 0 0.000757511167204
Gd3_2 0 n6 ni2 0 0.000315917309198
Gd3_3 0 n6 ni3 0 -0.00133534297282
Gd3_4 0 n6 ni4 0 0.000144002881421
Gd3_5 0 n6 ni5 0 0.000289381320077
Gd3_6 0 n6 ni6 0 -4.14097054281e-05
Gd3_7 0 n6 ni7 0 3.01232302647e-06
Gd3_8 0 n6 ni8 0 1.3045771699e-05
Gd3_9 0 n6 ni9 0 5.06716986895e-06
Gd3_10 0 n6 ni10 0 0.00253137732265
Gd3_11 0 n6 ni11 0 3.42237858476e-05
Gd3_12 0 n6 ni12 0 0.000283446559501
Gd3_13 0 n6 ni13 0 -1.45015742586e-05
Gd3_14 0 n6 ni14 0 -2.36829738593e-05
Gd3_15 0 n6 ni15 0 8.43232800288e-06
Gd3_16 0 n6 ni16 0 6.69100849414e-06
Gc4_1 0 n8 ns1 0 6.19520587657e-06
Gc4_2 0 n8 ns2 0 2.3784522811e-07
Gc4_3 0 n8 ns3 0 4.43393574485e-07
Gc4_4 0 n8 ns4 0 -5.71073410869e-06
Gc4_5 0 n8 ns5 0 -7.17293235846e-06
Gc4_6 0 n8 ns6 0 8.20625932242e-06
Gc4_7 0 n8 ns7 0 -1.44159389408e-07
Gc4_8 0 n8 ns8 0 -8.97282516464e-07
Gc4_9 0 n8 ns9 0 -0.0001769890814
Gc4_10 0 n8 ns10 0 3.86264013441e-06
Gc4_11 0 n8 ns11 0 -2.48379927635e-05
Gc4_12 0 n8 ns12 0 -4.88702866317e-05
Gc4_13 0 n8 ns13 0 -4.94357623498e-05
Gc4_14 0 n8 ns14 0 -1.30485639412e-05
Gc4_15 0 n8 ns15 0 -6.63418616448e-06
Gc4_16 0 n8 ns16 0 -1.48935406905e-05
Gc4_17 0 n8 ns17 0 0.000279634092761
Gc4_18 0 n8 ns18 0 -6.48976219973e-06
Gc4_19 0 n8 ns19 0 1.56566215486e-05
Gc4_20 0 n8 ns20 0 1.532421475e-05
Gc4_21 0 n8 ns21 0 -7.12432987436e-05
Gc4_22 0 n8 ns22 0 -6.47325068318e-05
Gc4_23 0 n8 ns23 0 7.25159927378e-06
Gc4_24 0 n8 ns24 0 1.3190210159e-06
Gc4_25 0 n8 ns25 0 0.00260067351357
Gc4_26 0 n8 ns26 0 -4.43719147818e-05
Gc4_27 0 n8 ns27 0 0.000264825364094
Gc4_28 0 n8 ns28 0 0.000566471566705
Gc4_29 0 n8 ns29 0 0.000160267196087
Gc4_30 0 n8 ns30 0 -8.62548657242e-05
Gc4_31 0 n8 ns31 0 -4.8023306723e-05
Gc4_32 0 n8 ns32 0 0.000381388984162
Gc4_33 0 n8 ns33 0 -4.07948267591e-05
Gc4_34 0 n8 ns34 0 9.31279645013e-07
Gc4_35 0 n8 ns35 0 -3.32638008652e-05
Gc4_36 0 n8 ns36 0 -5.163337651e-05
Gc4_37 0 n8 ns37 0 -8.82407690562e-05
Gc4_38 0 n8 ns38 0 -6.48347931539e-05
Gc4_39 0 n8 ns39 0 3.57856040065e-06
Gc4_40 0 n8 ns40 0 -3.17977602097e-05
Gc4_41 0 n8 ns41 0 -0.000206485326768
Gc4_42 0 n8 ns42 0 4.60971571495e-06
Gc4_43 0 n8 ns43 0 -2.94298226141e-05
Gc4_44 0 n8 ns44 0 -5.09703183045e-05
Gc4_45 0 n8 ns45 0 -4.60828786203e-05
Gc4_46 0 n8 ns46 0 -9.95306725945e-06
Gc4_47 0 n8 ns47 0 -6.92366866195e-06
Gc4_48 0 n8 ns48 0 -1.77704474297e-05
Gc4_49 0 n8 ns49 0 4.3280521616e-05
Gc4_50 0 n8 ns50 0 -6.98886134231e-07
Gc4_51 0 n8 ns51 0 5.65606584615e-06
Gc4_52 0 n8 ns52 0 1.37652488969e-06
Gc4_53 0 n8 ns53 0 3.73145319615e-06
Gc4_54 0 n8 ns54 0 5.55296473603e-06
Gc4_55 0 n8 ns55 0 1.43839252755e-06
Gc4_56 0 n8 ns56 0 2.99980129396e-06
Gc4_57 0 n8 ns57 0 -6.79808647133e-06
Gc4_58 0 n8 ns58 0 1.93351006335e-07
Gc4_59 0 n8 ns59 0 -8.43279871695e-07
Gc4_60 0 n8 ns60 0 -5.14154465606e-06
Gc4_61 0 n8 ns61 0 -4.11077977791e-06
Gc4_62 0 n8 ns62 0 -1.50817841073e-08
Gc4_63 0 n8 ns63 0 -3.21519209221e-07
Gc4_64 0 n8 ns64 0 -5.24812425234e-07
Gc4_65 0 n8 ns65 0 -1.74728450152e-05
Gc4_66 0 n8 ns66 0 3.67151640903e-07
Gc4_67 0 n8 ns67 0 -2.09229230608e-06
Gc4_68 0 n8 ns68 0 -4.2837217456e-06
Gc4_69 0 n8 ns69 0 -6.77155368265e-06
Gc4_70 0 n8 ns70 0 -6.34773702603e-07
Gc4_71 0 n8 ns71 0 -9.60648440033e-07
Gc4_72 0 n8 ns72 0 -1.30456977862e-06
Gc4_73 0 n8 ns73 0 -0.000528989617471
Gc4_74 0 n8 ns74 0 1.12284364269e-05
Gc4_75 0 n8 ns75 0 -7.89151534504e-05
Gc4_76 0 n8 ns76 0 -0.00012915155275
Gc4_77 0 n8 ns77 0 -0.000113282011914
Gc4_78 0 n8 ns78 0 -4.54158863742e-05
Gc4_79 0 n8 ns79 0 -1.49383207297e-05
Gc4_80 0 n8 ns80 0 -4.94848425366e-05
Gc4_81 0 n8 ns81 0 0.00168679657982
Gc4_82 0 n8 ns82 0 -2.68448755633e-05
Gc4_83 0 n8 ns83 0 8.02085238536e-06
Gc4_84 0 n8 ns84 0 0.000337410115542
Gc4_85 0 n8 ns85 0 1.13479066436e-05
Gc4_86 0 n8 ns86 0 -7.58389803008e-05
Gc4_87 0 n8 ns87 0 8.25271002342e-05
Gc4_88 0 n8 ns88 0 -6.61406514889e-05
Gc4_89 0 n8 ns89 0 0.00174050680003
Gc4_90 0 n8 ns90 0 -3.32490526527e-05
Gc4_91 0 n8 ns91 0 0.000133089643448
Gc4_92 0 n8 ns92 0 0.0004330019464
Gc4_93 0 n8 ns93 0 1.83869460392e-05
Gc4_94 0 n8 ns94 0 -2.46137986848e-05
Gc4_95 0 n8 ns95 0 3.57447983553e-05
Gc4_96 0 n8 ns96 0 6.74656402172e-05
Gc4_97 0 n8 ns97 0 -0.000225357024387
Gc4_98 0 n8 ns98 0 4.37159219207e-06
Gc4_99 0 n8 ns99 0 -3.37666355749e-05
Gc4_100 0 n8 ns100 0 -7.20047533642e-05
Gc4_101 0 n8 ns101 0 -8.81755207605e-05
Gc4_102 0 n8 ns102 0 -4.33214105264e-05
Gc4_103 0 n8 ns103 0 -9.6701621047e-06
Gc4_104 0 n8 ns104 0 -1.93393953924e-05
Gc4_105 0 n8 ns105 0 1.78065239761e-05
Gc4_106 0 n8 ns106 0 -1.25395336539e-07
Gc4_107 0 n8 ns107 0 2.05102572646e-06
Gc4_108 0 n8 ns108 0 -7.4312727416e-06
Gc4_109 0 n8 ns109 0 -3.66998409759e-06
Gc4_110 0 n8 ns110 0 3.18402644594e-06
Gc4_111 0 n8 ns111 0 5.12260365718e-07
Gc4_112 0 n8 ns112 0 1.01091470225e-06
Gc4_113 0 n8 ns113 0 3.03775569146e-05
Gc4_114 0 n8 ns114 0 -5.44309186014e-07
Gc4_115 0 n8 ns115 0 4.19204876073e-06
Gc4_116 0 n8 ns116 0 -8.76958685759e-07
Gc4_117 0 n8 ns117 0 9.41694995034e-07
Gc4_118 0 n8 ns118 0 1.97596118906e-06
Gc4_119 0 n8 ns119 0 9.24058503081e-07
Gc4_120 0 n8 ns120 0 2.4279042646e-06
Gc4_121 0 n8 ns121 0 -1.33757747242e-05
Gc4_122 0 n8 ns122 0 2.90673759896e-07
Gc4_123 0 n8 ns123 0 -1.58852394086e-06
Gc4_124 0 n8 ns124 0 -5.104172281e-06
Gc4_125 0 n8 ns125 0 -5.90425640655e-06
Gc4_126 0 n8 ns126 0 -8.75761924157e-07
Gc4_127 0 n8 ns127 0 -7.06633272464e-07
Gc4_128 0 n8 ns128 0 -9.30544897281e-07
Gd4_1 0 n8 ni1 0 1.04371483175e-05
Gd4_2 0 n8 ni2 0 0.000216076688167
Gd4_3 0 n8 ni3 0 0.000144002881421
Gd4_4 0 n8 ni4 0 -0.00111345938045
Gd4_5 0 n8 ni5 0 0.000548549085442
Gd4_6 0 n8 ni6 0 0.000250444533447
Gd4_7 0 n8 ni7 0 -3.4805545205e-05
Gd4_8 0 n8 ni8 0 9.63805909615e-06
Gd4_9 0 n8 ni9 0 1.64120887921e-05
Gd4_10 0 n8 ni10 0 0.000689640310647
Gd4_11 0 n8 ni11 0 0.00195227228226
Gd4_12 0 n8 ni12 0 -3.99250798225e-05
Gd4_13 0 n8 ni13 0 0.000324198017446
Gd4_14 0 n8 ni14 0 -2.14075632551e-06
Gd4_15 0 n8 ni15 0 -2.65146579729e-05
Gd4_16 0 n8 ni16 0 1.36673536186e-05
Gc5_1 0 n10 ns1 0 1.20370228915e-05
Gc5_2 0 n10 ns2 0 -1.22155562566e-07
Gc5_3 0 n10 ns3 0 1.70327311833e-06
Gc5_4 0 n10 ns4 0 -1.59210198577e-06
Gc5_5 0 n10 ns5 0 -2.74622201324e-06
Gc5_6 0 n10 ns6 0 3.41159763809e-06
Gc5_7 0 n10 ns7 0 1.06493496518e-07
Gc5_8 0 n10 ns8 0 6.31246642884e-07
Gc5_9 0 n10 ns9 0 3.99528001588e-05
Gc5_10 0 n10 ns10 0 -6.26679121221e-07
Gc5_11 0 n10 ns11 0 5.33199386441e-06
Gc5_12 0 n10 ns12 0 3.11141579631e-06
Gc5_13 0 n10 ns13 0 1.98244796347e-06
Gc5_14 0 n10 ns14 0 6.546770846e-06
Gc5_15 0 n10 ns15 0 1.02194771538e-06
Gc5_16 0 n10 ns16 0 2.66323791257e-06
Gc5_17 0 n10 ns17 0 -0.000243981691387
Gc5_18 0 n10 ns18 0 5.45955876037e-06
Gc5_19 0 n10 ns19 0 -3.46841541441e-05
Gc5_20 0 n10 ns20 0 -5.60766663964e-05
Gc5_21 0 n10 ns21 0 -4.87489289226e-05
Gc5_22 0 n10 ns22 0 -9.12308526774e-06
Gc5_23 0 n10 ns23 0 -7.86672946601e-06
Gc5_24 0 n10 ns24 0 -2.10525569138e-05
Gc5_25 0 n10 ns25 0 -4.0794826759e-05
Gc5_26 0 n10 ns26 0 9.31279645013e-07
Gc5_27 0 n10 ns27 0 -3.32638008652e-05
Gc5_28 0 n10 ns28 0 -5.163337651e-05
Gc5_29 0 n10 ns29 0 -8.82407690562e-05
Gc5_30 0 n10 ns30 0 -6.48347931539e-05
Gc5_31 0 n10 ns31 0 3.57856040065e-06
Gc5_32 0 n10 ns32 0 -3.17977602097e-05
Gc5_33 0 n10 ns33 0 0.00175013082332
Gc5_34 0 n10 ns34 0 -2.69569089188e-05
Gc5_35 0 n10 ns35 0 0.000193708702732
Gc5_36 0 n10 ns36 0 0.000557633004378
Gc5_37 0 n10 ns37 0 5.64627387586e-05
Gc5_38 0 n10 ns38 0 -3.65753770581e-05
Gc5_39 0 n10 ns39 0 -0.000105415606068
Gc5_40 0 n10 ns40 0 0.000370626805168
Gc5_41 0 n10 ns41 0 0.000412259160408
Gc5_42 0 n10 ns42 0 -9.48240577252e-06
Gc5_43 0 n10 ns43 0 3.33999673102e-05
Gc5_44 0 n10 ns44 0 3.78587860917e-05
Gc5_45 0 n10 ns45 0 -6.33930904236e-05
Gc5_46 0 n10 ns46 0 -6.75827939395e-05
Gc5_47 0 n10 ns47 0 1.02435553187e-05
Gc5_48 0 n10 ns48 0 1.22495099161e-05
Gc5_49 0 n10 ns49 0 -0.000185335650556
Gc5_50 0 n10 ns50 0 3.96983473583e-06
Gc5_51 0 n10 ns51 0 -2.59514998832e-05
Gc5_52 0 n10 ns52 0 -5.36050550876e-05
Gc5_53 0 n10 ns53 0 -5.19036319829e-05
Gc5_54 0 n10 ns54 0 -1.67076827822e-05
Gc5_55 0 n10 ns55 0 -6.74781351401e-06
Gc5_56 0 n10 ns56 0 -1.53385987311e-05
Gc5_57 0 n10 ns57 0 5.02184661993e-05
Gc5_58 0 n10 ns58 0 -8.49006009216e-07
Gc5_59 0 n10 ns59 0 6.75616558048e-06
Gc5_60 0 n10 ns60 0 3.45485942299e-06
Gc5_61 0 n10 ns61 0 3.43105159953e-06
Gc5_62 0 n10 ns62 0 6.30534242317e-06
Gc5_63 0 n10 ns63 0 1.44222411758e-06
Gc5_64 0 n10 ns64 0 3.55333625778e-06
Gc5_65 0 n10 ns65 0 2.35174293607e-06
Gc5_66 0 n10 ns66 0 -2.08109595048e-08
Gc5_67 0 n10 ns67 0 7.20481168481e-07
Gc5_68 0 n10 ns68 0 -4.07483878871e-06
Gc5_69 0 n10 ns69 0 -6.22805854561e-06
Gc5_70 0 n10 ns70 0 1.01369202911e-07
Gc5_71 0 n10 ns71 0 -3.80974860043e-07
Gc5_72 0 n10 ns72 0 2.89974094324e-07
Gc5_73 0 n10 ns73 0 -7.09137768122e-05
Gc5_74 0 n10 ns74 0 1.94024935126e-06
Gc5_75 0 n10 ns75 0 -1.06275646452e-05
Gc5_76 0 n10 ns76 0 -1.3552784779e-05
Gc5_77 0 n10 ns77 0 -1.02410512869e-05
Gc5_78 0 n10 ns78 0 8.57758204151e-06
Gc5_79 0 n10 ns79 0 -2.10086364247e-06
Gc5_80 0 n10 ns80 0 -7.35502662103e-06
Gc5_81 0 n10 ns81 0 -0.000583120781668
Gc5_82 0 n10 ns82 0 1.24796099228e-05
Gc5_83 0 n10 ns83 0 -8.69690055429e-05
Gc5_84 0 n10 ns84 0 -0.000140598714665
Gc5_85 0 n10 ns85 0 -0.000114830909271
Gc5_86 0 n10 ns86 0 -4.53618394728e-05
Gc5_87 0 n10 ns87 0 -1.55582568209e-05
Gc5_88 0 n10 ns88 0 -5.46568832722e-05
Gc5_89 0 n10 ns89 0 0.00203041538367
Gc5_90 0 n10 ns90 0 -3.29455410893e-05
Gc5_91 0 n10 ns91 0 8.31761413782e-06
Gc5_92 0 n10 ns92 0 0.000266181855967
Gc5_93 0 n10 ns93 0 7.56587628206e-05
Gc5_94 0 n10 ns94 0 -0.00011785218718
Gc5_95 0 n10 ns95 0 0.000129453843313
Gc5_96 0 n10 ns96 0 -0.00010318538896
Gc5_97 0 n10 ns97 0 0.00233822841415
Gc5_98 0 n10 ns98 0 -4.63278519359e-05
Gc5_99 0 n10 ns99 0 0.000214754458055
Gc5_100 0 n10 ns100 0 0.000544871474744
Gc5_101 0 n10 ns101 0 7.40170166462e-05
Gc5_102 0 n10 ns102 0 -1.94298070595e-05
Gc5_103 0 n10 ns103 0 4.90021007107e-05
Gc5_104 0 n10 ns104 0 0.00011947861877
Gc5_105 0 n10 ns105 0 -0.000203988445157
Gc5_106 0 n10 ns106 0 3.7940735961e-06
Gc5_107 0 n10 ns107 0 -3.0472158993e-05
Gc5_108 0 n10 ns108 0 -7.15652636847e-05
Gc5_109 0 n10 ns109 0 -9.12514232437e-05
Gc5_110 0 n10 ns110 0 -4.75841721521e-05
Gc5_111 0 n10 ns111 0 -9.55089307198e-06
Gc5_112 0 n10 ns112 0 -1.68764038398e-05
Gc5_113 0 n10 ns113 0 3.81124211666e-05
Gc5_114 0 n10 ns114 0 -6.06500104008e-07
Gc5_115 0 n10 ns115 0 5.21287235809e-06
Gc5_116 0 n10 ns116 0 -6.59245038961e-06
Gc5_117 0 n10 ns117 0 -4.56097985542e-06
Gc5_118 0 n10 ns118 0 1.95281954917e-06
Gc5_119 0 n10 ns119 0 8.9217208181e-07
Gc5_120 0 n10 ns120 0 2.96175337955e-06
Gc5_121 0 n10 ns121 0 3.36720091403e-05
Gc5_122 0 n10 ns122 0 -6.24253823121e-07
Gc5_123 0 n10 ns123 0 4.86138862183e-06
Gc5_124 0 n10 ns124 0 9.45181086767e-07
Gc5_125 0 n10 ns125 0 -7.84318096147e-07
Gc5_126 0 n10 ns126 0 2.58471141307e-06
Gc5_127 0 n10 ns127 0 6.76330586715e-07
Gc5_128 0 n10 ns128 0 2.72312753278e-06
Gd5_1 0 n10 ni1 0 -8.10531801031e-06
Gd5_2 0 n10 ni2 0 -3.37144605455e-05
Gd5_3 0 n10 ni3 0 0.000289381320077
Gd5_4 0 n10 ni4 0 0.000548549085442
Gd5_5 0 n10 ni5 0 -0.00102650589762
Gd5_6 0 n10 ni6 0 1.85714678132e-05
Gd5_7 0 n10 ni7 0 0.00022598784627
Gd5_8 0 n10 ni8 0 -4.40192767264e-05
Gd5_9 0 n10 ni9 0 -2.64877748396e-06
Gd5_10 0 n10 ni10 0 9.17481698985e-05
Gd5_11 0 n10 ni11 0 0.00075391676804
Gd5_12 0 n10 ni12 0 0.00239421290958
Gd5_13 0 n10 ni13 0 -0.000645710813608
Gd5_14 0 n10 ni14 0 0.000300400610231
Gd5_15 0 n10 ni15 0 -2.61303007592e-05
Gd5_16 0 n10 ni16 0 -3.27183378631e-05
Gc6_1 0 n12 ns1 0 -2.45215524068e-05
Gc6_2 0 n12 ns2 0 5.30778522145e-07
Gc6_3 0 n12 ns3 0 -3.08396167442e-06
Gc6_4 0 n12 ns4 0 -7.06056896579e-06
Gc6_5 0 n12 ns5 0 -8.13413540933e-06
Gc6_6 0 n12 ns6 0 -1.08609338201e-06
Gc6_7 0 n12 ns7 0 -1.11224817746e-06
Gc6_8 0 n12 ns8 0 -1.866996702e-06
Gc6_9 0 n12 ns9 0 -5.87851167022e-06
Gc6_10 0 n12 ns10 0 1.66872821775e-07
Gc6_11 0 n12 ns11 0 -6.18210754769e-07
Gc6_12 0 n12 ns12 0 -4.87381382673e-06
Gc6_13 0 n12 ns13 0 -4.97813371834e-06
Gc6_14 0 n12 ns14 0 -8.00957143502e-09
Gc6_15 0 n12 ns15 0 -4.23845974177e-07
Gc6_16 0 n12 ns16 0 -4.02718130643e-07
Gc6_17 0 n12 ns17 0 4.96728515638e-05
Gc6_18 0 n12 ns18 0 -8.24559214036e-07
Gc6_19 0 n12 ns19 0 6.51862176208e-06
Gc6_20 0 n12 ns20 0 2.67618678468e-06
Gc6_21 0 n12 ns21 0 4.92694351455e-06
Gc6_22 0 n12 ns22 0 6.1317161694e-06
Gc6_23 0 n12 ns23 0 1.637804931e-06
Gc6_24 0 n12 ns24 0 3.5120663778e-06
Gc6_25 0 n12 ns25 0 -0.000206485326768
Gc6_26 0 n12 ns26 0 4.60971571495e-06
Gc6_27 0 n12 ns27 0 -2.94298226141e-05
Gc6_28 0 n12 ns28 0 -5.09703183045e-05
Gc6_29 0 n12 ns29 0 -4.60828786203e-05
Gc6_30 0 n12 ns30 0 -9.95306725945e-06
Gc6_31 0 n12 ns31 0 -6.92366866195e-06
Gc6_32 0 n12 ns32 0 -1.77704474297e-05
Gc6_33 0 n12 ns33 0 0.000412259160408
Gc6_34 0 n12 ns34 0 -9.48240577252e-06
Gc6_35 0 n12 ns35 0 3.33999673102e-05
Gc6_36 0 n12 ns36 0 3.78587860917e-05
Gc6_37 0 n12 ns37 0 -6.33930904236e-05
Gc6_38 0 n12 ns38 0 -6.75827939395e-05
Gc6_39 0 n12 ns39 0 1.02435553187e-05
Gc6_40 0 n12 ns40 0 1.22495099161e-05
Gc6_41 0 n12 ns41 0 0.00265761189786
Gc6_42 0 n12 ns42 0 -4.57646122076e-05
Gc6_43 0 n12 ns43 0 0.000280457536726
Gc6_44 0 n12 ns44 0 0.000591784924693
Gc6_45 0 n12 ns45 0 0.000167355020856
Gc6_46 0 n12 ns46 0 -7.81141672533e-05
Gc6_47 0 n12 ns47 0 -5.21956918871e-05
Gc6_48 0 n12 ns48 0 0.000398136080107
Gc6_49 0 n12 ns49 0 0.000265667925407
Gc6_50 0 n12 ns50 0 -6.05006730401e-06
Gc6_51 0 n12 ns51 0 1.29188054699e-05
Gc6_52 0 n12 ns52 0 1.26795103389e-05
Gc6_53 0 n12 ns53 0 -6.41898569531e-05
Gc6_54 0 n12 ns54 0 -5.99813016744e-05
Gc6_55 0 n12 ns55 0 8.51129878975e-06
Gc6_56 0 n12 ns56 0 -1.87342241056e-06
Gc6_57 0 n12 ns57 0 -0.00020740116331
Gc6_58 0 n12 ns58 0 4.60119408212e-06
Gc6_59 0 n12 ns59 0 -2.94944542424e-05
Gc6_60 0 n12 ns60 0 -4.99524118779e-05
Gc6_61 0 n12 ns61 0 -4.74496175099e-05
Gc6_62 0 n12 ns62 0 -9.9856156687e-06
Gc6_63 0 n12 ns63 0 -7.04326277586e-06
Gc6_64 0 n12 ns64 0 -1.81008981411e-05
Gc6_65 0 n12 ns65 0 6.31549198078e-05
Gc6_66 0 n12 ns66 0 -1.13676191605e-06
Gc6_67 0 n12 ns67 0 8.72455823149e-06
Gc6_68 0 n12 ns68 0 4.21748439968e-06
Gc6_69 0 n12 ns69 0 2.16334025006e-06
Gc6_70 0 n12 ns70 0 6.34016736344e-06
Gc6_71 0 n12 ns71 0 1.66622588384e-06
Gc6_72 0 n12 ns72 0 4.52368549783e-06
Gc6_73 0 n12 ns73 0 1.22499948205e-05
Gc6_74 0 n12 ns74 0 -1.19278604293e-07
Gc6_75 0 n12 ns75 0 1.54394149213e-06
Gc6_76 0 n12 ns76 0 -1.45605242078e-06
Gc6_77 0 n12 ns77 0 -2.22156682214e-07
Gc6_78 0 n12 ns78 0 3.2872473059e-06
Gc6_79 0 n12 ns79 0 3.6405420909e-07
Gc6_80 0 n12 ns80 0 6.75091556278e-07
Gc6_81 0 n12 ns81 0 -2.78564405109e-05
Gc6_82 0 n12 ns82 0 9.40051105009e-07
Gc6_83 0 n12 ns83 0 -4.48509036758e-06
Gc6_84 0 n12 ns84 0 -1.11321965317e-05
Gc6_85 0 n12 ns85 0 -8.18315057366e-06
Gc6_86 0 n12 ns86 0 5.86589387302e-06
Gc6_87 0 n12 ns87 0 -8.57782587434e-07
Gc6_88 0 n12 ns88 0 -3.44105375606e-06
Gc6_89 0 n12 ns89 0 -0.000640052099338
Gc6_90 0 n12 ns90 0 1.38358711651e-05
Gc6_91 0 n12 ns91 0 -9.48126522045e-05
Gc6_92 0 n12 ns92 0 -0.000152983194766
Gc6_93 0 n12 ns93 0 -0.000114445239096
Gc6_94 0 n12 ns94 0 -4.37858698061e-05
Gc6_95 0 n12 ns95 0 -1.64589791744e-05
Gc6_96 0 n12 ns96 0 -5.8956597428e-05
Gc6_97 0 n12 ns97 0 0.00132828207303
Gc6_98 0 n12 ns98 0 -1.86033709536e-05
Gc6_99 0 n12 ns99 0 -5.03807738877e-05
Gc6_100 0 n12 ns100 0 0.000256954961272
Gc6_101 0 n12 ns101 0 -2.19729899184e-05
Gc6_102 0 n12 ns102 0 -8.67709110063e-05
Gc6_103 0 n12 ns103 0 7.86687932152e-05
Gc6_104 0 n12 ns104 0 -0.000106804328432
Gc6_105 0 n12 ns105 0 0.00149707817867
Gc6_106 0 n12 ns106 0 -2.77376184344e-05
Gc6_107 0 n12 ns107 0 9.56192774145e-05
Gc6_108 0 n12 ns108 0 0.000365635111469
Gc6_109 0 n12 ns109 0 6.29306681565e-06
Gc6_110 0 n12 ns110 0 -3.13979568489e-05
Gc6_111 0 n12 ns111 0 3.55055239812e-05
Gc6_112 0 n12 ns112 0 4.02693941813e-05
Gc6_113 0 n12 ns113 0 -0.000197644096907
Gc6_114 0 n12 ns114 0 3.71856038516e-06
Gc6_115 0 n12 ns115 0 -2.96761530611e-05
Gc6_116 0 n12 ns116 0 -6.84239109954e-05
Gc6_117 0 n12 ns117 0 -8.72545595793e-05
Gc6_118 0 n12 ns118 0 -4.44639783948e-05
Gc6_119 0 n12 ns119 0 -9.11733947175e-06
Gc6_120 0 n12 ns120 0 -1.67098809391e-05
Gc6_121 0 n12 ns121 0 2.49742273719e-05
Gc6_122 0 n12 ns122 0 -3.0343412114e-07
Gc6_123 0 n12 ns123 0 3.28404612067e-06
Gc6_124 0 n12 ns124 0 -6.65294054959e-06
Gc6_125 0 n12 ns125 0 -5.68851717827e-06
Gc6_126 0 n12 ns126 0 2.88112556534e-06
Gc6_127 0 n12 ns127 0 4.36333198941e-07
Gc6_128 0 n12 ns128 0 1.67218921582e-06
Gd6_1 0 n12 ni1 0 2.51435809681e-05
Gd6_2 0 n12 ni2 0 7.60703473324e-06
Gd6_3 0 n12 ni3 0 -4.14097054281e-05
Gd6_4 0 n12 ni4 0 0.000250444533447
Gd6_5 0 n12 ni5 0 1.85714678132e-05
Gd6_6 0 n12 ni6 0 -0.00130410328626
Gd6_7 0 n12 ni7 0 0.000167381039216
Gd6_8 0 n12 ni8 0 0.000250438701042
Gd6_9 0 n12 ni9 0 -5.81284818004e-05
Gd6_10 0 n12 ni10 0 -6.80860260315e-06
Gd6_11 0 n12 ni11 0 4.7284329438e-05
Gd6_12 0 n12 ni12 0 0.000810857298176
Gd6_13 0 n12 ni13 0 0.0024732842148
Gd6_14 0 n12 ni14 0 0.00027836586366
Gd6_15 0 n12 ni15 0 0.000292672877309
Gd6_16 0 n12 ni16 0 -1.17284404978e-05
Gc7_1 0 n14 ns1 0 -1.32249483454e-05
Gc7_2 0 n14 ns2 0 2.83410547229e-07
Gc7_3 0 n14 ns3 0 -1.61625567114e-06
Gc7_4 0 n14 ns4 0 -2.84037829234e-06
Gc7_5 0 n14 ns5 0 -4.75881817387e-06
Gc7_6 0 n14 ns6 0 -1.80587315176e-07
Gc7_7 0 n14 ns7 0 -7.15829998279e-07
Gc7_8 0 n14 ns8 0 -1.02093447752e-06
Gc7_9 0 n14 ns9 0 -1.43956027769e-05
Gc7_10 0 n14 ns10 0 3.07874694091e-07
Gc7_11 0 n14 ns11 0 -1.77502818613e-06
Gc7_12 0 n14 ns12 0 -4.1324000856e-06
Gc7_13 0 n14 ns13 0 -5.13919841725e-06
Gc7_14 0 n14 ns14 0 -6.7150129803e-07
Gc7_15 0 n14 ns15 0 -7.04269457944e-07
Gc7_16 0 n14 ns16 0 -1.06363861359e-06
Gc7_17 0 n14 ns17 0 4.59036299543e-07
Gc7_18 0 n14 ns18 0 4.08272732409e-08
Gc7_19 0 n14 ns19 0 1.15919400617e-07
Gc7_20 0 n14 ns20 0 -5.11515573862e-06
Gc7_21 0 n14 ns21 0 -2.70796449419e-06
Gc7_22 0 n14 ns22 0 -1.89877957179e-07
Gc7_23 0 n14 ns23 0 3.38233236775e-08
Gc7_24 0 n14 ns24 0 9.13761507797e-08
Gc7_25 0 n14 ns25 0 4.3280521616e-05
Gc7_26 0 n14 ns26 0 -6.98886134231e-07
Gc7_27 0 n14 ns27 0 5.65606584615e-06
Gc7_28 0 n14 ns28 0 1.37652488969e-06
Gc7_29 0 n14 ns29 0 3.73145319615e-06
Gc7_30 0 n14 ns30 0 5.55296473603e-06
Gc7_31 0 n14 ns31 0 1.43839252755e-06
Gc7_32 0 n14 ns32 0 2.99980129396e-06
Gc7_33 0 n14 ns33 0 -0.000185335650556
Gc7_34 0 n14 ns34 0 3.96983473583e-06
Gc7_35 0 n14 ns35 0 -2.59514998832e-05
Gc7_36 0 n14 ns36 0 -5.36050550876e-05
Gc7_37 0 n14 ns37 0 -5.19036319829e-05
Gc7_38 0 n14 ns38 0 -1.67076827822e-05
Gc7_39 0 n14 ns39 0 -6.74781351401e-06
Gc7_40 0 n14 ns40 0 -1.53385987311e-05
Gc7_41 0 n14 ns41 0 0.000265667925407
Gc7_42 0 n14 ns42 0 -6.05006730401e-06
Gc7_43 0 n14 ns43 0 1.29188054699e-05
Gc7_44 0 n14 ns44 0 1.26795103389e-05
Gc7_45 0 n14 ns45 0 -6.41898569531e-05
Gc7_46 0 n14 ns46 0 -5.99813016744e-05
Gc7_47 0 n14 ns47 0 8.51129878975e-06
Gc7_48 0 n14 ns48 0 -1.87342241057e-06
Gc7_49 0 n14 ns49 0 0.00252672950751
Gc7_50 0 n14 ns50 0 -4.23427435523e-05
Gc7_51 0 n14 ns51 0 0.000247422522001
Gc7_52 0 n14 ns52 0 0.000561916613217
Gc7_53 0 n14 ns53 0 0.00014366750007
Gc7_54 0 n14 ns54 0 -8.95220590544e-05
Gc7_55 0 n14 ns55 0 -5.08809757423e-05
Gc7_56 0 n14 ns56 0 0.000370950151909
Gc7_57 0 n14 ns57 0 7.49175096802e-05
Gc7_58 0 n14 ns58 0 -1.73642781081e-06
Gc7_59 0 n14 ns59 0 -1.52967060364e-05
Gc7_60 0 n14 ns60 0 -3.06961507089e-05
Gc7_61 0 n14 ns61 0 -7.64195587177e-05
Gc7_62 0 n14 ns62 0 -6.15082011574e-05
Gc7_63 0 n14 ns63 0 6.6173309757e-06
Gc7_64 0 n14 ns64 0 -2.16660931945e-05
Gc7_65 0 n14 ns65 0 -0.000164031663959
Gc7_66 0 n14 ns66 0 3.61425644525e-06
Gc7_67 0 n14 ns67 0 -2.30213813331e-05
Gc7_68 0 n14 ns68 0 -4.55445940404e-05
Gc7_69 0 n14 ns69 0 -5.00342643617e-05
Gc7_70 0 n14 ns70 0 -1.02271746557e-05
Gc7_71 0 n14 ns71 0 -6.20572113447e-06
Gc7_72 0 n14 ns72 0 -1.48916458481e-05
Gc7_73 0 n14 ns73 0 -1.8158363826e-05
Gc7_74 0 n14 ns74 0 4.05326032232e-07
Gc7_75 0 n14 ns75 0 -2.35741384158e-06
Gc7_76 0 n14 ns76 0 -5.89937008003e-06
Gc7_77 0 n14 ns77 0 -5.52301346989e-06
Gc7_78 0 n14 ns78 0 -7.95713720175e-07
Gc7_79 0 n14 ns79 0 -7.23722378015e-07
Gc7_80 0 n14 ns80 0 -1.39876001982e-06
Gc7_81 0 n14 ns81 0 2.38015583146e-05
Gc7_82 0 n14 ns82 0 -3.69909008961e-07
Gc7_83 0 n14 ns83 0 3.1607323937e-06
Gc7_84 0 n14 ns84 0 -6.8273550187e-07
Gc7_85 0 n14 ns85 0 1.05209706713e-06
Gc7_86 0 n14 ns86 0 3.18284146995e-06
Gc7_87 0 n14 ns87 0 7.77163351346e-07
Gc7_88 0 n14 ns88 0 1.64429010908e-06
Gc7_89 0 n14 ns89 0 -3.71484658488e-05
Gc7_90 0 n14 ns90 0 1.19239921646e-06
Gc7_91 0 n14 ns91 0 -6.02747130247e-06
Gc7_92 0 n14 ns92 0 -1.02175138137e-05
Gc7_93 0 n14 ns93 0 -6.17739226687e-06
Gc7_94 0 n14 ns94 0 7.8737526254e-06
Gc7_95 0 n14 ns95 0 -9.3491035228e-07
Gc7_96 0 n14 ns96 0 -4.51265653881e-06
Gc7_97 0 n14 ns97 0 -0.000484216598759
Gc7_98 0 n14 ns98 0 1.02918651775e-05
Gc7_99 0 n14 ns99 0 -7.2965704598e-05
Gc7_100 0 n14 ns100 0 -0.000121637761668
Gc7_101 0 n14 ns101 0 -0.000105129323102
Gc7_102 0 n14 ns102 0 -4.37236830194e-05
Gc7_103 0 n14 ns103 0 -1.33430652445e-05
Gc7_104 0 n14 ns104 0 -4.59131508424e-05
Gc7_105 0 n14 ns105 0 0.00137176778548
Gc7_106 0 n14 ns106 0 -1.9904764203e-05
Gc7_107 0 n14 ns107 0 -3.52296360878e-05
Gc7_108 0 n14 ns108 0 0.000272558677495
Gc7_109 0 n14 ns109 0 -1.8018015396e-05
Gc7_110 0 n14 ns110 0 -8.26127163015e-05
Gc7_111 0 n14 ns111 0 7.5050040962e-05
Gc7_112 0 n14 ns112 0 -9.14140787572e-05
Gc7_113 0 n14 ns113 0 0.00165839741184
Gc7_114 0 n14 ns114 0 -3.12754648103e-05
Gc7_115 0 n14 ns115 0 0.000119646576834
Gc7_116 0 n14 ns116 0 0.000413688292917
Gc7_117 0 n14 ns117 0 1.10293839642e-05
Gc7_118 0 n14 ns118 0 -2.78062261647e-05
Gc7_119 0 n14 ns119 0 3.400431767e-05
Gc7_120 0 n14 ns120 0 6.01108407527e-05
Gc7_121 0 n14 ns121 0 -0.000256580224924
Gc7_122 0 n14 ns122 0 5.11243805401e-06
Gc7_123 0 n14 ns123 0 -3.79884825281e-05
Gc7_124 0 n14 ns124 0 -7.55284999659e-05
Gc7_125 0 n14 ns125 0 -9.15406838338e-05
Gc7_126 0 n14 ns126 0 -4.07896820163e-05
Gc7_127 0 n14 ns127 0 -1.05721660025e-05
Gc7_128 0 n14 ns128 0 -2.23556028986e-05
Gd7_1 0 n14 ni1 0 1.25802383049e-05
Gd7_2 0 n14 ni2 0 1.43812698675e-05
Gd7_3 0 n14 ni3 0 3.01232302647e-06
Gd7_4 0 n14 ni4 0 -3.4805545205e-05
Gd7_5 0 n14 ni5 0 0.00022598784627
Gd7_6 0 n14 ni6 0 0.000167381039216
Gd7_7 0 n14 ni7 0 -0.000918847890765
Gd7_8 0 n14 ni8 0 0.000395998249606
Gd7_9 0 n14 ni9 0 0.000203158931799
Gd7_10 0 n14 ni10 0 1.98783978471e-05
Gd7_11 0 n14 ni11 0 -1.85967621534e-05
Gd7_12 0 n14 ni12 0 5.84805551825e-05
Gd7_13 0 n14 ni13 0 0.000645280734517
Gd7_14 0 n14 ni14 0 0.00227778946994
Gd7_15 0 n14 ni15 0 8.12469634996e-05
Gd7_16 0 n14 ni16 0 0.000354792270976
Gc8_1 0 n16 ns1 0 -3.79933865695e-06
Gc8_2 0 n16 ns2 0 9.26575079366e-08
Gc8_3 0 n16 ns3 0 -4.6585241826e-07
Gc8_4 0 n16 ns4 0 -6.70550860828e-07
Gc8_5 0 n16 ns5 0 -1.59604541563e-06
Gc8_6 0 n16 ns6 0 4.38427267323e-07
Gc8_7 0 n16 ns7 0 -2.49472249676e-07
Gc8_8 0 n16 ns8 0 -3.31086261474e-07
Gc8_9 0 n16 ns9 0 -5.92132847777e-06
Gc8_10 0 n16 ns10 0 1.33479806124e-07
Gc8_11 0 n16 ns11 0 -7.19054638995e-07
Gc8_12 0 n16 ns12 0 -1.18706051592e-06
Gc8_13 0 n16 ns13 0 -2.33458023821e-06
Gc8_14 0 n16 ns14 0 2.06921765449e-07
Gc8_15 0 n16 ns15 0 -3.57348366654e-07
Gc8_16 0 n16 ns16 0 -4.71494958902e-07
Gc8_17 0 n16 ns17 0 -1.19625816287e-05
Gc8_18 0 n16 ns18 0 2.62646452171e-07
Gc8_19 0 n16 ns19 0 -1.52906907275e-06
Gc8_20 0 n16 ns20 0 -4.34176643557e-06
Gc8_21 0 n16 ns21 0 -3.90455962093e-06
Gc8_22 0 n16 ns22 0 -7.43265055281e-07
Gc8_23 0 n16 ns23 0 -4.77460262438e-07
Gc8_24 0 n16 ns24 0 -8.86443564675e-07
Gc8_25 0 n16 ns25 0 -6.79808647133e-06
Gc8_26 0 n16 ns26 0 1.93351006335e-07
Gc8_27 0 n16 ns27 0 -8.43279871695e-07
Gc8_28 0 n16 ns28 0 -5.14154465606e-06
Gc8_29 0 n16 ns29 0 -4.11077977791e-06
Gc8_30 0 n16 ns30 0 -1.50817841073e-08
Gc8_31 0 n16 ns31 0 -3.21519209221e-07
Gc8_32 0 n16 ns32 0 -5.24812425234e-07
Gc8_33 0 n16 ns33 0 5.02184661993e-05
Gc8_34 0 n16 ns34 0 -8.49006009216e-07
Gc8_35 0 n16 ns35 0 6.75616558048e-06
Gc8_36 0 n16 ns36 0 3.45485942298e-06
Gc8_37 0 n16 ns37 0 3.43105159953e-06
Gc8_38 0 n16 ns38 0 6.30534242317e-06
Gc8_39 0 n16 ns39 0 1.44222411758e-06
Gc8_40 0 n16 ns40 0 3.55333625778e-06
Gc8_41 0 n16 ns41 0 -0.00020740116331
Gc8_42 0 n16 ns42 0 4.60119408212e-06
Gc8_43 0 n16 ns43 0 -2.94944542424e-05
Gc8_44 0 n16 ns44 0 -4.99524118779e-05
Gc8_45 0 n16 ns45 0 -4.74496175099e-05
Gc8_46 0 n16 ns46 0 -9.9856156687e-06
Gc8_47 0 n16 ns47 0 -7.04326277586e-06
Gc8_48 0 n16 ns48 0 -1.81008981411e-05
Gc8_49 0 n16 ns49 0 7.49175096802e-05
Gc8_50 0 n16 ns50 0 -1.73642781081e-06
Gc8_51 0 n16 ns51 0 -1.52967060364e-05
Gc8_52 0 n16 ns52 0 -3.06961507089e-05
Gc8_53 0 n16 ns53 0 -7.64195587177e-05
Gc8_54 0 n16 ns54 0 -6.15082011574e-05
Gc8_55 0 n16 ns55 0 6.6173309757e-06
Gc8_56 0 n16 ns56 0 -2.16660931945e-05
Gc8_57 0 n16 ns57 0 0.00265068571292
Gc8_58 0 n16 ns58 0 -4.63422067564e-05
Gc8_59 0 n16 ns59 0 0.000301883953253
Gc8_60 0 n16 ns60 0 0.000682405277562
Gc8_61 0 n16 ns61 0 0.000135725260441
Gc8_62 0 n16 ns62 0 -4.9571669476e-05
Gc8_63 0 n16 ns63 0 -7.46922885996e-05
Gc8_64 0 n16 ns64 0 0.000428364502461
Gc8_65 0 n16 ns65 0 0.000330002744625
Gc8_66 0 n16 ns66 0 -8.13869525014e-06
Gc8_67 0 n16 ns67 0 2.18106063738e-05
Gc8_68 0 n16 ns68 0 -8.63739854298e-06
Gc8_69 0 n16 ns69 0 -8.93356830086e-05
Gc8_70 0 n16 ns70 0 -8.68911670181e-05
Gc8_71 0 n16 ns71 0 1.17945666e-05
Gc8_72 0 n16 ns72 0 4.16393846586e-09
Gc8_73 0 n16 ns73 0 -1.18704870009e-05
Gc8_74 0 n16 ns74 0 2.59611373042e-07
Gc8_75 0 n16 ns75 0 -1.50881676156e-06
Gc8_76 0 n16 ns76 0 -2.4640876965e-06
Gc8_77 0 n16 ns77 0 -3.6464821954e-06
Gc8_78 0 n16 ns78 0 -8.27375125007e-08
Gc8_79 0 n16 ns79 0 -5.7864499779e-07
Gc8_80 0 n16 ns80 0 -9.37000376159e-07
Gc8_81 0 n16 ns81 0 -1.76714168234e-05
Gc8_82 0 n16 ns82 0 3.94205703298e-07
Gc8_83 0 n16 ns83 0 -2.27381542719e-06
Gc8_84 0 n16 ns84 0 -5.76759359869e-06
Gc8_85 0 n16 ns85 0 -5.63545858265e-06
Gc8_86 0 n16 ns86 0 -7.51815963e-07
Gc8_87 0 n16 ns87 0 -7.31729746798e-07
Gc8_88 0 n16 ns88 0 -1.35997020768e-06
Gc8_89 0 n16 ns89 0 3.21564792953e-06
Gc8_90 0 n16 ns90 0 7.31680437336e-08
Gc8_91 0 n16 ns91 0 2.31976484929e-07
Gc8_92 0 n16 ns92 0 -3.09292155676e-06
Gc8_93 0 n16 ns93 0 -8.90160615925e-07
Gc8_94 0 n16 ns94 0 2.85923054656e-06
Gc8_95 0 n16 ns95 0 1.77014318363e-07
Gc8_96 0 n16 ns96 0 -9.74156757754e-08
Gc8_97 0 n16 ns97 0 -5.80713728419e-05
Gc8_98 0 n16 ns98 0 1.62707471882e-06
Gc8_99 0 n16 ns99 0 -8.8035330078e-06
Gc8_100 0 n16 ns100 0 -1.3610215698e-05
Gc8_101 0 n16 ns101 0 -9.89053589508e-06
Gc8_102 0 n16 ns102 0 7.05833321937e-06
Gc8_103 0 n16 ns103 0 -1.67633297849e-06
Gc8_104 0 n16 ns104 0 -6.17803511118e-06
Gc8_105 0 n16 ns105 0 -0.000509645790512
Gc8_106 0 n16 ns106 0 1.08935729103e-05
Gc8_107 0 n16 ns107 0 -7.66570916483e-05
Gc8_108 0 n16 ns108 0 -0.000126985881327
Gc8_109 0 n16 ns109 0 -0.000105475676385
Gc8_110 0 n16 ns110 0 -4.23687299047e-05
Gc8_111 0 n16 ns111 0 -1.34163503852e-05
Gc8_112 0 n16 ns112 0 -4.87964106455e-05
Gc8_113 0 n16 ns113 0 0.00144473529064
Gc8_114 0 n16 ns114 0 -2.05880173706e-05
Gc8_115 0 n16 ns115 0 -5.54711214874e-05
Gc8_116 0 n16 ns116 0 0.000188893872145
Gc8_117 0 n16 ns117 0 1.04584877974e-05
Gc8_118 0 n16 ns118 0 -0.000114412392334
Gc8_119 0 n16 ns119 0 0.00010295429238
Gc8_120 0 n16 ns120 0 -0.000128225056716
Gc8_121 0 n16 ns121 0 0.00174499801323
Gc8_122 0 n16 ns122 0 -3.3215408067e-05
Gc8_123 0 n16 ns123 0 0.000130973727851
Gc8_124 0 n16 ns124 0 0.000449511823642
Gc8_125 0 n16 ns125 0 -3.95091382585e-06
Gc8_126 0 n16 ns126 0 -2.86444539224e-05
Gc8_127 0 n16 ns127 0 3.08449940804e-05
Gc8_128 0 n16 ns128 0 6.94405872255e-05
Gd8_1 0 n16 ni1 0 3.78622145149e-06
Gd8_2 0 n16 ni2 0 5.68761425467e-06
Gd8_3 0 n16 ni3 0 1.3045771699e-05
Gd8_4 0 n16 ni4 0 9.63805909615e-06
Gd8_5 0 n16 ni5 0 -4.40192767264e-05
Gd8_6 0 n16 ni6 0 0.000250438701042
Gd8_7 0 n16 ni7 0 0.000395998249606
Gd8_8 0 n16 ni8 0 -0.00167941484723
Gd8_9 0 n16 ni9 0 0.000129164128304
Gd8_10 0 n16 ni10 0 1.18410244839e-05
Gd8_11 0 n16 ni11 0 1.91867465127e-05
Gd8_12 0 n16 ni12 0 3.40773102046e-06
Gd8_13 0 n16 ni13 0 7.9012564602e-05
Gd8_14 0 n16 ni14 0 0.000673903454497
Gd8_15 0 n16 ni15 0 0.00271939044449
Gd8_16 0 n16 ni16 0 5.70965984872e-06
Gc9_1 0 n18 ns1 0 5.10187713518e-07
Gc9_2 0 n18 ns2 0 5.26057012904e-09
Gc9_3 0 n18 ns3 0 6.29743488324e-08
Gc9_4 0 n18 ns4 0 -2.93206361134e-07
Gc9_5 0 n18 ns5 0 -2.77246705676e-07
Gc9_6 0 n18 ns6 0 5.26181318434e-07
Gc9_7 0 n18 ns7 0 -4.56625062906e-09
Gc9_8 0 n18 ns8 0 -1.91908117476e-09
Gc9_9 0 n18 ns9 0 -1.69854637436e-06
Gc9_10 0 n18 ns10 0 4.8167449143e-08
Gc9_11 0 n18 ns11 0 -1.92968863617e-07
Gc9_12 0 n18 ns12 0 -2.43468214806e-07
Gc9_13 0 n18 ns13 0 -1.05675369117e-06
Gc9_14 0 n18 ns14 0 5.24336706599e-07
Gc9_15 0 n18 ns15 0 -1.60597604508e-07
Gc9_16 0 n18 ns16 0 -1.67112279397e-07
Gc9_17 0 n18 ns17 0 -5.38569718614e-06
Gc9_18 0 n18 ns18 0 1.20928343182e-07
Gc9_19 0 n18 ns19 0 -6.19617568441e-07
Gc9_20 0 n18 ns20 0 -1.42170536585e-06
Gc9_21 0 n18 ns21 0 -2.61192606132e-06
Gc9_22 0 n18 ns22 0 1.45873987595e-07
Gc9_23 0 n18 ns23 0 -3.55447237246e-07
Gc9_24 0 n18 ns24 0 -4.19395235924e-07
Gc9_25 0 n18 ns25 0 -1.74728450152e-05
Gc9_26 0 n18 ns26 0 3.67151640903e-07
Gc9_27 0 n18 ns27 0 -2.09229230608e-06
Gc9_28 0 n18 ns28 0 -4.2837217456e-06
Gc9_29 0 n18 ns29 0 -6.77155368265e-06
Gc9_30 0 n18 ns30 0 -6.34773702603e-07
Gc9_31 0 n18 ns31 0 -9.60648440033e-07
Gc9_32 0 n18 ns32 0 -1.30456977862e-06
Gc9_33 0 n18 ns33 0 2.35174293607e-06
Gc9_34 0 n18 ns34 0 -2.08109595048e-08
Gc9_35 0 n18 ns35 0 7.20481168481e-07
Gc9_36 0 n18 ns36 0 -4.07483878871e-06
Gc9_37 0 n18 ns37 0 -6.22805854561e-06
Gc9_38 0 n18 ns38 0 1.01369202911e-07
Gc9_39 0 n18 ns39 0 -3.80974860043e-07
Gc9_40 0 n18 ns40 0 2.89974094324e-07
Gc9_41 0 n18 ns41 0 6.31549198078e-05
Gc9_42 0 n18 ns42 0 -1.13676191605e-06
Gc9_43 0 n18 ns43 0 8.72455823149e-06
Gc9_44 0 n18 ns44 0 4.21748439968e-06
Gc9_45 0 n18 ns45 0 2.16334025006e-06
Gc9_46 0 n18 ns46 0 6.34016736344e-06
Gc9_47 0 n18 ns47 0 1.66622588384e-06
Gc9_48 0 n18 ns48 0 4.52368549783e-06
Gc9_49 0 n18 ns49 0 -0.000164031663959
Gc9_50 0 n18 ns50 0 3.61425644525e-06
Gc9_51 0 n18 ns51 0 -2.30213813331e-05
Gc9_52 0 n18 ns52 0 -4.55445940404e-05
Gc9_53 0 n18 ns53 0 -5.00342643617e-05
Gc9_54 0 n18 ns54 0 -1.02271746557e-05
Gc9_55 0 n18 ns55 0 -6.20572113447e-06
Gc9_56 0 n18 ns56 0 -1.48916458481e-05
Gc9_57 0 n18 ns57 0 0.000330002744625
Gc9_58 0 n18 ns58 0 -8.13869525014e-06
Gc9_59 0 n18 ns59 0 2.18106063738e-05
Gc9_60 0 n18 ns60 0 -8.63739854298e-06
Gc9_61 0 n18 ns61 0 -8.93356830086e-05
Gc9_62 0 n18 ns62 0 -8.68911670181e-05
Gc9_63 0 n18 ns63 0 1.17945666e-05
Gc9_64 0 n18 ns64 0 4.16393846541e-09
Gc9_65 0 n18 ns65 0 0.00447103859283
Gc9_66 0 n18 ns66 0 -8.71355693377e-05
Gc9_67 0 n18 ns67 0 0.000544719039683
Gc9_68 0 n18 ns68 0 0.00104224456672
Gc9_69 0 n18 ns69 0 0.000245662679521
Gc9_70 0 n18 ns70 0 -4.61696271876e-05
Gc9_71 0 n18 ns71 0 -3.16758643009e-05
Gc9_72 0 n18 ns72 0 0.000563097946123
Gc9_73 0 n18 ns73 0 -5.92409363623e-06
Gc9_74 0 n18 ns74 0 1.35162811158e-07
Gc9_75 0 n18 ns75 0 -7.14935622347e-07
Gc9_76 0 n18 ns76 0 -4.59570842479e-07
Gc9_77 0 n18 ns77 0 -2.30809716247e-06
Gc9_78 0 n18 ns78 0 5.47373051715e-07
Gc9_79 0 n18 ns79 0 -4.06415858044e-07
Gc9_80 0 n18 ns80 0 -5.02294444305e-07
Gc9_81 0 n18 ns81 0 -1.5419832129e-05
Gc9_82 0 n18 ns82 0 3.25292769669e-07
Gc9_83 0 n18 ns83 0 -1.85335220289e-06
Gc9_84 0 n18 ns84 0 -2.63829970893e-06
Gc9_85 0 n18 ns85 0 -5.70944781269e-06
Gc9_86 0 n18 ns86 0 -9.73234243709e-08
Gc9_87 0 n18 ns87 0 -8.99775786879e-07
Gc9_88 0 n18 ns88 0 -1.19271034738e-06
Gc9_89 0 n18 ns89 0 -2.49793592217e-05
Gc9_90 0 n18 ns90 0 5.40516314283e-07
Gc9_91 0 n18 ns91 0 -3.14309379312e-06
Gc9_92 0 n18 ns92 0 -6.68313219359e-06
Gc9_93 0 n18 ns93 0 -8.24037559619e-06
Gc9_94 0 n18 ns94 0 -9.10413982197e-07
Gc9_95 0 n18 ns95 0 -1.15451486137e-06
Gc9_96 0 n18 ns96 0 -1.94041204534e-06
Gc9_97 0 n18 ns97 0 1.88210583904e-05
Gc9_98 0 n18 ns98 0 -2.69854602772e-07
Gc9_99 0 n18 ns99 0 2.66949826623e-06
Gc9_100 0 n18 ns100 0 -1.07677517272e-06
Gc9_101 0 n18 ns101 0 -2.10239898931e-06
Gc9_102 0 n18 ns102 0 3.41959928295e-06
Gc9_103 0 n18 ns103 0 3.41659712889e-07
Gc9_104 0 n18 ns104 0 1.18079277049e-06
Gc9_105 0 n18 ns105 0 -5.0365213296e-07
Gc9_106 0 n18 ns106 0 3.51908736282e-07
Gc9_107 0 n18 ns107 0 -4.39712265447e-07
Gc9_108 0 n18 ns108 0 -6.51743635438e-06
Gc9_109 0 n18 ns109 0 -9.05676342661e-06
Gc9_110 0 n18 ns110 0 7.47567841332e-06
Gc9_111 0 n18 ns111 0 -3.8913972992e-07
Gc9_112 0 n18 ns112 0 -1.57067038167e-06
Gc9_113 0 n18 ns113 0 -0.000554674208466
Gc9_114 0 n18 ns114 0 1.188018418e-05
Gc9_115 0 n18 ns115 0 -8.29650683047e-05
Gc9_116 0 n18 ns116 0 -0.000143447072203
Gc9_117 0 n18 ns117 0 -0.000114352221074
Gc9_118 0 n18 ns118 0 -4.40566211289e-05
Gc9_119 0 n18 ns119 0 -1.35817526434e-05
Gc9_120 0 n18 ns120 0 -5.43520905485e-05
Gc9_121 0 n18 ns121 0 0.00234877905334
Gc9_122 0 n18 ns122 0 -4.17321968383e-05
Gc9_123 0 n18 ns123 0 7.28214005941e-05
Gc9_124 0 n18 ns124 0 0.000252875440643
Gc9_125 0 n18 ns125 0 9.52922970868e-05
Gc9_126 0 n18 ns126 0 -0.000147858583895
Gc9_127 0 n18 ns127 0 0.000139262885025
Gc9_128 0 n18 ns128 0 -6.09760253552e-05
Gd9_1 0 n18 ni1 0 7.03349055233e-08
Gd9_2 0 n18 ni2 0 1.67449036216e-06
Gd9_3 0 n18 ni3 0 5.06716986895e-06
Gd9_4 0 n18 ni4 0 1.64120887921e-05
Gd9_5 0 n18 ni5 0 -2.64877748396e-06
Gd9_6 0 n18 ni6 0 -5.81284818004e-05
Gd9_7 0 n18 ni7 0 0.000203158931799
Gd9_8 0 n18 ni8 0 0.000129164128304
Gd9_9 0 n18 ni9 0 -0.00341147906647
Gd9_10 0 n18 ni10 0 5.28783804493e-06
Gd9_11 0 n18 ni11 0 1.39314255723e-05
Gd9_12 0 n18 ni12 0 2.5381392322e-05
Gd9_13 0 n18 ni13 0 -1.52609614812e-05
Gd9_14 0 n18 ni14 0 1.70281693251e-05
Gd9_15 0 n18 ni15 0 0.000728441936391
Gd9_16 0 n18 ni16 0 0.0017656377046
Gc10_1 0 n20 ns1 0 0.000255627852429
Gc10_2 0 n20 ns2 0 -6.42873416842e-06
Gc10_3 0 n20 ns3 0 1.23217762639e-05
Gc10_4 0 n20 ns4 0 2.02328290634e-06
Gc10_5 0 n20 ns5 0 -0.000111142392723
Gc10_6 0 n20 ns6 0 -8.6404752839e-05
Gc10_7 0 n20 ns7 0 3.3281281639e-06
Gc10_8 0 n20 ns8 0 3.28649442323e-07
Gc10_9 0 n20 ns9 0 0.00200724653791
Gc10_10 0 n20 ns10 0 -3.91419194742e-05
Gc10_11 0 n20 ns11 0 0.000172003051018
Gc10_12 0 n20 ns12 0 0.000506691300361
Gc10_13 0 n20 ns13 0 2.3999336226e-05
Gc10_14 0 n20 ns14 0 -1.98679104574e-05
Gc10_15 0 n20 ns15 0 3.49336170623e-05
Gc10_16 0 n20 ns16 0 9.69560154653e-05
Gc10_17 0 n20 ns17 0 0.00146919185322
Gc10_18 0 n20 ns18 0 -2.12857910264e-05
Gc10_19 0 n20 ns19 0 -4.2977754716e-05
Gc10_20 0 n20 ns20 0 0.000246698064877
Gc10_21 0 n20 ns21 0 1.24625551941e-06
Gc10_22 0 n20 ns22 0 -9.54218550464e-05
Gc10_23 0 n20 ns23 0 9.24107291793e-05
Gc10_24 0 n20 ns24 0 -0.000112217613401
Gc10_25 0 n20 ns25 0 -0.000528989617471
Gc10_26 0 n20 ns26 0 1.12284364269e-05
Gc10_27 0 n20 ns27 0 -7.89151534504e-05
Gc10_28 0 n20 ns28 0 -0.00012915155275
Gc10_29 0 n20 ns29 0 -0.000113282011914
Gc10_30 0 n20 ns30 0 -4.54158863742e-05
Gc10_31 0 n20 ns31 0 -1.49383207297e-05
Gc10_32 0 n20 ns32 0 -4.94848425366e-05
Gc10_33 0 n20 ns33 0 -7.09137768122e-05
Gc10_34 0 n20 ns34 0 1.94024935126e-06
Gc10_35 0 n20 ns35 0 -1.06275646452e-05
Gc10_36 0 n20 ns36 0 -1.3552784779e-05
Gc10_37 0 n20 ns37 0 -1.02410512869e-05
Gc10_38 0 n20 ns38 0 8.57758204151e-06
Gc10_39 0 n20 ns39 0 -2.10086364247e-06
Gc10_40 0 n20 ns40 0 -7.35502662103e-06
Gc10_41 0 n20 ns41 0 1.22499948205e-05
Gc10_42 0 n20 ns42 0 -1.19278604293e-07
Gc10_43 0 n20 ns43 0 1.54394149213e-06
Gc10_44 0 n20 ns44 0 -1.45605242078e-06
Gc10_45 0 n20 ns45 0 -2.22156682214e-07
Gc10_46 0 n20 ns46 0 3.2872473059e-06
Gc10_47 0 n20 ns47 0 3.6405420909e-07
Gc10_48 0 n20 ns48 0 6.75091556278e-07
Gc10_49 0 n20 ns49 0 -1.8158363826e-05
Gc10_50 0 n20 ns50 0 4.05326032232e-07
Gc10_51 0 n20 ns51 0 -2.35741384158e-06
Gc10_52 0 n20 ns52 0 -5.89937008003e-06
Gc10_53 0 n20 ns53 0 -5.52301346989e-06
Gc10_54 0 n20 ns54 0 -7.95713720175e-07
Gc10_55 0 n20 ns55 0 -7.23722378015e-07
Gc10_56 0 n20 ns56 0 -1.39876001982e-06
Gc10_57 0 n20 ns57 0 -1.18704870009e-05
Gc10_58 0 n20 ns58 0 2.59611373042e-07
Gc10_59 0 n20 ns59 0 -1.50881676156e-06
Gc10_60 0 n20 ns60 0 -2.4640876965e-06
Gc10_61 0 n20 ns61 0 -3.6464821954e-06
Gc10_62 0 n20 ns62 0 -8.27375125007e-08
Gc10_63 0 n20 ns63 0 -5.7864499779e-07
Gc10_64 0 n20 ns64 0 -9.37000376159e-07
Gc10_65 0 n20 ns65 0 -5.92409363623e-06
Gc10_66 0 n20 ns66 0 1.35162811158e-07
Gc10_67 0 n20 ns67 0 -7.14935622347e-07
Gc10_68 0 n20 ns68 0 -4.59570842479e-07
Gc10_69 0 n20 ns69 0 -2.30809716247e-06
Gc10_70 0 n20 ns70 0 5.47373051715e-07
Gc10_71 0 n20 ns71 0 -4.06415858044e-07
Gc10_72 0 n20 ns72 0 -5.02294444305e-07
Gc10_73 0 n20 ns73 0 0.00277867191432
Gc10_74 0 n20 ns74 0 -4.90370137607e-05
Gc10_75 0 n20 ns75 0 0.000306089266341
Gc10_76 0 n20 ns76 0 0.000618440345291
Gc10_77 0 n20 ns77 0 0.00018735318894
Gc10_78 0 n20 ns78 0 -6.33849028944e-05
Gc10_79 0 n20 ns79 0 -4.67054713485e-05
Gc10_80 0 n20 ns80 0 0.000406953470228
Gc10_81 0 n20 ns81 0 9.8716610638e-05
Gc10_82 0 n20 ns82 0 -2.20861565649e-06
Gc10_83 0 n20 ns83 0 -1.2704020243e-05
Gc10_84 0 n20 ns84 0 -1.50693969712e-05
Gc10_85 0 n20 ns85 0 -8.27057918031e-05
Gc10_86 0 n20 ns86 0 -6.16506050773e-05
Gc10_87 0 n20 ns87 0 4.35468589959e-06
Gc10_88 0 n20 ns88 0 -1.78615327291e-05
Gc10_89 0 n20 ns89 0 -0.000215394845714
Gc10_90 0 n20 ns90 0 4.7261540694e-06
Gc10_91 0 n20 ns91 0 -3.03242023269e-05
Gc10_92 0 n20 ns92 0 -5.47917689852e-05
Gc10_93 0 n20 ns93 0 -5.11803003723e-05
Gc10_94 0 n20 ns94 0 -1.30055756667e-05
Gc10_95 0 n20 ns95 0 -7.48432894173e-06
Gc10_96 0 n20 ns96 0 -1.81064561441e-05
Gc10_97 0 n20 ns97 0 4.47462542728e-05
Gc10_98 0 n20 ns98 0 -7.25285384624e-07
Gc10_99 0 n20 ns99 0 5.94633949626e-06
Gc10_100 0 n20 ns100 0 3.06074772357e-06
Gc10_101 0 n20 ns101 0 3.33752671339e-06
Gc10_102 0 n20 ns102 0 6.42849685484e-06
Gc10_103 0 n20 ns103 0 1.3036293483e-06
Gc10_104 0 n20 ns104 0 3.08200797288e-06
Gc10_105 0 n20 ns105 0 -6.14856044072e-06
Gc10_106 0 n20 ns106 0 1.77772609317e-07
Gc10_107 0 n20 ns107 0 -7.47838813868e-07
Gc10_108 0 n20 ns108 0 -5.11477848383e-06
Gc10_109 0 n20 ns109 0 -4.07381072025e-06
Gc10_110 0 n20 ns110 0 -7.82809232336e-08
Gc10_111 0 n20 ns111 0 -3.0519607436e-07
Gc10_112 0 n20 ns112 0 -4.54462245249e-07
Gc10_113 0 n20 ns113 0 -1.21323220079e-05
Gc10_114 0 n20 ns114 0 2.63607267151e-07
Gc10_115 0 n20 ns115 0 -1.52679921289e-06
Gc10_116 0 n20 ns116 0 -4.29227603052e-06
Gc10_117 0 n20 ns117 0 -4.18063444018e-06
Gc10_118 0 n20 ns118 0 -7.67292975811e-07
Gc10_119 0 n20 ns119 0 -5.19017068953e-07
Gc10_120 0 n20 ns120 0 -8.87190430273e-07
Gc10_121 0 n20 ns121 0 -6.7935037963e-06
Gc10_122 0 n20 ns122 0 1.51215699355e-07
Gc10_123 0 n20 ns123 0 -8.21800021607e-07
Gc10_124 0 n20 ns124 0 -1.08234753819e-06
Gc10_125 0 n20 ns125 0 -2.62261287762e-06
Gc10_126 0 n20 ns126 0 2.64589779324e-07
Gc10_127 0 n20 ns127 0 -4.23445235459e-07
Gc10_128 0 n20 ns128 0 -5.4146526617e-07
Gd10_1 0 n20 ni1 0 0.000191911773795
Gd10_2 0 n20 ni2 0 -0.000349284122458
Gd10_3 0 n20 ni3 0 0.00253137732265
Gd10_4 0 n20 ni4 0 0.000689640310647
Gd10_5 0 n20 ni5 0 9.17481698985e-05
Gd10_6 0 n20 ni6 0 -6.80860260315e-06
Gd10_7 0 n20 ni7 0 1.98783978471e-05
Gd10_8 0 n20 ni8 0 1.18410244839e-05
Gd10_9 0 n20 ni9 0 5.28783804493e-06
Gd10_10 0 n20 ni10 0 -0.00158142851514
Gd10_11 0 n20 ni11 0 0.000382491287589
Gd10_12 0 n20 ni12 0 0.000257282980409
Gd10_13 0 n20 ni13 0 -3.79931894344e-05
Gd10_14 0 n20 ni14 0 8.92046372427e-06
Gd10_15 0 n20 ni15 0 1.29121964224e-05
Gd10_16 0 n20 ni16 0 6.30326646412e-06
Gc11_1 0 n22 ns1 0 -0.000193365998062
Gc11_2 0 n22 ns2 0 4.30579104473e-06
Gc11_3 0 n22 ns3 0 -2.71300115619e-05
Gc11_4 0 n22 ns4 0 -5.13233030284e-05
Gc11_5 0 n22 ns5 0 -5.19808613777e-05
Gc11_6 0 n22 ns6 0 -1.02447817267e-05
Gc11_7 0 n22 ns7 0 -7.07990052351e-06
Gc11_8 0 n22 ns8 0 -1.68316835908e-05
Gc11_9 0 n22 ns9 0 -0.000252088360404
Gc11_10 0 n22 ns10 0 4.93715114592e-06
Gc11_11 0 n22 ns11 0 -3.70945505007e-05
Gc11_12 0 n22 ns12 0 -7.48361684392e-05
Gc11_13 0 n22 ns13 0 -9.53200089991e-05
Gc11_14 0 n22 ns14 0 -4.33828894287e-05
Gc11_15 0 n22 ns15 0 -1.10705058984e-05
Gc11_16 0 n22 ns16 0 -2.13691782657e-05
Gc11_17 0 n22 ns17 0 0.0017314763145
Gc11_18 0 n22 ns18 0 -3.29028759871e-05
Gc11_19 0 n22 ns19 0 0.00012794972743
Gc11_20 0 n22 ns20 0 0.000424052302862
Gc11_21 0 n22 ns21 0 1.94550881083e-05
Gc11_22 0 n22 ns22 0 -2.65260469772e-05
Gc11_23 0 n22 ns23 0 3.83172714771e-05
Gc11_24 0 n22 ns24 0 6.11434746033e-05
Gc11_25 0 n22 ns25 0 0.00168679657982
Gc11_26 0 n22 ns26 0 -2.68448755633e-05
Gc11_27 0 n22 ns27 0 8.02085238536e-06
Gc11_28 0 n22 ns28 0 0.000337410115542
Gc11_29 0 n22 ns29 0 1.13479066436e-05
Gc11_30 0 n22 ns30 0 -7.58389803008e-05
Gc11_31 0 n22 ns31 0 8.25271002342e-05
Gc11_32 0 n22 ns32 0 -6.61406514889e-05
Gc11_33 0 n22 ns33 0 -0.000583120781668
Gc11_34 0 n22 ns34 0 1.24796099228e-05
Gc11_35 0 n22 ns35 0 -8.69690055429e-05
Gc11_36 0 n22 ns36 0 -0.000140598714665
Gc11_37 0 n22 ns37 0 -0.000114830909271
Gc11_38 0 n22 ns38 0 -4.53618394728e-05
Gc11_39 0 n22 ns39 0 -1.55582568209e-05
Gc11_40 0 n22 ns40 0 -5.46568832722e-05
Gc11_41 0 n22 ns41 0 -2.78564405109e-05
Gc11_42 0 n22 ns42 0 9.40051105009e-07
Gc11_43 0 n22 ns43 0 -4.48509036758e-06
Gc11_44 0 n22 ns44 0 -1.11321965317e-05
Gc11_45 0 n22 ns45 0 -8.18315057366e-06
Gc11_46 0 n22 ns46 0 5.86589387302e-06
Gc11_47 0 n22 ns47 0 -8.57782587434e-07
Gc11_48 0 n22 ns48 0 -3.44105375606e-06
Gc11_49 0 n22 ns49 0 2.38015583146e-05
Gc11_50 0 n22 ns50 0 -3.69909008961e-07
Gc11_51 0 n22 ns51 0 3.1607323937e-06
Gc11_52 0 n22 ns52 0 -6.8273550187e-07
Gc11_53 0 n22 ns53 0 1.05209706713e-06
Gc11_54 0 n22 ns54 0 3.18284146995e-06
Gc11_55 0 n22 ns55 0 7.77163351346e-07
Gc11_56 0 n22 ns56 0 1.64429010908e-06
Gc11_57 0 n22 ns57 0 -1.76714168234e-05
Gc11_58 0 n22 ns58 0 3.94205703298e-07
Gc11_59 0 n22 ns59 0 -2.27381542719e-06
Gc11_60 0 n22 ns60 0 -5.76759359869e-06
Gc11_61 0 n22 ns61 0 -5.63545858265e-06
Gc11_62 0 n22 ns62 0 -7.51815963e-07
Gc11_63 0 n22 ns63 0 -7.31729746798e-07
Gc11_64 0 n22 ns64 0 -1.35997020768e-06
Gc11_65 0 n22 ns65 0 -1.5419832129e-05
Gc11_66 0 n22 ns66 0 3.25292769669e-07
Gc11_67 0 n22 ns67 0 -1.85335220289e-06
Gc11_68 0 n22 ns68 0 -2.63829970893e-06
Gc11_69 0 n22 ns69 0 -5.70944781269e-06
Gc11_70 0 n22 ns70 0 -9.73234243709e-08
Gc11_71 0 n22 ns71 0 -8.99775786879e-07
Gc11_72 0 n22 ns72 0 -1.19271034738e-06
Gc11_73 0 n22 ns73 0 9.8716610638e-05
Gc11_74 0 n22 ns74 0 -2.20861565649e-06
Gc11_75 0 n22 ns75 0 -1.2704020243e-05
Gc11_76 0 n22 ns76 0 -1.50693969712e-05
Gc11_77 0 n22 ns77 0 -8.27057918031e-05
Gc11_78 0 n22 ns78 0 -6.16506050773e-05
Gc11_79 0 n22 ns79 0 4.35468589959e-06
Gc11_80 0 n22 ns80 0 -1.78615327291e-05
Gc11_81 0 n22 ns81 0 0.00270610029933
Gc11_82 0 n22 ns82 0 -4.69117304286e-05
Gc11_83 0 n22 ns83 0 0.000283163837132
Gc11_84 0 n22 ns84 0 0.000583960012308
Gc11_85 0 n22 ns85 0 0.000176696066992
Gc11_86 0 n22 ns86 0 -8.074103127e-05
Gc11_87 0 n22 ns87 0 -4.43041364769e-05
Gc11_88 0 n22 ns88 0 0.000390875404432
Gc11_89 0 n22 ns89 0 0.000442116787992
Gc11_90 0 n22 ns90 0 -1.01443573133e-05
Gc11_91 0 n22 ns91 0 3.83547234951e-05
Gc11_92 0 n22 ns92 0 5.04203755973e-05
Gc11_93 0 n22 ns93 0 -6.22391668012e-05
Gc11_94 0 n22 ns94 0 -6.44308210856e-05
Gc11_95 0 n22 ns95 0 9.7304023389e-06
Gc11_96 0 n22 ns96 0 1.58972729012e-05
Gc11_97 0 n22 ns97 0 -0.000190048829312
Gc11_98 0 n22 ns98 0 4.11001605983e-06
Gc11_99 0 n22 ns99 0 -2.66944890208e-05
Gc11_100 0 n22 ns100 0 -5.22496521261e-05
Gc11_101 0 n22 ns101 0 -5.09581626108e-05
Gc11_102 0 n22 ns102 0 -1.49314791451e-05
Gc11_103 0 n22 ns103 0 -6.87506922985e-06
Gc11_104 0 n22 ns104 0 -1.59122708761e-05
Gc11_105 0 n22 ns105 0 4.91963294168e-05
Gc11_106 0 n22 ns106 0 -8.28221363194e-07
Gc11_107 0 n22 ns107 0 6.51603091445e-06
Gc11_108 0 n22 ns108 0 2.33706720415e-06
Gc11_109 0 n22 ns109 0 4.10044312229e-06
Gc11_110 0 n22 ns110 0 5.69762813597e-06
Gc11_111 0 n22 ns111 0 1.56609725449e-06
Gc11_112 0 n22 ns112 0 3.50889444873e-06
Gc11_113 0 n22 ns113 0 3.46770648464e-06
Gc11_114 0 n22 ns114 0 -2.6788672598e-08
Gc11_115 0 n22 ns115 0 5.8011941478e-07
Gc11_116 0 n22 ns116 0 -4.57129846502e-06
Gc11_117 0 n22 ns117 0 -2.7914896606e-06
Gc11_118 0 n22 ns118 0 -1.04224118437e-07
Gc11_119 0 n22 ns119 0 6.42489359127e-08
Gc11_120 0 n22 ns120 0 3.55594397611e-07
Gc11_121 0 n22 ns121 0 -1.56385244704e-05
Gc11_122 0 n22 ns122 0 3.32252237804e-07
Gc11_123 0 n22 ns123 0 -1.91200169939e-06
Gc11_124 0 n22 ns124 0 -4.03261200512e-06
Gc11_125 0 n22 ns125 0 -5.66003742796e-06
Gc11_126 0 n22 ns126 0 -6.18188926581e-07
Gc11_127 0 n22 ns127 0 -8.07335886215e-07
Gc11_128 0 n22 ns128 0 -1.1585456105e-06
Gd11_1 0 n22 ni1 0 0.00023448060264
Gd11_2 0 n22 ni2 0 0.000347779628347
Gd11_3 0 n22 ni3 0 3.42237858478e-05
Gd11_4 0 n22 ni4 0 0.00195227228226
Gd11_5 0 n22 ni5 0 0.00075391676804
Gd11_6 0 n22 ni6 0 4.7284329438e-05
Gd11_7 0 n22 ni7 0 -1.85967621534e-05
Gd11_8 0 n22 ni8 0 1.91867465127e-05
Gd11_9 0 n22 ni9 0 1.39314255723e-05
Gd11_10 0 n22 ni10 0 0.000382491287589
Gd11_11 0 n22 ni11 0 -0.00128687178965
Gd11_12 0 n22 ni12 0 -2.77832584681e-05
Gd11_13 0 n22 ni13 0 0.00023077462273
Gd11_14 0 n22 ni14 0 -4.14425446025e-05
Gd11_15 0 n22 ni15 0 -6.65569976706e-07
Gd11_16 0 n22 ni16 0 1.51900969614e-05
Gc12_1 0 n24 ns1 0 7.63131403312e-05
Gc12_2 0 n24 ns2 0 -1.40056905352e-06
Gc12_3 0 n24 ns3 0 1.0545317299e-05
Gc12_4 0 n24 ns4 0 6.49273343603e-06
Gc12_5 0 n24 ns5 0 4.21332579687e-06
Gc12_6 0 n24 ns6 0 7.20418779089e-06
Gc12_7 0 n24 ns7 0 2.02985677331e-06
Gc12_8 0 n24 ns8 0 5.6811216195e-06
Gc12_9 0 n24 ns9 0 3.93712811119e-05
Gc12_10 0 n24 ns10 0 -6.35542271504e-07
Gc12_11 0 n24 ns11 0 5.44236055417e-06
Gc12_12 0 n24 ns12 0 -5.25514533149e-06
Gc12_13 0 n24 ns13 0 -5.4450295489e-06
Gc12_14 0 n24 ns14 0 2.39747494239e-06
Gc12_15 0 n24 ns15 0 7.29437069202e-07
Gc12_16 0 n24 ns16 0 3.03402833101e-06
Gc12_17 0 n24 ns17 0 -0.000190010036797
Gc12_18 0 n24 ns18 0 3.49364153638e-06
Gc12_19 0 n24 ns19 0 -2.83968096019e-05
Gc12_20 0 n24 ns20 0 -6.85762365233e-05
Gc12_21 0 n24 ns21 0 -8.98826290617e-05
Gc12_22 0 n24 ns22 0 -4.70144525347e-05
Gc12_23 0 n24 ns23 0 -9.36190505878e-06
Gc12_24 0 n24 ns24 0 -1.54310405027e-05
Gc12_25 0 n24 ns25 0 0.00174050680003
Gc12_26 0 n24 ns26 0 -3.32490526527e-05
Gc12_27 0 n24 ns27 0 0.000133089643448
Gc12_28 0 n24 ns28 0 0.0004330019464
Gc12_29 0 n24 ns29 0 1.83869460392e-05
Gc12_30 0 n24 ns30 0 -2.46137986848e-05
Gc12_31 0 n24 ns31 0 3.57447983553e-05
Gc12_32 0 n24 ns32 0 6.74656402172e-05
Gc12_33 0 n24 ns33 0 0.00203041538367
Gc12_34 0 n24 ns34 0 -3.29455410893e-05
Gc12_35 0 n24 ns35 0 8.31761413782e-06
Gc12_36 0 n24 ns36 0 0.000266181855967
Gc12_37 0 n24 ns37 0 7.56587628206e-05
Gc12_38 0 n24 ns38 0 -0.00011785218718
Gc12_39 0 n24 ns39 0 0.000129453843313
Gc12_40 0 n24 ns40 0 -0.00010318538896
Gc12_41 0 n24 ns41 0 -0.000640052099338
Gc12_42 0 n24 ns42 0 1.38358711651e-05
Gc12_43 0 n24 ns43 0 -9.48126522045e-05
Gc12_44 0 n24 ns44 0 -0.000152983194766
Gc12_45 0 n24 ns45 0 -0.000114445239096
Gc12_46 0 n24 ns46 0 -4.37858698061e-05
Gc12_47 0 n24 ns47 0 -1.64589791744e-05
Gc12_48 0 n24 ns48 0 -5.8956597428e-05
Gc12_49 0 n24 ns49 0 -3.71484658488e-05
Gc12_50 0 n24 ns50 0 1.19239921646e-06
Gc12_51 0 n24 ns51 0 -6.02747130247e-06
Gc12_52 0 n24 ns52 0 -1.02175138137e-05
Gc12_53 0 n24 ns53 0 -6.17739226687e-06
Gc12_54 0 n24 ns54 0 7.8737526254e-06
Gc12_55 0 n24 ns55 0 -9.3491035228e-07
Gc12_56 0 n24 ns56 0 -4.51265653881e-06
Gc12_57 0 n24 ns57 0 3.21564792954e-06
Gc12_58 0 n24 ns58 0 7.31680437336e-08
Gc12_59 0 n24 ns59 0 2.31976484929e-07
Gc12_60 0 n24 ns60 0 -3.09292155676e-06
Gc12_61 0 n24 ns61 0 -8.90160615925e-07
Gc12_62 0 n24 ns62 0 2.85923054656e-06
Gc12_63 0 n24 ns63 0 1.77014318363e-07
Gc12_64 0 n24 ns64 0 -9.74156757753e-08
Gc12_65 0 n24 ns65 0 -2.49793592217e-05
Gc12_66 0 n24 ns66 0 5.40516314283e-07
Gc12_67 0 n24 ns67 0 -3.14309379312e-06
Gc12_68 0 n24 ns68 0 -6.68313219359e-06
Gc12_69 0 n24 ns69 0 -8.24037559619e-06
Gc12_70 0 n24 ns70 0 -9.10413982197e-07
Gc12_71 0 n24 ns71 0 -1.15451486137e-06
Gc12_72 0 n24 ns72 0 -1.94041204534e-06
Gc12_73 0 n24 ns73 0 -0.000215394845714
Gc12_74 0 n24 ns74 0 4.7261540694e-06
Gc12_75 0 n24 ns75 0 -3.03242023269e-05
Gc12_76 0 n24 ns76 0 -5.47917689852e-05
Gc12_77 0 n24 ns77 0 -5.11803003723e-05
Gc12_78 0 n24 ns78 0 -1.30055756667e-05
Gc12_79 0 n24 ns79 0 -7.48432894173e-06
Gc12_80 0 n24 ns80 0 -1.81064561441e-05
Gc12_81 0 n24 ns81 0 0.000442116787992
Gc12_82 0 n24 ns82 0 -1.01443573133e-05
Gc12_83 0 n24 ns83 0 3.83547234951e-05
Gc12_84 0 n24 ns84 0 5.04203755973e-05
Gc12_85 0 n24 ns85 0 -6.22391668012e-05
Gc12_86 0 n24 ns86 0 -6.44308210856e-05
Gc12_87 0 n24 ns87 0 9.7304023389e-06
Gc12_88 0 n24 ns88 0 1.58972729012e-05
Gc12_89 0 n24 ns89 0 0.00210263191196
Gc12_90 0 n24 ns90 0 -3.45662798555e-05
Gc12_91 0 n24 ns91 0 0.000238262980473
Gc12_92 0 n24 ns92 0 0.0005979504105
Gc12_93 0 n24 ns93 0 8.99621590683e-05
Gc12_94 0 n24 ns94 0 -4.65148045809e-05
Gc12_95 0 n24 ns95 0 -9.48461846857e-05
Gc12_96 0 n24 ns96 0 0.000399396725469
Gc12_97 0 n24 ns97 0 1.60406145504e-05
Gc12_98 0 n24 ns98 0 -5.72203239681e-07
Gc12_99 0 n24 ns99 0 -2.22505051487e-05
Gc12_100 0 n24 ns100 0 -4.78414496104e-05
Gc12_101 0 n24 ns101 0 -8.54177109659e-05
Gc12_102 0 n24 ns102 0 -6.90632814616e-05
Gc12_103 0 n24 ns103 0 4.2598702461e-06
Gc12_104 0 n24 ns104 0 -2.34683894221e-05
Gc12_105 0 n24 ns105 0 -0.000228273047408
Gc12_106 0 n24 ns106 0 5.18469384487e-06
Gc12_107 0 n24 ns107 0 -3.27309473507e-05
Gc12_108 0 n24 ns108 0 -5.20933660223e-05
Gc12_109 0 n24 ns109 0 -4.34633951021e-05
Gc12_110 0 n24 ns110 0 -6.49607632722e-06
Gc12_111 0 n24 ns111 0 -7.1539270336e-06
Gc12_112 0 n24 ns112 0 -1.99755101652e-05
Gc12_113 0 n24 ns113 0 4.66276625029e-05
Gc12_114 0 n24 ns114 0 -7.57751593694e-07
Gc12_115 0 n24 ns115 0 6.05151415499e-06
Gc12_116 0 n24 ns116 0 2.41905797902e-06
Gc12_117 0 n24 ns117 0 4.98379548237e-06
Gc12_118 0 n24 ns118 0 6.13636581096e-06
Gc12_119 0 n24 ns119 0 1.59028475404e-06
Gc12_120 0 n24 ns120 0 3.22243250139e-06
Gc12_121 0 n24 ns121 0 -1.11237243648e-05
Gc12_122 0 n24 ns122 0 2.79959089757e-07
Gc12_123 0 n24 ns123 0 -1.37553880987e-06
Gc12_124 0 n24 ns124 0 -5.60188077136e-06
Gc12_125 0 n24 ns125 0 -5.3899480184e-06
Gc12_126 0 n24 ns126 0 -1.45298456569e-07
Gc12_127 0 n24 ns127 0 -5.57201898676e-07
Gc12_128 0 n24 ns128 0 -8.48493898313e-07
Gd12_1 0 n24 ni1 0 -7.20545335786e-05
Gd12_2 0 n24 ni2 0 -2.82324269035e-05
Gd12_3 0 n24 ni3 0 0.000283446559501
Gd12_4 0 n24 ni4 0 -3.99250798225e-05
Gd12_5 0 n24 ni5 0 0.00239421290958
Gd12_6 0 n24 ni6 0 0.000810857298176
Gd12_7 0 n24 ni7 0 5.84805551825e-05
Gd12_8 0 n24 ni8 0 3.40773102046e-06
Gd12_9 0 n24 ni9 0 2.5381392322e-05
Gd12_10 0 n24 ni10 0 0.000257282980409
Gd12_11 0 n24 ni11 0 -2.77832584681e-05
Gd12_12 0 n24 ni12 0 -0.00131492091039
Gd12_13 0 n24 ni13 0 0.000442301655671
Gd12_14 0 n24 ni14 0 0.000274292104387
Gd12_15 0 n24 ni15 0 -3.7857361774e-05
Gd12_16 0 n24 ni16 0 1.33928222059e-05
Gc13_1 0 n26 ns1 0 -3.20265433397e-06
Gc13_2 0 n26 ns2 0 1.01729570115e-07
Gc13_3 0 n26 ns3 0 -1.13660528189e-07
Gc13_4 0 n26 ns4 0 -5.15790751499e-06
Gc13_5 0 n26 ns5 0 -6.28834330417e-06
Gc13_6 0 n26 ns6 0 -1.50893624818e-07
Gc13_7 0 n26 ns7 0 -4.67872151664e-07
Gc13_8 0 n26 ns8 0 -1.57725381117e-07
Gc13_9 0 n26 ns9 0 3.07376504922e-05
Gc13_10 0 n26 ns10 0 -5.61900590216e-07
Gc13_11 0 n26 ns11 0 4.42595244919e-06
Gc13_12 0 n26 ns12 0 4.81790138288e-07
Gc13_13 0 n26 ns13 0 -8.57540513525e-07
Gc13_14 0 n26 ns14 0 2.45427058053e-06
Gc13_15 0 n26 ns15 0 6.28826906924e-07
Gc13_16 0 n26 ns16 0 2.46635985147e-06
Gc13_17 0 n26 ns17 0 2.82408980511e-05
Gc13_18 0 n26 ns18 0 -3.7441614715e-07
Gc13_19 0 n26 ns19 0 3.67738043991e-06
Gc13_20 0 n26 ns20 0 -6.85504679692e-06
Gc13_21 0 n26 ns21 0 -4.24614979483e-06
Gc13_22 0 n26 ns22 0 2.56667383025e-06
Gc13_23 0 n26 ns23 0 6.93161381618e-07
Gc13_24 0 n26 ns24 0 1.99197980264e-06
Gc13_25 0 n26 ns25 0 -0.000225357024387
Gc13_26 0 n26 ns26 0 4.37159219207e-06
Gc13_27 0 n26 ns27 0 -3.37666355749e-05
Gc13_28 0 n26 ns28 0 -7.20047533642e-05
Gc13_29 0 n26 ns29 0 -8.81755207605e-05
Gc13_30 0 n26 ns30 0 -4.33214105264e-05
Gc13_31 0 n26 ns31 0 -9.6701621047e-06
Gc13_32 0 n26 ns32 0 -1.93393953924e-05
Gc13_33 0 n26 ns33 0 0.00233822841415
Gc13_34 0 n26 ns34 0 -4.63278519359e-05
Gc13_35 0 n26 ns35 0 0.000214754458055
Gc13_36 0 n26 ns36 0 0.000544871474744
Gc13_37 0 n26 ns37 0 7.40170166462e-05
Gc13_38 0 n26 ns38 0 -1.94298070595e-05
Gc13_39 0 n26 ns39 0 4.90021007107e-05
Gc13_40 0 n26 ns40 0 0.00011947861877
Gc13_41 0 n26 ns41 0 0.00132828207303
Gc13_42 0 n26 ns42 0 -1.86033709536e-05
Gc13_43 0 n26 ns43 0 -5.03807738877e-05
Gc13_44 0 n26 ns44 0 0.000256954961272
Gc13_45 0 n26 ns45 0 -2.19729899184e-05
Gc13_46 0 n26 ns46 0 -8.67709110063e-05
Gc13_47 0 n26 ns47 0 7.86687932152e-05
Gc13_48 0 n26 ns48 0 -0.000106804328432
Gc13_49 0 n26 ns49 0 -0.000484216598759
Gc13_50 0 n26 ns50 0 1.02918651775e-05
Gc13_51 0 n26 ns51 0 -7.2965704598e-05
Gc13_52 0 n26 ns52 0 -0.000121637761668
Gc13_53 0 n26 ns53 0 -0.000105129323102
Gc13_54 0 n26 ns54 0 -4.37236830194e-05
Gc13_55 0 n26 ns55 0 -1.33430652445e-05
Gc13_56 0 n26 ns56 0 -4.59131508424e-05
Gc13_57 0 n26 ns57 0 -5.80713728419e-05
Gc13_58 0 n26 ns58 0 1.62707471882e-06
Gc13_59 0 n26 ns59 0 -8.8035330078e-06
Gc13_60 0 n26 ns60 0 -1.3610215698e-05
Gc13_61 0 n26 ns61 0 -9.89053589507e-06
Gc13_62 0 n26 ns62 0 7.05833321937e-06
Gc13_63 0 n26 ns63 0 -1.67633297849e-06
Gc13_64 0 n26 ns64 0 -6.17803511118e-06
Gc13_65 0 n26 ns65 0 1.88210583904e-05
Gc13_66 0 n26 ns66 0 -2.69854602772e-07
Gc13_67 0 n26 ns67 0 2.66949826623e-06
Gc13_68 0 n26 ns68 0 -1.07677517272e-06
Gc13_69 0 n26 ns69 0 -2.10239898931e-06
Gc13_70 0 n26 ns70 0 3.41959928295e-06
Gc13_71 0 n26 ns71 0 3.41659712889e-07
Gc13_72 0 n26 ns72 0 1.18079277049e-06
Gc13_73 0 n26 ns73 0 4.47462542728e-05
Gc13_74 0 n26 ns74 0 -7.25285384624e-07
Gc13_75 0 n26 ns75 0 5.94633949626e-06
Gc13_76 0 n26 ns76 0 3.06074772357e-06
Gc13_77 0 n26 ns77 0 3.33752671339e-06
Gc13_78 0 n26 ns78 0 6.42849685484e-06
Gc13_79 0 n26 ns79 0 1.3036293483e-06
Gc13_80 0 n26 ns80 0 3.08200797288e-06
Gc13_81 0 n26 ns81 0 -0.000190048829312
Gc13_82 0 n26 ns82 0 4.11001605983e-06
Gc13_83 0 n26 ns83 0 -2.66944890208e-05
Gc13_84 0 n26 ns84 0 -5.22496521261e-05
Gc13_85 0 n26 ns85 0 -5.09581626108e-05
Gc13_86 0 n26 ns86 0 -1.49314791451e-05
Gc13_87 0 n26 ns87 0 -6.87506922985e-06
Gc13_88 0 n26 ns88 0 -1.59122708761e-05
Gc13_89 0 n26 ns89 0 1.60406145504e-05
Gc13_90 0 n26 ns90 0 -5.7220323968e-07
Gc13_91 0 n26 ns91 0 -2.22505051487e-05
Gc13_92 0 n26 ns92 0 -4.78414496104e-05
Gc13_93 0 n26 ns93 0 -8.54177109659e-05
Gc13_94 0 n26 ns94 0 -6.90632814616e-05
Gc13_95 0 n26 ns95 0 4.2598702461e-06
Gc13_96 0 n26 ns96 0 -2.34683894221e-05
Gc13_97 0 n26 ns97 0 0.0025469467149
Gc13_98 0 n26 ns98 0 -4.33278185875e-05
Gc13_99 0 n26 ns99 0 0.000261017080668
Gc13_100 0 n26 ns100 0 0.000574315892517
Gc13_101 0 n26 ns101 0 0.000154952677753
Gc13_102 0 n26 ns102 0 -7.67602754687e-05
Gc13_103 0 n26 ns103 0 -5.11098019689e-05
Gc13_104 0 n26 ns104 0 0.000378363617353
Gc13_105 0 n26 ns105 0 5.31578661348e-05
Gc13_106 0 n26 ns106 0 -1.16830536178e-06
Gc13_107 0 n26 ns107 0 -1.82357850945e-05
Gc13_108 0 n26 ns108 0 -2.46139290322e-05
Gc13_109 0 n26 ns109 0 -8.26733788104e-05
Gc13_110 0 n26 ns110 0 -6.1195500916e-05
Gc13_111 0 n26 ns111 0 3.10870055311e-06
Gc13_112 0 n26 ns112 0 -1.99657902181e-05
Gc13_113 0 n26 ns113 0 -0.000208889870213
Gc13_114 0 n26 ns114 0 4.61338535753e-06
Gc13_115 0 n26 ns115 0 -2.95621812087e-05
Gc13_116 0 n26 ns116 0 -5.39493415237e-05
Gc13_117 0 n26 ns117 0 -4.82907398443e-05
Gc13_118 0 n26 ns118 0 -1.21872391384e-05
Gc13_119 0 n26 ns119 0 -7.03765194992e-06
Gc13_120 0 n26 ns120 0 -1.76715311934e-05
Gc13_121 0 n26 ns121 0 4.05970019201e-05
Gc13_122 0 n26 ns122 0 -6.34302000833e-07
Gc13_123 0 n26 ns123 0 5.39799963533e-06
Gc13_124 0 n26 ns124 0 2.24503323336e-06
Gc13_125 0 n26 ns125 0 2.40750278052e-06
Gc13_126 0 n26 ns126 0 6.34026864403e-06
Gc13_127 0 n26 ns127 0 1.13257555334e-06
Gc13_128 0 n26 ns128 0 2.76603721958e-06
Gd13_1 0 n26 ni1 0 3.92471066114e-06
Gd13_2 0 n26 ni2 0 -2.93691804214e-05
Gd13_3 0 n26 ni3 0 -1.45015742586e-05
Gd13_4 0 n26 ni4 0 0.000324198017446
Gd13_5 0 n26 ni5 0 -0.000645710813608
Gd13_6 0 n26 ni6 0 0.0024732842148
Gd13_7 0 n26 ni7 0 0.000645280734517
Gd13_8 0 n26 ni8 0 7.9012564602e-05
Gd13_9 0 n26 ni9 0 -1.52609614812e-05
Gd13_10 0 n26 ni10 0 -3.79931894344e-05
Gd13_11 0 n26 ni11 0 0.00023077462273
Gd13_12 0 n26 ni12 0 0.000442301655671
Gd13_13 0 n26 ni13 0 -0.0011235830978
Gd13_14 0 n26 ni14 0 0.000415939186152
Gd13_15 0 n26 ni15 0 0.000251733576029
Gd13_16 0 n26 ni16 0 -3.37447092617e-05
Gc14_1 0 n28 ns1 0 -1.61502683143e-05
Gc14_2 0 n28 ns2 0 3.42125010003e-07
Gc14_3 0 n28 ns3 0 -1.95785849689e-06
Gc14_4 0 n28 ns4 0 -4.58958248434e-06
Gc14_5 0 n28 ns5 0 -6.11549326171e-06
Gc14_6 0 n28 ns6 0 -7.62966198547e-07
Gc14_7 0 n28 ns7 0 -8.29055558816e-07
Gc14_8 0 n28 ns8 0 -1.19183030654e-06
Gc14_9 0 n28 ns9 0 -1.19920105989e-05
Gc14_10 0 n28 ns10 0 2.61321680393e-07
Gc14_11 0 n28 ns11 0 -1.41279687907e-06
Gc14_12 0 n28 ns12 0 -5.16645518409e-06
Gc14_13 0 n28 ns13 0 -5.55650341292e-06
Gc14_14 0 n28 ns14 0 -9.49498283206e-07
Gc14_15 0 n28 ns15 0 -6.23081541388e-07
Gc14_16 0 n28 ns16 0 -8.14458859871e-07
Gc14_17 0 n28 ns17 0 2.80279685742e-05
Gc14_18 0 n28 ns18 0 -4.93144821695e-07
Gc14_19 0 n28 ns19 0 3.83671043534e-06
Gc14_20 0 n28 ns20 0 -1.36289478433e-06
Gc14_21 0 n28 ns21 0 9.09554492912e-07
Gc14_22 0 n28 ns22 0 1.84427314005e-06
Gc14_23 0 n28 ns23 0 8.92518168504e-07
Gc14_24 0 n28 ns24 0 2.23198932125e-06
Gc14_25 0 n28 ns25 0 1.78065239761e-05
Gc14_26 0 n28 ns26 0 -1.25395336539e-07
Gc14_27 0 n28 ns27 0 2.05102572646e-06
Gc14_28 0 n28 ns28 0 -7.4312727416e-06
Gc14_29 0 n28 ns29 0 -3.66998409759e-06
Gc14_30 0 n28 ns30 0 3.18402644594e-06
Gc14_31 0 n28 ns31 0 5.12260365718e-07
Gc14_32 0 n28 ns32 0 1.01091470225e-06
Gc14_33 0 n28 ns33 0 -0.000203988445157
Gc14_34 0 n28 ns34 0 3.7940735961e-06
Gc14_35 0 n28 ns35 0 -3.0472158993e-05
Gc14_36 0 n28 ns36 0 -7.15652636847e-05
Gc14_37 0 n28 ns37 0 -9.12514232437e-05
Gc14_38 0 n28 ns38 0 -4.75841721521e-05
Gc14_39 0 n28 ns39 0 -9.55089307198e-06
Gc14_40 0 n28 ns40 0 -1.68764038398e-05
Gc14_41 0 n28 ns41 0 0.00149707817867
Gc14_42 0 n28 ns42 0 -2.77376184344e-05
Gc14_43 0 n28 ns43 0 9.56192774145e-05
Gc14_44 0 n28 ns44 0 0.000365635111469
Gc14_45 0 n28 ns45 0 6.29306681561e-06
Gc14_46 0 n28 ns46 0 -3.13979568489e-05
Gc14_47 0 n28 ns47 0 3.55055239812e-05
Gc14_48 0 n28 ns48 0 4.02693941813e-05
Gc14_49 0 n28 ns49 0 0.00137176778548
Gc14_50 0 n28 ns50 0 -1.9904764203e-05
Gc14_51 0 n28 ns51 0 -3.52296360878e-05
Gc14_52 0 n28 ns52 0 0.000272558677495
Gc14_53 0 n28 ns53 0 -1.8018015396e-05
Gc14_54 0 n28 ns54 0 -8.26127163015e-05
Gc14_55 0 n28 ns55 0 7.5050040962e-05
Gc14_56 0 n28 ns56 0 -9.14140787572e-05
Gc14_57 0 n28 ns57 0 -0.000509645790512
Gc14_58 0 n28 ns58 0 1.08935729103e-05
Gc14_59 0 n28 ns59 0 -7.66570916483e-05
Gc14_60 0 n28 ns60 0 -0.000126985881327
Gc14_61 0 n28 ns61 0 -0.000105475676385
Gc14_62 0 n28 ns62 0 -4.23687299047e-05
Gc14_63 0 n28 ns63 0 -1.34163503852e-05
Gc14_64 0 n28 ns64 0 -4.87964106455e-05
Gc14_65 0 n28 ns65 0 -5.03652132962e-07
Gc14_66 0 n28 ns66 0 3.51908736282e-07
Gc14_67 0 n28 ns67 0 -4.39712265447e-07
Gc14_68 0 n28 ns68 0 -6.51743635438e-06
Gc14_69 0 n28 ns69 0 -9.05676342661e-06
Gc14_70 0 n28 ns70 0 7.47567841332e-06
Gc14_71 0 n28 ns71 0 -3.8913972992e-07
Gc14_72 0 n28 ns72 0 -1.57067038167e-06
Gc14_73 0 n28 ns73 0 -6.14856044072e-06
Gc14_74 0 n28 ns74 0 1.77772609317e-07
Gc14_75 0 n28 ns75 0 -7.47838813868e-07
Gc14_76 0 n28 ns76 0 -5.11477848383e-06
Gc14_77 0 n28 ns77 0 -4.07381072025e-06
Gc14_78 0 n28 ns78 0 -7.82809232336e-08
Gc14_79 0 n28 ns79 0 -3.0519607436e-07
Gc14_80 0 n28 ns80 0 -4.54462245249e-07
Gc14_81 0 n28 ns81 0 4.91963294168e-05
Gc14_82 0 n28 ns82 0 -8.28221363194e-07
Gc14_83 0 n28 ns83 0 6.51603091445e-06
Gc14_84 0 n28 ns84 0 2.33706720415e-06
Gc14_85 0 n28 ns85 0 4.10044312229e-06
Gc14_86 0 n28 ns86 0 5.69762813597e-06
Gc14_87 0 n28 ns87 0 1.56609725449e-06
Gc14_88 0 n28 ns88 0 3.50889444873e-06
Gc14_89 0 n28 ns89 0 -0.000228273047408
Gc14_90 0 n28 ns90 0 5.18469384487e-06
Gc14_91 0 n28 ns91 0 -3.27309473507e-05
Gc14_92 0 n28 ns92 0 -5.20933660223e-05
Gc14_93 0 n28 ns93 0 -4.34633951021e-05
Gc14_94 0 n28 ns94 0 -6.49607632722e-06
Gc14_95 0 n28 ns95 0 -7.1539270336e-06
Gc14_96 0 n28 ns96 0 -1.99755101652e-05
Gc14_97 0 n28 ns97 0 5.31578661348e-05
Gc14_98 0 n28 ns98 0 -1.16830536178e-06
Gc14_99 0 n28 ns99 0 -1.82357850945e-05
Gc14_100 0 n28 ns100 0 -2.46139290322e-05
Gc14_101 0 n28 ns101 0 -8.26733788104e-05
Gc14_102 0 n28 ns102 0 -6.1195500916e-05
Gc14_103 0 n28 ns103 0 3.10870055311e-06
Gc14_104 0 n28 ns104 0 -1.99657902181e-05
Gc14_105 0 n28 ns105 0 0.00281894723746
Gc14_106 0 n28 ns106 0 -4.93644563446e-05
Gc14_107 0 n28 ns107 0 0.000296811160772
Gc14_108 0 n28 ns108 0 0.000607382731692
Gc14_109 0 n28 ns109 0 0.000176721858724
Gc14_110 0 n28 ns110 0 -8.52678870904e-05
Gc14_111 0 n28 ns111 0 -4.344757978e-05
Gc14_112 0 n28 ns112 0 0.000400967611515
Gc14_113 0 n28 ns113 0 0.00025016841377
Gc14_114 0 n28 ns114 0 -5.74675438485e-06
Gc14_115 0 n28 ns115 0 1.07226646033e-05
Gc14_116 0 n28 ns116 0 1.17624738297e-05
Gc14_117 0 n28 ns117 0 -7.52572256446e-05
Gc14_118 0 n28 ns118 0 -6.53609569062e-05
Gc14_119 0 n28 ns119 0 5.79820545389e-06
Gc14_120 0 n28 ns120 0 -5.61653505659e-07
Gc14_121 0 n28 ns121 0 -0.00019093895151
Gc14_122 0 n28 ns122 0 4.24002380102e-06
Gc14_123 0 n28 ns123 0 -2.70068504052e-05
Gc14_124 0 n28 ns124 0 -4.96837736737e-05
Gc14_125 0 n28 ns125 0 -4.77757426981e-05
Gc14_126 0 n28 ns126 0 -1.07232690763e-05
Gc14_127 0 n28 ns127 0 -6.77793784536e-06
Gc14_128 0 n28 ns128 0 -1.633912121e-05
Gd14_1 0 n28 ni1 0 1.57662550726e-05
Gd14_2 0 n28 ni2 0 1.24984800771e-05
Gd14_3 0 n28 ni3 0 -2.36829738593e-05
Gd14_4 0 n28 ni4 0 -2.14075632551e-06
Gd14_5 0 n28 ni5 0 0.000300400610231
Gd14_6 0 n28 ni6 0 0.00027836586366
Gd14_7 0 n28 ni7 0 0.00227778946994
Gd14_8 0 n28 ni8 0 0.000673903454497
Gd14_9 0 n28 ni9 0 1.70281693251e-05
Gd14_10 0 n28 ni10 0 8.92046372427e-06
Gd14_11 0 n28 ni11 0 -4.14425446025e-05
Gd14_12 0 n28 ni12 0 0.000274292104387
Gd14_13 0 n28 ni13 0 0.000415939186152
Gd14_14 0 n28 ni14 0 -0.00136811622842
Gd14_15 0 n28 ni15 0 0.000188722757427
Gd14_16 0 n28 ni16 0 0.000232336529133
Gc15_1 0 n30 ns1 0 -3.87286364384e-06
Gc15_2 0 n30 ns2 0 8.98701049763e-08
Gc15_3 0 n30 ns3 0 -4.3163990464e-07
Gc15_4 0 n30 ns4 0 -1.50958242733e-06
Gc15_5 0 n30 ns5 0 -2.20913932122e-06
Gc15_6 0 n30 ns6 0 8.02495980397e-08
Gc15_7 0 n30 ns7 0 -2.61380148037e-07
Gc15_8 0 n30 ns8 0 -2.92972664086e-07
Gc15_9 0 n30 ns9 0 -6.19618196583e-06
Gc15_10 0 n30 ns10 0 1.34841100182e-07
Gc15_11 0 n30 ns11 0 -7.18391090887e-07
Gc15_12 0 n30 ns12 0 -2.45395147122e-06
Gc15_13 0 n30 ns13 0 -2.96452147234e-06
Gc15_14 0 n30 ns14 0 -3.22964885518e-07
Gc15_15 0 n30 ns15 0 -3.47571912745e-07
Gc15_16 0 n30 ns16 0 -4.3294432116e-07
Gc15_17 0 n30 ns17 0 -6.24111369122e-06
Gc15_18 0 n30 ns18 0 1.4587871265e-07
Gc15_19 0 n30 ns19 0 -7.41931778459e-07
Gc15_20 0 n30 ns20 0 -5.71700638605e-06
Gc15_21 0 n30 ns21 0 -3.55787956916e-06
Gc15_22 0 n30 ns22 0 -1.26140224618e-06
Gc15_23 0 n30 ns23 0 -1.92929668152e-07
Gc15_24 0 n30 ns24 0 -3.46911814172e-07
Gc15_25 0 n30 ns25 0 3.03775569146e-05
Gc15_26 0 n30 ns26 0 -5.44309186014e-07
Gc15_27 0 n30 ns27 0 4.19204876073e-06
Gc15_28 0 n30 ns28 0 -8.76958685759e-07
Gc15_29 0 n30 ns29 0 9.41694995034e-07
Gc15_30 0 n30 ns30 0 1.97596118906e-06
Gc15_31 0 n30 ns31 0 9.24058503082e-07
Gc15_32 0 n30 ns32 0 2.4279042646e-06
Gc15_33 0 n30 ns33 0 3.81124211666e-05
Gc15_34 0 n30 ns34 0 -6.06500104008e-07
Gc15_35 0 n30 ns35 0 5.21287235809e-06
Gc15_36 0 n30 ns36 0 -6.59245038961e-06
Gc15_37 0 n30 ns37 0 -4.56097985542e-06
Gc15_38 0 n30 ns38 0 1.95281954917e-06
Gc15_39 0 n30 ns39 0 8.9217208181e-07
Gc15_40 0 n30 ns40 0 2.96175337955e-06
Gc15_41 0 n30 ns41 0 -0.000197644096907
Gc15_42 0 n30 ns42 0 3.71856038516e-06
Gc15_43 0 n30 ns43 0 -2.96761530611e-05
Gc15_44 0 n30 ns44 0 -6.84239109954e-05
Gc15_45 0 n30 ns45 0 -8.72545595793e-05
Gc15_46 0 n30 ns46 0 -4.44639783948e-05
Gc15_47 0 n30 ns47 0 -9.11733947175e-06
Gc15_48 0 n30 ns48 0 -1.67098809391e-05
Gc15_49 0 n30 ns49 0 0.00165839741184
Gc15_50 0 n30 ns50 0 -3.12754648103e-05
Gc15_51 0 n30 ns51 0 0.000119646576834
Gc15_52 0 n30 ns52 0 0.000413688292917
Gc15_53 0 n30 ns53 0 1.10293839642e-05
Gc15_54 0 n30 ns54 0 -2.78062261647e-05
Gc15_55 0 n30 ns55 0 3.400431767e-05
Gc15_56 0 n30 ns56 0 6.01108407528e-05
Gc15_57 0 n30 ns57 0 0.00144473529064
Gc15_58 0 n30 ns58 0 -2.05880173706e-05
Gc15_59 0 n30 ns59 0 -5.54711214874e-05
Gc15_60 0 n30 ns60 0 0.000188893872145
Gc15_61 0 n30 ns61 0 1.04584877974e-05
Gc15_62 0 n30 ns62 0 -0.000114412392334
Gc15_63 0 n30 ns63 0 0.00010295429238
Gc15_64 0 n30 ns64 0 -0.000128225056716
Gc15_65 0 n30 ns65 0 -0.000554674208466
Gc15_66 0 n30 ns66 0 1.188018418e-05
Gc15_67 0 n30 ns67 0 -8.29650683047e-05
Gc15_68 0 n30 ns68 0 -0.000143447072203
Gc15_69 0 n30 ns69 0 -0.000114352221074
Gc15_70 0 n30 ns70 0 -4.40566211289e-05
Gc15_71 0 n30 ns71 0 -1.35817526434e-05
Gc15_72 0 n30 ns72 0 -5.43520905485e-05
Gc15_73 0 n30 ns73 0 -1.21323220079e-05
Gc15_74 0 n30 ns74 0 2.63607267151e-07
Gc15_75 0 n30 ns75 0 -1.52679921289e-06
Gc15_76 0 n30 ns76 0 -4.29227603052e-06
Gc15_77 0 n30 ns77 0 -4.18063444018e-06
Gc15_78 0 n30 ns78 0 -7.67292975811e-07
Gc15_79 0 n30 ns79 0 -5.19017068953e-07
Gc15_80 0 n30 ns80 0 -8.87190430273e-07
Gc15_81 0 n30 ns81 0 3.46770648464e-06
Gc15_82 0 n30 ns82 0 -2.6788672598e-08
Gc15_83 0 n30 ns83 0 5.8011941478e-07
Gc15_84 0 n30 ns84 0 -4.57129846502e-06
Gc15_85 0 n30 ns85 0 -2.7914896606e-06
Gc15_86 0 n30 ns86 0 -1.04224118437e-07
Gc15_87 0 n30 ns87 0 6.42489359127e-08
Gc15_88 0 n30 ns88 0 3.55594397611e-07
Gc15_89 0 n30 ns89 0 4.66276625029e-05
Gc15_90 0 n30 ns90 0 -7.57751593694e-07
Gc15_91 0 n30 ns91 0 6.05151415499e-06
Gc15_92 0 n30 ns92 0 2.41905797902e-06
Gc15_93 0 n30 ns93 0 4.98379548237e-06
Gc15_94 0 n30 ns94 0 6.13636581096e-06
Gc15_95 0 n30 ns95 0 1.59028475404e-06
Gc15_96 0 n30 ns96 0 3.22243250139e-06
Gc15_97 0 n30 ns97 0 -0.000208889870213
Gc15_98 0 n30 ns98 0 4.61338535753e-06
Gc15_99 0 n30 ns99 0 -2.95621812087e-05
Gc15_100 0 n30 ns100 0 -5.39493415237e-05
Gc15_101 0 n30 ns101 0 -4.82907398443e-05
Gc15_102 0 n30 ns102 0 -1.21872391384e-05
Gc15_103 0 n30 ns103 0 -7.03765194992e-06
Gc15_104 0 n30 ns104 0 -1.76715311934e-05
Gc15_105 0 n30 ns105 0 0.00025016841377
Gc15_106 0 n30 ns106 0 -5.74675438485e-06
Gc15_107 0 n30 ns107 0 1.07226646033e-05
Gc15_108 0 n30 ns108 0 1.17624738298e-05
Gc15_109 0 n30 ns109 0 -7.52572256446e-05
Gc15_110 0 n30 ns110 0 -6.53609569062e-05
Gc15_111 0 n30 ns111 0 5.79820545389e-06
Gc15_112 0 n30 ns112 0 -5.61653505657e-07
Gc15_113 0 n30 ns113 0 0.00276250834897
Gc15_114 0 n30 ns114 0 -4.895253666e-05
Gc15_115 0 n30 ns115 0 0.000315005711916
Gc15_116 0 n30 ns116 0 0.000691106004899
Gc15_117 0 n30 ns117 0 0.000147949499178
Gc15_118 0 n30 ns118 0 -5.28501695499e-05
Gc15_119 0 n30 ns119 0 -6.76203404696e-05
Gc15_120 0 n30 ns120 0 0.000430568400451
Gc15_121 0 n30 ns121 0 -8.65359600959e-05
Gc15_122 0 n30 ns122 0 1.87447368562e-06
Gc15_123 0 n30 ns123 0 -3.82167884149e-05
Gc15_124 0 n30 ns124 0 -5.52911282617e-05
Gc15_125 0 n30 ns125 0 -0.000102786248558
Gc15_126 0 n30 ns126 0 -6.66314239375e-05
Gc15_127 0 n30 ns127 0 -1.43666512578e-07
Gc15_128 0 n30 ns128 0 -3.28464651165e-05
Gd15_1 0 n30 ni1 0 3.85756382057e-06
Gd15_2 0 n30 ni2 0 6.23069991758e-06
Gd15_3 0 n30 ni3 0 8.43232800288e-06
Gd15_4 0 n30 ni4 0 -2.65146579729e-05
Gd15_5 0 n30 ni5 0 -2.61303007592e-05
Gd15_6 0 n30 ni6 0 0.000292672877309
Gd15_7 0 n30 ni7 0 8.12469634995e-05
Gd15_8 0 n30 ni8 0 0.00271939044449
Gd15_9 0 n30 ni9 0 0.000728441936391
Gd15_10 0 n30 ni10 0 1.29121964224e-05
Gd15_11 0 n30 ni11 0 -6.65569976706e-07
Gd15_12 0 n30 ni12 0 -3.7857361774e-05
Gd15_13 0 n30 ni13 0 0.000251733576029
Gd15_14 0 n30 ni14 0 0.000188722757427
Gd15_15 0 n30 ni15 0 -0.00175519352731
Gd15_16 0 n30 ni16 0 0.000577771786353
Gc16_1 0 n32 ns1 0 -4.57363747615e-07
Gc16_2 0 n32 ns2 0 2.31169762556e-08
Gc16_3 0 n32 ns3 0 -4.45258905153e-08
Gc16_4 0 n32 ns4 0 -3.66780861288e-07
Gc16_5 0 n32 ns5 0 -6.7277140007e-07
Gc16_6 0 n32 ns6 0 4.58997778174e-07
Gc16_7 0 n32 ns7 0 -7.27149246216e-08
Gc16_8 0 n32 ns8 0 -6.5843443029e-08
Gc16_9 0 n32 ns9 0 -2.51080993227e-06
Gc16_10 0 n32 ns10 0 6.2873687703e-08
Gc16_11 0 n32 ns11 0 -2.83810068169e-07
Gc16_12 0 n32 ns12 0 -4.83521858314e-07
Gc16_13 0 n32 ns13 0 -1.4035843426e-06
Gc16_14 0 n32 ns14 0 3.89496879272e-07
Gc16_15 0 n32 ns15 0 -2.07335119414e-07
Gc16_16 0 n32 ns16 0 -2.12477278762e-07
Gc16_17 0 n32 ns17 0 -6.61507577058e-06
Gc16_18 0 n32 ns18 0 1.44858704987e-07
Gc16_19 0 n32 ns19 0 -7.81728229064e-07
Gc16_20 0 n32 ns20 0 -2.43268002078e-06
Gc16_21 0 n32 ns21 0 -2.96651042326e-06
Gc16_22 0 n32 ns22 0 -2.80914841197e-07
Gc16_23 0 n32 ns23 0 -3.61299282375e-07
Gc16_24 0 n32 ns24 0 -4.72741089205e-07
Gc16_25 0 n32 ns25 0 -1.33757747242e-05
Gc16_26 0 n32 ns26 0 2.90673759896e-07
Gc16_27 0 n32 ns27 0 -1.58852394086e-06
Gc16_28 0 n32 ns28 0 -5.104172281e-06
Gc16_29 0 n32 ns29 0 -5.90425640655e-06
Gc16_30 0 n32 ns30 0 -8.75761924157e-07
Gc16_31 0 n32 ns31 0 -7.06633272464e-07
Gc16_32 0 n32 ns32 0 -9.30544897281e-07
Gc16_33 0 n32 ns33 0 3.36720091403e-05
Gc16_34 0 n32 ns34 0 -6.24253823121e-07
Gc16_35 0 n32 ns35 0 4.86138862183e-06
Gc16_36 0 n32 ns36 0 9.45181086767e-07
Gc16_37 0 n32 ns37 0 -7.84318096147e-07
Gc16_38 0 n32 ns38 0 2.58471141307e-06
Gc16_39 0 n32 ns39 0 6.76330586715e-07
Gc16_40 0 n32 ns40 0 2.72312753278e-06
Gc16_41 0 n32 ns41 0 2.49742273719e-05
Gc16_42 0 n32 ns42 0 -3.0343412114e-07
Gc16_43 0 n32 ns43 0 3.28404612067e-06
Gc16_44 0 n32 ns44 0 -6.65294054959e-06
Gc16_45 0 n32 ns45 0 -5.68851717827e-06
Gc16_46 0 n32 ns46 0 2.88112556534e-06
Gc16_47 0 n32 ns47 0 4.36333198941e-07
Gc16_48 0 n32 ns48 0 1.67218921582e-06
Gc16_49 0 n32 ns49 0 -0.000256580224924
Gc16_50 0 n32 ns50 0 5.11243805401e-06
Gc16_51 0 n32 ns51 0 -3.79884825281e-05
Gc16_52 0 n32 ns52 0 -7.55284999659e-05
Gc16_53 0 n32 ns53 0 -9.15406838338e-05
Gc16_54 0 n32 ns54 0 -4.07896820163e-05
Gc16_55 0 n32 ns55 0 -1.05721660025e-05
Gc16_56 0 n32 ns56 0 -2.23556028986e-05
Gc16_57 0 n32 ns57 0 0.00174499801323
Gc16_58 0 n32 ns58 0 -3.3215408067e-05
Gc16_59 0 n32 ns59 0 0.000130973727851
Gc16_60 0 n32 ns60 0 0.000449511823642
Gc16_61 0 n32 ns61 0 -3.95091382586e-06
Gc16_62 0 n32 ns62 0 -2.86444539224e-05
Gc16_63 0 n32 ns63 0 3.08449940804e-05
Gc16_64 0 n32 ns64 0 6.94405872255e-05
Gc16_65 0 n32 ns65 0 0.00234877905334
Gc16_66 0 n32 ns66 0 -4.17321968383e-05
Gc16_67 0 n32 ns67 0 7.28214005941e-05
Gc16_68 0 n32 ns68 0 0.000252875440643
Gc16_69 0 n32 ns69 0 9.52922970868e-05
Gc16_70 0 n32 ns70 0 -0.000147858583895
Gc16_71 0 n32 ns71 0 0.000139262885025
Gc16_72 0 n32 ns72 0 -6.09760253552e-05
Gc16_73 0 n32 ns73 0 -6.7935037963e-06
Gc16_74 0 n32 ns74 0 1.51215699355e-07
Gc16_75 0 n32 ns75 0 -8.21800021607e-07
Gc16_76 0 n32 ns76 0 -1.08234753819e-06
Gc16_77 0 n32 ns77 0 -2.62261287762e-06
Gc16_78 0 n32 ns78 0 2.64589779324e-07
Gc16_79 0 n32 ns79 0 -4.23445235459e-07
Gc16_80 0 n32 ns80 0 -5.4146526617e-07
Gc16_81 0 n32 ns81 0 -1.56385244704e-05
Gc16_82 0 n32 ns82 0 3.32252237804e-07
Gc16_83 0 n32 ns83 0 -1.91200169939e-06
Gc16_84 0 n32 ns84 0 -4.03261200512e-06
Gc16_85 0 n32 ns85 0 -5.66003742796e-06
Gc16_86 0 n32 ns86 0 -6.18188926581e-07
Gc16_87 0 n32 ns87 0 -8.07335886215e-07
Gc16_88 0 n32 ns88 0 -1.1585456105e-06
Gc16_89 0 n32 ns89 0 -1.11237243648e-05
Gc16_90 0 n32 ns90 0 2.79959089757e-07
Gc16_91 0 n32 ns91 0 -1.37553880987e-06
Gc16_92 0 n32 ns92 0 -5.60188077136e-06
Gc16_93 0 n32 ns93 0 -5.3899480184e-06
Gc16_94 0 n32 ns94 0 -1.45298456569e-07
Gc16_95 0 n32 ns95 0 -5.57201898676e-07
Gc16_96 0 n32 ns96 0 -8.48493898313e-07
Gc16_97 0 n32 ns97 0 4.05970019201e-05
Gc16_98 0 n32 ns98 0 -6.34302000833e-07
Gc16_99 0 n32 ns99 0 5.39799963533e-06
Gc16_100 0 n32 ns100 0 2.24503323336e-06
Gc16_101 0 n32 ns101 0 2.40750278052e-06
Gc16_102 0 n32 ns102 0 6.34026864403e-06
Gc16_103 0 n32 ns103 0 1.13257555334e-06
Gc16_104 0 n32 ns104 0 2.76603721958e-06
Gc16_105 0 n32 ns105 0 -0.00019093895151
Gc16_106 0 n32 ns106 0 4.24002380102e-06
Gc16_107 0 n32 ns107 0 -2.70068504052e-05
Gc16_108 0 n32 ns108 0 -4.96837736737e-05
Gc16_109 0 n32 ns109 0 -4.77757426981e-05
Gc16_110 0 n32 ns110 0 -1.07232690763e-05
Gc16_111 0 n32 ns111 0 -6.77793784536e-06
Gc16_112 0 n32 ns112 0 -1.633912121e-05
Gc16_113 0 n32 ns113 0 -8.65359600959e-05
Gc16_114 0 n32 ns114 0 1.87447368562e-06
Gc16_115 0 n32 ns115 0 -3.82167884149e-05
Gc16_116 0 n32 ns116 0 -5.52911282617e-05
Gc16_117 0 n32 ns117 0 -0.000102786248558
Gc16_118 0 n32 ns118 0 -6.66314239375e-05
Gc16_119 0 n32 ns119 0 -1.43666512579e-07
Gc16_120 0 n32 ns120 0 -3.28464651165e-05
Gc16_121 0 n32 ns121 0 0.00282249924087
Gc16_122 0 n32 ns122 0 -5.05484740722e-05
Gc16_123 0 n32 ns123 0 0.000325218471957
Gc16_124 0 n32 ns124 0 0.000771010954176
Gc16_125 0 n32 ns125 0 0.000101627014436
Gc16_126 0 n32 ns126 0 -4.6150936829e-05
Gc16_127 0 n32 ns127 0 -8.00632257186e-05
Gc16_128 0 n32 ns128 0 0.000441381778948
Gd16_1 0 n32 ni1 0 7.68098493696e-07
Gd16_2 0 n32 ni2 0 2.35642833709e-06
Gd16_3 0 n32 ni3 0 6.69100849414e-06
Gd16_4 0 n32 ni4 0 1.36673536186e-05
Gd16_5 0 n32 ni5 0 -3.27183378631e-05
Gd16_6 0 n32 ni6 0 -1.17284404978e-05
Gd16_7 0 n32 ni7 0 0.000354792270976
Gd16_8 0 n32 ni8 0 5.70965984879e-06
Gd16_9 0 n32 ni9 0 0.0017656377046
Gd16_10 0 n32 ni10 0 6.30326646412e-06
Gd16_11 0 n32 ni11 0 1.51900969614e-05
Gd16_12 0 n32 ni12 0 1.33928222059e-05
Gd16_13 0 n32 ni13 0 -3.37447092617e-05
Gd16_14 0 n32 ni14 0 0.000232336529133
Gd16_15 0 n32 ni15 0 0.000577771786353
Gd16_16 0 n32 ni16 0 -0.00185055972006
Gc17_129 0 n34 ns129 0 0.00443033184969
Gc17_130 0 n34 ns130 0 -8.53987184957e-05
Gc17_131 0 n34 ns131 0 0.000513583097002
Gc17_132 0 n34 ns132 0 0.000887926660691
Gc17_133 0 n34 ns133 0 0.000298967663366
Gc17_134 0 n34 ns134 0 -8.38898663078e-05
Gc17_135 0 n34 ns135 0 8.08483507646e-07
Gc17_136 0 n34 ns136 0 0.000520141047351
Gc17_137 0 n34 ns137 0 0.00197538164282
Gc17_138 0 n34 ns138 0 -3.38766779844e-05
Gc17_139 0 n34 ns139 0 4.27405051916e-05
Gc17_140 0 n34 ns140 0 0.000327267498887
Gc17_141 0 n34 ns141 0 1.27742523074e-05
Gc17_142 0 n34 ns142 0 -0.000112985473158
Gc17_143 0 n34 ns143 0 9.76066802375e-05
Gc17_144 0 n34 ns144 0 -5.34835783035e-05
Gc17_145 0 n34 ns145 0 -0.00052107230389
Gc17_146 0 n34 ns146 0 1.09531391784e-05
Gc17_147 0 n34 ns147 0 -7.74932498464e-05
Gc17_148 0 n34 ns148 0 -0.000135459896804
Gc17_149 0 n34 ns149 0 -0.000123470489552
Gc17_150 0 n34 ns150 0 -5.03518660533e-05
Gc17_151 0 n34 ns151 0 -1.5020583969e-05
Gc17_152 0 n34 ns152 0 -4.91949074398e-05
Gc17_153 0 n34 ns153 0 7.30196924656e-06
Gc17_154 0 n34 ns154 0 2.26492507689e-07
Gc17_155 0 n34 ns155 0 4.78812895107e-07
Gc17_156 0 n34 ns156 0 -6.60905021238e-06
Gc17_157 0 n34 ns157 0 -5.55830646295e-06
Gc17_158 0 n34 ns158 0 8.05618558295e-06
Gc17_159 0 n34 ns159 0 1.21803573774e-07
Gc17_160 0 n34 ns160 0 -7.92775181765e-07
Gc17_161 0 n34 ns161 0 1.35656372589e-05
Gc17_162 0 n34 ns162 0 -1.55764943396e-07
Gc17_163 0 n34 ns163 0 1.91771962977e-06
Gc17_164 0 n34 ns164 0 -1.52519381556e-06
Gc17_165 0 n34 ns165 0 -2.59970023172e-06
Gc17_166 0 n34 ns166 0 3.38282693512e-06
Gc17_167 0 n34 ns167 0 1.65053867196e-07
Gc17_168 0 n34 ns168 0 7.53025738557e-07
Gc17_169 0 n34 ns169 0 -3.06050536826e-05
Gc17_170 0 n34 ns170 0 6.60081195375e-07
Gc17_171 0 n34 ns171 0 -3.91670304776e-06
Gc17_172 0 n34 ns172 0 -7.07286218715e-06
Gc17_173 0 n34 ns173 0 -9.00732037322e-06
Gc17_174 0 n34 ns174 0 -9.24992987795e-07
Gc17_175 0 n34 ns175 0 -1.36981950601e-06
Gc17_176 0 n34 ns176 0 -2.40553908227e-06
Gc17_177 0 n34 ns177 0 -1.47916828061e-05
Gc17_178 0 n34 ns178 0 3.12076773426e-07
Gc17_179 0 n34 ns179 0 -1.77396695398e-06
Gc17_180 0 n34 ns180 0 -2.72953712497e-06
Gc17_181 0 n34 ns181 0 -5.5532784192e-06
Gc17_182 0 n34 ns182 0 -1.57461685514e-07
Gc17_183 0 n34 ns183 0 -8.5981085107e-07
Gc17_184 0 n34 ns184 0 -1.13303185558e-06
Gc17_185 0 n34 ns185 0 -1.25620906464e-06
Gc17_186 0 n34 ns186 0 4.08974149788e-08
Gc17_187 0 n34 ns187 0 -1.60982709195e-07
Gc17_188 0 n34 ns188 0 -9.16825760851e-07
Gc17_189 0 n34 ns189 0 -8.07864029922e-07
Gc17_190 0 n34 ns190 0 2.94648591741e-07
Gc17_191 0 n34 ns191 0 -6.87981632436e-08
Gc17_192 0 n34 ns192 0 -1.24079376585e-07
Gc17_193 0 n34 ns193 0 1.67725608497e-06
Gc17_194 0 n34 ns194 0 -1.89545011707e-08
Gc17_195 0 n34 ns195 0 2.08393457017e-07
Gc17_196 0 n34 ns196 0 -3.97220728029e-07
Gc17_197 0 n34 ns197 0 2.6606856596e-08
Gc17_198 0 n34 ns198 0 4.58268492725e-07
Gc17_199 0 n34 ns199 0 7.09971356125e-08
Gc17_200 0 n34 ns200 0 9.4965052511e-08
Gc17_201 0 n34 ns201 0 0.000310054649495
Gc17_202 0 n34 ns202 0 -7.5790263544e-06
Gc17_203 0 n34 ns203 0 1.94747088505e-05
Gc17_204 0 n34 ns204 0 -1.95408506006e-06
Gc17_205 0 n34 ns205 0 -9.17915853797e-05
Gc17_206 0 n34 ns206 0 -8.37137922697e-05
Gc17_207 0 n34 ns207 0 8.83866439149e-06
Gc17_208 0 n34 ns208 0 1.52706257142e-06
Gc17_209 0 n34 ns209 0 -0.000182158362103
Gc17_210 0 n34 ns210 0 4.02845363093e-06
Gc17_211 0 n34 ns211 0 -2.55371836663e-05
Gc17_212 0 n34 ns212 0 -4.97734747553e-05
Gc17_213 0 n34 ns213 0 -5.17000566399e-05
Gc17_214 0 n34 ns214 0 -1.10632181189e-05
Gc17_215 0 n34 ns215 0 -6.80721247628e-06
Gc17_216 0 n34 ns216 0 -1.58904781004e-05
Gc17_217 0 n34 ns217 0 7.733002638e-05
Gc17_218 0 n34 ns218 0 -1.42954198782e-06
Gc17_219 0 n34 ns219 0 1.07058650543e-05
Gc17_220 0 n34 ns220 0 6.19313766866e-06
Gc17_221 0 n34 ns221 0 4.05951133347e-06
Gc17_222 0 n34 ns222 0 6.9131254031e-06
Gc17_223 0 n34 ns223 0 2.07944567914e-06
Gc17_224 0 n34 ns224 0 5.76371935762e-06
Gc17_225 0 n34 ns225 0 4.9081659875e-06
Gc17_226 0 n34 ns226 0 -7.3050743847e-08
Gc17_227 0 n34 ns227 0 1.0356195598e-06
Gc17_228 0 n34 ns228 0 -4.51008781946e-06
Gc17_229 0 n34 ns229 0 -5.52285259528e-06
Gc17_230 0 n34 ns230 0 -1.29066089474e-07
Gc17_231 0 n34 ns231 0 -2.06717282931e-07
Gc17_232 0 n34 ns232 0 5.30744237983e-07
Gc17_233 0 n34 ns233 0 -1.69827161015e-05
Gc17_234 0 n34 ns234 0 3.59693814167e-07
Gc17_235 0 n34 ns235 0 -2.06151375346e-06
Gc17_236 0 n34 ns236 0 -4.41115606647e-06
Gc17_237 0 n34 ns237 0 -6.33549784162e-06
Gc17_238 0 n34 ns238 0 -6.60134767694e-07
Gc17_239 0 n34 ns239 0 -8.87678411229e-07
Gc17_240 0 n34 ns240 0 -1.27264896543e-06
Gc17_241 0 n34 ns241 0 -4.40896228817e-06
Gc17_242 0 n34 ns242 0 1.01540444749e-07
Gc17_243 0 n34 ns243 0 -5.04656543256e-07
Gc17_244 0 n34 ns244 0 -1.45244153256e-06
Gc17_245 0 n34 ns245 0 -2.28280679221e-06
Gc17_246 0 n34 ns246 0 1.22043923387e-07
Gc17_247 0 n34 ns247 0 -2.88582963005e-07
Gc17_248 0 n34 ns248 0 -3.41532995247e-07
Gc17_249 0 n34 ns249 0 5.47928584666e-08
Gc17_250 0 n34 ns250 0 1.23386166374e-08
Gc17_251 0 n34 ns251 0 1.87981375548e-08
Gc17_252 0 n34 ns252 0 -4.08227354013e-07
Gc17_253 0 n34 ns253 0 -5.29882634366e-07
Gc17_254 0 n34 ns254 0 4.24206541947e-07
Gc17_255 0 n34 ns255 0 -3.83760312087e-08
Gc17_256 0 n34 ns256 0 -2.36854284737e-08
Gd17_17 0 n34 ni17 0 -0.00292685887431
Gd17_18 0 n34 ni18 0 0.00177323231406
Gd17_19 0 n34 ni19 0 0.000685464803364
Gd17_20 0 n34 ni20 0 1.08444607516e-05
Gd17_21 0 n34 ni21 0 -9.64707390168e-06
Gd17_22 0 n34 ni22 0 3.09789765259e-05
Gd17_23 0 n34 ni23 0 1.34367946382e-05
Gd17_24 0 n34 ni24 0 1.91103853184e-06
Gd17_25 0 n34 ni25 0 -8.50607552001e-07
Gd17_26 0 n34 ni26 0 0.000139649861222
Gd17_27 0 n34 ni27 0 0.000222617609962
Gd17_28 0 n34 ni28 0 -7.31066984986e-05
Gd17_29 0 n34 ni29 0 -4.53758675177e-06
Gd17_30 0 n34 ni30 0 1.63795167917e-05
Gd17_31 0 n34 ni31 0 4.33983755983e-06
Gd17_32 0 n34 ni32 0 3.63182731526e-07
Gc18_129 0 n36 ns129 0 0.00197538164282
Gc18_130 0 n36 ns130 0 -3.38766779844e-05
Gc18_131 0 n36 ns131 0 4.27405051916e-05
Gc18_132 0 n36 ns132 0 0.000327267498887
Gc18_133 0 n36 ns133 0 1.27742523074e-05
Gc18_134 0 n36 ns134 0 -0.000112985473158
Gc18_135 0 n36 ns135 0 9.76066802375e-05
Gc18_136 0 n36 ns136 0 -5.34835783035e-05
Gc18_137 0 n36 ns137 0 0.00254605031782
Gc18_138 0 n36 ns138 0 -4.35452111609e-05
Gc18_139 0 n36 ns139 0 0.000260505239421
Gc18_140 0 n36 ns140 0 0.000604037708165
Gc18_141 0 n36 ns141 0 0.000119437019521
Gc18_142 0 n36 ns142 0 -7.83216495984e-05
Gc18_143 0 n36 ns143 0 -5.72402819756e-05
Gc18_144 0 n36 ns144 0 0.000377730845551
Gc18_145 0 n36 ns145 0 0.000113102852201
Gc18_146 0 n36 ns146 0 -2.61172163164e-06
Gc18_147 0 n36 ns147 0 -9.02201734479e-06
Gc18_148 0 n36 ns148 0 -1.2936376485e-05
Gc18_149 0 n36 ns149 0 -8.51461922694e-05
Gc18_150 0 n36 ns150 0 -6.26976309827e-05
Gc18_151 0 n36 ns151 0 3.52651246227e-06
Gc18_152 0 n36 ns152 0 -1.43076603524e-05
Gc18_153 0 n36 ns153 0 -0.000184758348528
Gc18_154 0 n36 ns154 0 4.11199442709e-06
Gc18_155 0 n36 ns155 0 -2.6203230319e-05
Gc18_156 0 n36 ns156 0 -4.98301491456e-05
Gc18_157 0 n36 ns157 0 -4.58661913378e-05
Gc18_158 0 n36 ns158 0 -1.10049878198e-05
Gc18_159 0 n36 ns159 0 -6.43795470912e-06
Gc18_160 0 n36 ns160 0 -1.56814799145e-05
Gc18_161 0 n36 ns161 0 3.53594576079e-05
Gc18_162 0 n36 ns162 0 -5.206497634e-07
Gc18_163 0 n36 ns163 0 4.64485168624e-06
Gc18_164 0 n36 ns164 0 2.38236722006e-06
Gc18_165 0 n36 ns165 0 1.93305676145e-06
Gc18_166 0 n36 ns166 0 6.57900395022e-06
Gc18_167 0 n36 ns167 0 9.42378552506e-07
Gc18_168 0 n36 ns168 0 2.26078242009e-06
Gc18_169 0 n36 ns169 0 -1.71945529931e-05
Gc18_170 0 n36 ns170 0 4.07382377781e-07
Gc18_171 0 n36 ns171 0 -2.2089364016e-06
Gc18_172 0 n36 ns172 0 -5.9138010829e-06
Gc18_173 0 n36 ns173 0 -6.2668396593e-06
Gc18_174 0 n36 ns174 0 -1.42431326888e-07
Gc18_175 0 n36 ns175 0 -7.92191301715e-07
Gc18_176 0 n36 ns176 0 -1.37370821033e-06
Gc18_177 0 n36 ns177 0 -1.50620155548e-05
Gc18_178 0 n36 ns178 0 3.19179100052e-07
Gc18_179 0 n36 ns179 0 -1.82797677892e-06
Gc18_180 0 n36 ns180 0 -4.00163507526e-06
Gc18_181 0 n36 ns181 0 -5.62410315084e-06
Gc18_182 0 n36 ns182 0 -6.3835544089e-07
Gc18_183 0 n36 ns183 0 -7.89271096538e-07
Gc18_184 0 n36 ns184 0 -1.10776446439e-06
Gc18_185 0 n36 ns185 0 -3.30015529186e-06
Gc18_186 0 n36 ns186 0 8.08517218538e-08
Gc18_187 0 n36 ns187 0 -4.1069396312e-07
Gc18_188 0 n36 ns188 0 -1.43027707199e-06
Gc18_189 0 n36 ns189 0 -1.4633355967e-06
Gc18_190 0 n36 ns190 0 7.52478281486e-08
Gc18_191 0 n36 ns191 0 -1.65319921253e-07
Gc18_192 0 n36 ns192 0 -2.61099207903e-07
Gc18_193 0 n36 ns193 0 1.14100323904e-10
Gc18_194 0 n36 ns194 0 1.31414501056e-08
Gc18_195 0 n36 ns195 0 1.66909831802e-08
Gc18_196 0 n36 ns196 0 -3.93996171683e-07
Gc18_197 0 n36 ns197 0 -5.95047448575e-07
Gc18_198 0 n36 ns198 0 4.29406188071e-07
Gc18_199 0 n36 ns199 0 -4.8404230285e-08
Gc18_200 0 n36 ns200 0 -2.71601396184e-08
Gc18_201 0 n36 ns201 0 0.00178206886175
Gc18_202 0 n36 ns202 0 -3.40637084719e-05
Gc18_203 0 n36 ns203 0 0.000135569811946
Gc18_204 0 n36 ns204 0 0.000416849249638
Gc18_205 0 n36 ns205 0 2.44606450996e-05
Gc18_206 0 n36 ns206 0 -3.22037957035e-05
Gc18_207 0 n36 ns207 0 4.05626890389e-05
Gc18_208 0 n36 ns208 0 6.66321845711e-05
Gc18_209 0 n36 ns209 0 -0.000267174996208
Gc18_210 0 n36 ns210 0 5.3447858213e-06
Gc18_211 0 n36 ns211 0 -3.94151121682e-05
Gc18_212 0 n36 ns212 0 -7.5982279035e-05
Gc18_213 0 n36 ns213 0 -9.31847931764e-05
Gc18_214 0 n36 ns214 0 -4.10644691591e-05
Gc18_215 0 n36 ns215 0 -1.12262584765e-05
Gc18_216 0 n36 ns216 0 -2.27800045622e-05
Gc18_217 0 n36 ns217 0 3.32870787667e-05
Gc18_218 0 n36 ns218 0 -5.00182165155e-07
Gc18_219 0 n36 ns219 0 4.54448540439e-06
Gc18_220 0 n36 ns220 0 -6.23033590648e-06
Gc18_221 0 n36 ns221 0 -5.70600452125e-06
Gc18_222 0 n36 ns222 0 2.33656965896e-06
Gc18_223 0 n36 ns223 0 6.18588789146e-07
Gc18_224 0 n36 ns224 0 2.48166174707e-06
Gc18_225 0 n36 ns225 0 3.79524285912e-05
Gc18_226 0 n36 ns226 0 -7.1416073835e-07
Gc18_227 0 n36 ns227 0 5.43240328863e-06
Gc18_228 0 n36 ns228 0 1.10493777751e-06
Gc18_229 0 n36 ns229 0 -1.3867833371e-08
Gc18_230 0 n36 ns230 0 2.55301134937e-06
Gc18_231 0 n36 ns231 0 8.72325500788e-07
Gc18_232 0 n36 ns232 0 3.07434730433e-06
Gc18_233 0 n36 ns233 0 -1.33355424201e-05
Gc18_234 0 n36 ns234 0 2.91817450727e-07
Gc18_235 0 n36 ns235 0 -1.60742569852e-06
Gc18_236 0 n36 ns236 0 -5.08720653946e-06
Gc18_237 0 n36 ns237 0 -5.64978307588e-06
Gc18_238 0 n36 ns238 0 -8.36443791649e-07
Gc18_239 0 n36 ns239 0 -6.7268816613e-07
Gc18_240 0 n36 ns240 0 -9.47913571328e-07
Gc18_241 0 n36 ns241 0 -6.21514766582e-06
Gc18_242 0 n36 ns242 0 1.36817946084e-07
Gc18_243 0 n36 ns243 0 -7.33781561121e-07
Gc18_244 0 n36 ns244 0 -2.38815207263e-06
Gc18_245 0 n36 ns245 0 -2.83567387845e-06
Gc18_246 0 n36 ns246 0 -2.699612921e-07
Gc18_247 0 n36 ns247 0 -3.37327672664e-07
Gc18_248 0 n36 ns248 0 -4.44846641079e-07
Gc18_249 0 n36 ns249 0 -1.57066795593e-06
Gc18_250 0 n36 ns250 0 4.35766279547e-08
Gc18_251 0 n36 ns251 0 -1.70641176063e-07
Gc18_252 0 n36 ns252 0 -5.68180280887e-07
Gc18_253 0 n36 ns253 0 -1.11537023788e-06
Gc18_254 0 n36 ns254 0 3.34263086421e-07
Gc18_255 0 n36 ns255 0 -1.40862230092e-07
Gc18_256 0 n36 ns256 0 -1.36606983246e-07
Gd18_17 0 n36 ni17 0 0.00177323231406
Gd18_18 0 n36 ni18 0 -0.00111091602565
Gd18_19 0 n36 ni19 0 0.000342607412087
Gd18_20 0 n36 ni20 0 0.000226568444921
Gd18_21 0 n36 ni21 0 -2.83614667589e-05
Gd18_22 0 n36 ni22 0 1.93801761121e-05
Gd18_23 0 n36 ni23 0 1.45647470786e-05
Gd18_24 0 n36 ni24 0 3.81327801596e-06
Gd18_25 0 n36 ni25 0 3.55350447338e-07
Gd18_26 0 n36 ni26 0 -2.12815643512e-05
Gd18_27 0 n36 ni27 0 0.000364881563081
Gd18_28 0 n36 ni28 0 -2.12523804366e-05
Gd18_29 0 n36 ni29 0 -3.67400193527e-05
Gd18_30 0 n36 ni30 0 1.38752198232e-05
Gd18_31 0 n36 ni31 0 6.35537833744e-06
Gd18_32 0 n36 ni32 0 1.65374822263e-06
Gc19_129 0 n38 ns129 0 -0.00052107230389
Gc19_130 0 n38 ns130 0 1.09531391784e-05
Gc19_131 0 n38 ns131 0 -7.74932498464e-05
Gc19_132 0 n38 ns132 0 -0.000135459896804
Gc19_133 0 n38 ns133 0 -0.000123470489552
Gc19_134 0 n38 ns134 0 -5.03518660533e-05
Gc19_135 0 n38 ns135 0 -1.5020583969e-05
Gc19_136 0 n38 ns136 0 -4.91949074398e-05
Gc19_137 0 n38 ns137 0 0.000113102852201
Gc19_138 0 n38 ns138 0 -2.61172163164e-06
Gc19_139 0 n38 ns139 0 -9.0220173448e-06
Gc19_140 0 n38 ns140 0 -1.2936376485e-05
Gc19_141 0 n38 ns141 0 -8.51461922694e-05
Gc19_142 0 n38 ns142 0 -6.26976309827e-05
Gc19_143 0 n38 ns143 0 3.52651246226e-06
Gc19_144 0 n38 ns144 0 -1.43076603524e-05
Gc19_145 0 n38 ns145 0 0.00249144406448
Gc19_146 0 n38 ns146 0 -4.19295944993e-05
Gc19_147 0 n38 ns147 0 0.000250599840449
Gc19_148 0 n38 ns148 0 0.000533653501263
Gc19_149 0 n38 ns149 0 0.000163977305428
Gc19_150 0 n38 ns150 0 -8.34235104616e-05
Gc19_151 0 n38 ns151 0 -4.69844576307e-05
Gc19_152 0 n38 ns152 0 0.000369931919853
Gc19_153 0 n38 ns153 0 0.00027547942249
Gc19_154 0 n38 ns154 0 -6.29743904079e-06
Gc19_155 0 n38 ns155 0 1.52662861889e-05
Gc19_156 0 n38 ns156 0 2.01455865057e-05
Gc19_157 0 n38 ns157 0 -7.13739157615e-05
Gc19_158 0 n38 ns158 0 -6.28060102586e-05
Gc19_159 0 n38 ns159 0 5.57531817177e-06
Gc19_160 0 n38 ns160 0 3.28812347368e-06
Gc19_161 0 n38 ns161 0 -0.000243806168314
Gc19_162 0 n38 ns162 0 5.42528677548e-06
Gc19_163 0 n38 ns163 0 -3.45521665106e-05
Gc19_164 0 n38 ns164 0 -5.68681852698e-05
Gc19_165 0 n38 ns165 0 -5.00437543758e-05
Gc19_166 0 n38 ns166 0 -1.02474333421e-05
Gc19_167 0 n38 ns167 0 -7.95365907297e-06
Gc19_168 0 n38 ns168 0 -2.08947327703e-05
Gc19_169 0 n38 ns169 0 3.59291539627e-05
Gc19_170 0 n38 ns170 0 -5.17275241691e-07
Gc19_171 0 n38 ns171 0 4.52266992836e-06
Gc19_172 0 n38 ns172 0 2.59033604094e-06
Gc19_173 0 n38 ns173 0 4.17125174957e-06
Gc19_174 0 n38 ns174 0 6.85511135141e-06
Gc19_175 0 n38 ns175 0 1.21378701607e-06
Gc19_176 0 n38 ns176 0 2.19875271132e-06
Gc19_177 0 n38 ns177 0 4.41802438122e-06
Gc19_178 0 n38 ns178 0 -4.89953204648e-08
Gc19_179 0 n38 ns179 0 7.48482092281e-07
Gc19_180 0 n38 ns180 0 -4.04150364066e-06
Gc19_181 0 n38 ns181 0 -3.0161971271e-06
Gc19_182 0 n38 ns182 0 5.65313466912e-08
Gc19_183 0 n38 ns183 0 2.48215745122e-08
Gc19_184 0 n38 ns184 0 4.33779109321e-07
Gc19_185 0 n38 ns185 0 -1.0728648796e-05
Gc19_186 0 n38 ns186 0 2.36920505096e-07
Gc19_187 0 n38 ns187 0 -1.37831665325e-06
Gc19_188 0 n38 ns188 0 -4.46597855045e-06
Gc19_189 0 n38 ns189 0 -3.54116510808e-06
Gc19_190 0 n38 ns190 0 -8.31523477795e-07
Gc19_191 0 n38 ns191 0 -3.92367661306e-07
Gc19_192 0 n38 ns192 0 -7.81671188253e-07
Gc19_193 0 n38 ns193 0 -5.16237636419e-06
Gc19_194 0 n38 ns194 0 1.15175557401e-07
Gc19_195 0 n38 ns195 0 -5.79125061106e-07
Gc19_196 0 n38 ns196 0 -1.38421003863e-06
Gc19_197 0 n38 ns197 0 -2.67882728836e-06
Gc19_198 0 n38 ns198 0 1.36255822705e-07
Gc19_199 0 n38 ns199 0 -3.60297080737e-07
Gc19_200 0 n38 ns200 0 -3.95732490212e-07
Gc19_201 0 n38 ns201 0 0.00127287147905
Gc19_202 0 n38 ns202 0 -1.70232403006e-05
Gc19_203 0 n38 ns203 0 -6.09795598044e-05
Gc19_204 0 n38 ns204 0 0.000267415140037
Gc19_205 0 n38 ns205 0 -3.50050203318e-05
Gc19_206 0 n38 ns206 0 -8.29567995603e-05
Gc19_207 0 n38 ns207 0 7.31693981773e-05
Gc19_208 0 n38 ns208 0 -0.000109603359805
Gc19_209 0 n38 ns209 0 0.00166906749824
Gc19_210 0 n38 ns210 0 -3.15684708875e-05
Gc19_211 0 n38 ns211 0 0.000122405720945
Gc19_212 0 n38 ns212 0 0.000417289081472
Gc19_213 0 n38 ns213 0 1.90010912889e-05
Gc19_214 0 n38 ns214 0 -2.18361121753e-05
Gc19_215 0 n38 ns215 0 3.58491100484e-05
Gc19_216 0 n38 ns216 0 5.92064875233e-05
Gc19_217 0 n38 ns217 0 -0.00017177073103
Gc19_218 0 n38 ns218 0 3.03997583428e-06
Gc19_219 0 n38 ns219 0 -2.5688780132e-05
Gc19_220 0 n38 ns220 0 -6.60011769802e-05
Gc19_221 0 n38 ns221 0 -8.99652185167e-05
Gc19_222 0 n38 ns222 0 -4.82944389287e-05
Gc19_223 0 n38 ns223 0 -9.03026798271e-06
Gc19_224 0 n38 ns224 0 -1.37709351205e-05
Gc19_225 0 n38 ns225 0 3.84017844558e-05
Gc19_226 0 n38 ns226 0 -6.21160805768e-07
Gc19_227 0 n38 ns227 0 5.29937603072e-06
Gc19_228 0 n38 ns228 0 -7.1009321353e-06
Gc19_229 0 n38 ns229 0 -5.09336172222e-06
Gc19_230 0 n38 ns230 0 1.553232906e-06
Gc19_231 0 n38 ns231 0 8.77393960938e-07
Gc19_232 0 n38 ns232 0 3.03333521248e-06
Gc19_233 0 n38 ns233 0 2.60666358716e-05
Gc19_234 0 n38 ns234 0 -4.51887875034e-07
Gc19_235 0 n38 ns235 0 3.58886350753e-06
Gc19_236 0 n38 ns236 0 -1.08883575176e-06
Gc19_237 0 n38 ns237 0 4.3894775372e-07
Gc19_238 0 n38 ns238 0 2.0404767572e-06
Gc19_239 0 n38 ns239 0 7.75710499288e-07
Gc19_240 0 n38 ns240 0 2.03417517817e-06
Gc19_241 0 n38 ns241 0 -7.87620638845e-06
Gc19_242 0 n38 ns242 0 1.79741965036e-07
Gc19_243 0 n38 ns243 0 -9.4776889781e-07
Gc19_244 0 n38 ns244 0 -5.50734435248e-06
Gc19_245 0 n38 ns245 0 -3.96035923335e-06
Gc19_246 0 n38 ns246 0 -1.14493889138e-06
Gc19_247 0 n38 ns247 0 -2.98283274329e-07
Gc19_248 0 n38 ns248 0 -4.90177944627e-07
Gc19_249 0 n38 ns249 0 -7.00660133042e-06
Gc19_250 0 n38 ns250 0 1.5167016135e-07
Gc19_251 0 n38 ns251 0 -8.20297489284e-07
Gc19_252 0 n38 ns252 0 -2.35232568451e-06
Gc19_253 0 n38 ns253 0 -3.1640734489e-06
Gc19_254 0 n38 ns254 0 -2.66343538937e-07
Gc19_255 0 n38 ns255 0 -4.00116692533e-07
Gc19_256 0 n38 ns256 0 -5.02843839907e-07
Gd19_17 0 n38 ni17 0 0.000685464803364
Gd19_18 0 n38 ni18 0 0.000342607412087
Gd19_19 0 n38 ni19 0 -0.00101587046647
Gd19_20 0 n38 ni20 0 0.000143379554203
Gd19_21 0 n38 ni21 0 0.000288419473067
Gd19_22 0 n38 ni22 0 -2.69957025158e-05
Gd19_23 0 n38 ni23 0 -2.22104834109e-06
Gd19_24 0 n38 ni24 0 1.21001062324e-05
Gd19_25 0 n38 ni25 0 4.73051916026e-06
Gd19_26 0 n38 ni26 0 0.00257494590141
Gd19_27 0 n38 ni27 0 4.47447586163e-05
Gd19_28 0 n38 ni28 0 0.000262585654946
Gd19_29 0 n38 ni29 0 -2.66429824283e-05
Gd19_30 0 n38 ni30 0 -2.21435560549e-05
Gd19_31 0 n38 ni31 0 9.71314523216e-06
Gd19_32 0 n38 ni32 0 6.86507352528e-06
Gc20_129 0 n40 ns129 0 7.30196924656e-06
Gc20_130 0 n40 ns130 0 2.26492507689e-07
Gc20_131 0 n40 ns131 0 4.78812895108e-07
Gc20_132 0 n40 ns132 0 -6.60905021238e-06
Gc20_133 0 n40 ns133 0 -5.55830646295e-06
Gc20_134 0 n40 ns134 0 8.05618558295e-06
Gc20_135 0 n40 ns135 0 1.21803573774e-07
Gc20_136 0 n40 ns136 0 -7.92775181765e-07
Gc20_137 0 n40 ns137 0 -0.000184758348528
Gc20_138 0 n40 ns138 0 4.11199442709e-06
Gc20_139 0 n40 ns139 0 -2.6203230319e-05
Gc20_140 0 n40 ns140 0 -4.98301491456e-05
Gc20_141 0 n40 ns141 0 -4.58661913378e-05
Gc20_142 0 n40 ns142 0 -1.10049878198e-05
Gc20_143 0 n40 ns143 0 -6.43795470912e-06
Gc20_144 0 n40 ns144 0 -1.56814799145e-05
Gc20_145 0 n40 ns145 0 0.00027547942249
Gc20_146 0 n40 ns146 0 -6.29743904079e-06
Gc20_147 0 n40 ns147 0 1.52662861889e-05
Gc20_148 0 n40 ns148 0 2.01455865057e-05
Gc20_149 0 n40 ns149 0 -7.13739157615e-05
Gc20_150 0 n40 ns150 0 -6.28060102586e-05
Gc20_151 0 n40 ns151 0 5.57531817178e-06
Gc20_152 0 n40 ns152 0 3.28812347368e-06
Gc20_153 0 n40 ns153 0 0.0024572540604
Gc20_154 0 n40 ns154 0 -4.0459220001e-05
Gc20_155 0 n40 ns155 0 0.000221395085557
Gc20_156 0 n40 ns156 0 0.000490730578254
Gc20_157 0 n40 ns157 0 0.000149198354389
Gc20_158 0 n40 ns158 0 -0.000109132557453
Gc20_159 0 n40 ns159 0 -3.61241046186e-05
Gc20_160 0 n40 ns160 0 0.000338292800983
Gc20_161 0 n40 ns161 0 -0.000119041320448
Gc20_162 0 n40 ns162 0 2.72638953624e-06
Gc20_163 0 n40 ns163 0 -4.40067390766e-05
Gc20_164 0 n40 ns164 0 -6.97532768023e-05
Gc20_165 0 n40 ns165 0 -9.10102852696e-05
Gc20_166 0 n40 ns166 0 -6.4947936202e-05
Gc20_167 0 n40 ns167 0 2.22791825878e-06
Gc20_168 0 n40 ns168 0 -3.78747576339e-05
Gc20_169 0 n40 ns169 0 -0.000276443662959
Gc20_170 0 n40 ns170 0 6.38875514535e-06
Gc20_171 0 n40 ns171 0 -3.98279121712e-05
Gc20_172 0 n40 ns172 0 -5.63517492063e-05
Gc20_173 0 n40 ns173 0 -4.12273649965e-05
Gc20_174 0 n40 ns174 0 -1.21031662736e-06
Gc20_175 0 n40 ns175 0 -7.84964740317e-06
Gc20_176 0 n40 ns176 0 -2.47619898646e-05
Gc20_177 0 n40 ns177 0 5.17091479984e-05
Gc20_178 0 n40 ns178 0 -8.82283467562e-07
Gc20_179 0 n40 ns179 0 6.80720005299e-06
Gc20_180 0 n40 ns180 0 1.78669389651e-06
Gc20_181 0 n40 ns181 0 4.97113112419e-06
Gc20_182 0 n40 ns182 0 5.34172995064e-06
Gc20_183 0 n40 ns183 0 1.77878004493e-06
Gc20_184 0 n40 ns184 0 3.72902072723e-06
Gc20_185 0 n40 ns185 0 -5.38563464307e-06
Gc20_186 0 n40 ns186 0 1.7010665414e-07
Gc20_187 0 n40 ns187 0 -7.84867720737e-07
Gc20_188 0 n40 ns188 0 -6.40379803217e-06
Gc20_189 0 n40 ns189 0 -2.54063903107e-06
Gc20_190 0 n40 ns190 0 -4.99140861372e-07
Gc20_191 0 n40 ns191 0 -8.31991487463e-09
Gc20_192 0 n40 ns192 0 -4.06454994006e-07
Gc20_193 0 n40 ns193 0 -1.29585490452e-05
Gc20_194 0 n40 ns194 0 2.78515819321e-07
Gc20_195 0 n40 ns195 0 -1.59040419369e-06
Gc20_196 0 n40 ns196 0 -4.93828053284e-06
Gc20_197 0 n40 ns197 0 -4.97049521728e-06
Gc20_198 0 n40 ns198 0 -9.34367104711e-07
Gc20_199 0 n40 ns199 0 -5.80137857788e-07
Gc20_200 0 n40 ns200 0 -9.40202246415e-07
Gc20_201 0 n40 ns201 0 -0.000508213037802
Gc20_202 0 n40 ns202 0 1.08195802248e-05
Gc20_203 0 n40 ns203 0 -7.58612447122e-05
Gc20_204 0 n40 ns204 0 -0.000126150320067
Gc20_205 0 n40 ns205 0 -0.00010990400649
Gc20_206 0 n40 ns206 0 -4.52722846055e-05
Gc20_207 0 n40 ns207 0 -1.48603195403e-05
Gc20_208 0 n40 ns208 0 -4.63364501973e-05
Gc20_209 0 n40 ns209 0 0.00130887914861
Gc20_210 0 n40 ns210 0 -1.8676172166e-05
Gc20_211 0 n40 ns211 0 -3.47104426868e-05
Gc20_212 0 n40 ns212 0 0.000290435613173
Gc20_213 0 n40 ns213 0 -2.68253148113e-05
Gc20_214 0 n40 ns214 0 -7.24735164399e-05
Gc20_215 0 n40 ns215 0 6.49422394252e-05
Gc20_216 0 n40 ns216 0 -8.1551587668e-05
Gc20_217 0 n40 ns217 0 0.00156320061994
Gc20_218 0 n40 ns218 0 -2.93045088013e-05
Gc20_219 0 n40 ns219 0 0.000109309459108
Gc20_220 0 n40 ns220 0 0.000391708020177
Gc20_221 0 n40 ns221 0 8.39797280059e-06
Gc20_222 0 n40 ns222 0 -2.70096610872e-05
Gc20_223 0 n40 ns223 0 3.25200382389e-05
Gc20_224 0 n40 ns224 0 5.36158478825e-05
Gc20_225 0 n40 ns225 0 -0.000170186034785
Gc20_226 0 n40 ns226 0 3.03358613983e-06
Gc20_227 0 n40 ns227 0 -2.58088438595e-05
Gc20_228 0 n40 ns228 0 -6.8780230585e-05
Gc20_229 0 n40 ns229 0 -8.72485474163e-05
Gc20_230 0 n40 ns230 0 -4.85698399507e-05
Gc20_231 0 n40 ns231 0 -8.30723890537e-06
Gc20_232 0 n40 ns232 0 -1.40684582433e-05
Gc20_233 0 n40 ns233 0 1.06417417816e-05
Gc20_234 0 n40 ns234 0 4.49536344769e-08
Gc20_235 0 n40 ns235 0 8.87549088776e-07
Gc20_236 0 n40 ns236 0 -7.92784942294e-06
Gc20_237 0 n40 ns237 0 -2.86039764916e-06
Gc20_238 0 n40 ns238 0 3.62068457176e-06
Gc20_239 0 n40 ns239 0 4.89944621164e-07
Gc20_240 0 n40 ns240 0 2.27252652544e-07
Gc20_241 0 n40 ns241 0 2.41720982126e-05
Gc20_242 0 n40 ns242 0 -4.07348547403e-07
Gc20_243 0 n40 ns243 0 3.21228125022e-06
Gc20_244 0 n40 ns244 0 -2.60139744367e-06
Gc20_245 0 n40 ns245 0 1.30438576621e-06
Gc20_246 0 n40 ns246 0 1.48443556621e-06
Gc20_247 0 n40 ns247 0 9.30459771362e-07
Gc20_248 0 n40 ns248 0 1.89943721576e-06
Gc20_249 0 n40 ns249 0 -1.00470253424e-05
Gc20_250 0 n40 ns250 0 2.26299914288e-07
Gc20_251 0 n40 ns251 0 -1.23212275319e-06
Gc20_252 0 n40 ns252 0 -5.53469931986e-06
Gc20_253 0 n40 ns253 0 -4.41550244487e-06
Gc20_254 0 n40 ns254 0 -1.05923420368e-06
Gc20_255 0 n40 ns255 0 -4.07754826767e-07
Gc20_256 0 n40 ns256 0 -6.7638426384e-07
Gd20_17 0 n40 ni17 0 1.08444607516e-05
Gd20_18 0 n40 ni18 0 0.000226568444921
Gd20_19 0 n40 ni19 0 0.000143379554203
Gd20_20 0 n40 ni20 0 -0.000564979949688
Gd20_21 0 n40 ni21 0 0.000628164002486
Gd20_22 0 n40 ni22 0 0.000326244483298
Gd20_23 0 n40 ni23 0 -4.30734856707e-05
Gd20_24 0 n40 ni24 0 1.02280488526e-05
Gd20_25 0 n40 ni25 0 1.35884040403e-05
Gd20_26 0 n40 ni26 0 0.000665020699165
Gd20_27 0 n40 ni27 0 0.00218462950339
Gd20_28 0 n40 ni28 0 0.000133009848401
Gd20_29 0 n40 ni29 0 0.000266384621423
Gd20_30 0 n40 ni30 0 6.88572029591e-06
Gd20_31 0 n40 ni31 0 -1.84350154855e-05
Gd20_32 0 n40 ni32 0 1.1690764446e-05
Gc21_129 0 n42 ns129 0 1.35656372589e-05
Gc21_130 0 n42 ns130 0 -1.55764943396e-07
Gc21_131 0 n42 ns131 0 1.91771962977e-06
Gc21_132 0 n42 ns132 0 -1.52519381556e-06
Gc21_133 0 n42 ns133 0 -2.59970023172e-06
Gc21_134 0 n42 ns134 0 3.38282693512e-06
Gc21_135 0 n42 ns135 0 1.65053867196e-07
Gc21_136 0 n42 ns136 0 7.53025738557e-07
Gc21_137 0 n42 ns137 0 3.53594576079e-05
Gc21_138 0 n42 ns138 0 -5.206497634e-07
Gc21_139 0 n42 ns139 0 4.64485168624e-06
Gc21_140 0 n42 ns140 0 2.38236722006e-06
Gc21_141 0 n42 ns141 0 1.93305676145e-06
Gc21_142 0 n42 ns142 0 6.57900395022e-06
Gc21_143 0 n42 ns143 0 9.42378552506e-07
Gc21_144 0 n42 ns144 0 2.26078242009e-06
Gc21_145 0 n42 ns145 0 -0.000243806168314
Gc21_146 0 n42 ns146 0 5.42528677548e-06
Gc21_147 0 n42 ns147 0 -3.45521665106e-05
Gc21_148 0 n42 ns148 0 -5.68681852698e-05
Gc21_149 0 n42 ns149 0 -5.00437543758e-05
Gc21_150 0 n42 ns150 0 -1.02474333421e-05
Gc21_151 0 n42 ns151 0 -7.95365907297e-06
Gc21_152 0 n42 ns152 0 -2.08947327703e-05
Gc21_153 0 n42 ns153 0 -0.000119041320448
Gc21_154 0 n42 ns154 0 2.72638953624e-06
Gc21_155 0 n42 ns155 0 -4.40067390766e-05
Gc21_156 0 n42 ns156 0 -6.97532768023e-05
Gc21_157 0 n42 ns157 0 -9.10102852696e-05
Gc21_158 0 n42 ns158 0 -6.4947936202e-05
Gc21_159 0 n42 ns159 0 2.22791825878e-06
Gc21_160 0 n42 ns160 0 -3.78747576339e-05
Gc21_161 0 n42 ns161 0 0.00172172114502
Gc21_162 0 n42 ns162 0 -2.6499236605e-05
Gc21_163 0 n42 ns163 0 0.000191290459621
Gc21_164 0 n42 ns164 0 0.000550391788158
Gc21_165 0 n42 ns165 0 4.93026521333e-05
Gc21_166 0 n42 ns166 0 -4.02652266577e-05
Gc21_167 0 n42 ns167 0 -0.000106733143589
Gc21_168 0 n42 ns168 0 0.000369682696091
Gc21_169 0 n42 ns169 0 -4.57559205108e-05
Gc21_170 0 n42 ns170 0 7.67095408912e-07
Gc21_171 0 n42 ns171 0 -3.37241918926e-05
Gc21_172 0 n42 ns172 0 -7.9743616577e-05
Gc21_173 0 n42 ns173 0 -8.58979938445e-05
Gc21_174 0 n42 ns174 0 -7.56112191811e-05
Gc21_175 0 n42 ns175 0 7.92636106253e-06
Gc21_176 0 n42 ns176 0 -3.54730129274e-05
Gc21_177 0 n42 ns177 0 -0.000157891414269
Gc21_178 0 n42 ns178 0 3.308961004e-06
Gc21_179 0 n42 ns179 0 -2.1950177423e-05
Gc21_180 0 n42 ns180 0 -4.96536090927e-05
Gc21_181 0 n42 ns181 0 -5.23795027206e-05
Gc21_182 0 n42 ns182 0 -1.81648417013e-05
Gc21_183 0 n42 ns183 0 -6.29681737742e-06
Gc21_184 0 n42 ns184 0 -1.29235588521e-05
Gc21_185 0 n42 ns185 0 4.98858490247e-05
Gc21_186 0 n42 ns186 0 -8.41613722655e-07
Gc21_187 0 n42 ns187 0 6.67519611143e-06
Gc21_188 0 n42 ns188 0 2.85917292361e-06
Gc21_189 0 n42 ns189 0 3.77290856164e-06
Gc21_190 0 n42 ns190 0 6.04942341069e-06
Gc21_191 0 n42 ns191 0 1.51283826448e-06
Gc21_192 0 n42 ns192 0 3.54572171625e-06
Gc21_193 0 n42 ns193 0 3.07314839005e-06
Gc21_194 0 n42 ns194 0 -3.63272599161e-08
Gc21_195 0 n42 ns195 0 8.08308920139e-07
Gc21_196 0 n42 ns196 0 -4.29492203614e-06
Gc21_197 0 n42 ns197 0 -6.0311872348e-06
Gc21_198 0 n42 ns198 0 -3.37206458522e-08
Gc21_199 0 n42 ns199 0 -3.27225691668e-07
Gc21_200 0 n42 ns200 0 3.68825479228e-07
Gc21_201 0 n42 ns201 0 -6.17816254036e-05
Gc21_202 0 n42 ns202 0 1.74986330091e-06
Gc21_203 0 n42 ns203 0 -9.40333936283e-06
Gc21_204 0 n42 ns204 0 -1.34449001868e-05
Gc21_205 0 n42 ns205 0 -8.54082041553e-06
Gc21_206 0 n42 ns206 0 8.35419128121e-06
Gc21_207 0 n42 ns207 0 -1.70450106561e-06
Gc21_208 0 n42 ns208 0 -6.49632100499e-06
Gc21_209 0 n42 ns209 0 -0.000531780502685
Gc21_210 0 n42 ns210 0 1.13471956681e-05
Gc21_211 0 n42 ns211 0 -7.97480222113e-05
Gc21_212 0 n42 ns212 0 -0.000129903300348
Gc21_213 0 n42 ns213 0 -0.000109889199387
Gc21_214 0 n42 ns214 0 -4.42226622106e-05
Gc21_215 0 n42 ns215 0 -1.4473930927e-05
Gc21_216 0 n42 ns216 0 -5.0179212223e-05
Gc21_217 0 n42 ns217 0 0.00199390528219
Gc21_218 0 n42 ns218 0 -3.21546787817e-05
Gc21_219 0 n42 ns219 0 3.61632466146e-06
Gc21_220 0 n42 ns220 0 0.000264246952066
Gc21_221 0 n42 ns221 0 6.7218883078e-05
Gc21_222 0 n42 ns222 0 -0.000119199496022
Gc21_223 0 n42 ns223 0 0.000126839976001
Gc21_224 0 n42 ns224 0 -0.000104421539545
Gc21_225 0 n42 ns225 0 0.00285122941534
Gc21_226 0 n42 ns226 0 -5.76952618647e-05
Gc21_227 0 n42 ns227 0 0.000287364733151
Gc21_228 0 n42 ns228 0 0.000666227611578
Gc21_229 0 n42 ns229 0 0.000107110229529
Gc21_230 0 n42 ns230 0 -1.04027360321e-05
Gc21_231 0 n42 ns231 0 5.52341999835e-05
Gc21_232 0 n42 ns232 0 0.000167912032143
Gc21_233 0 n42 ns233 0 -0.000173215164082
Gc21_234 0 n42 ns234 0 3.18960499216e-06
Gc21_235 0 n42 ns235 0 -2.6785850694e-05
Gc21_236 0 n42 ns236 0 -6.44675872247e-05
Gc21_237 0 n42 ns237 0 -8.34645613861e-05
Gc21_238 0 n42 ns238 0 -4.36229344444e-05
Gc21_239 0 n42 ns239 0 -7.80898851309e-06
Gc21_240 0 n42 ns240 0 -1.59229212503e-05
Gc21_241 0 n42 ns241 0 3.18982930675e-05
Gc21_242 0 n42 ns242 0 -4.60668994107e-07
Gc21_243 0 n42 ns243 0 4.2504089657e-06
Gc21_244 0 n42 ns244 0 -6.23127892136e-06
Gc21_245 0 n42 ns245 0 -4.47765563216e-06
Gc21_246 0 n42 ns246 0 2.56348621427e-06
Gc21_247 0 n42 ns247 0 7.30172313007e-07
Gc21_248 0 n42 ns248 0 2.30131295973e-06
Gc21_249 0 n42 ns249 0 3.35154064557e-05
Gc21_250 0 n42 ns250 0 -6.2324267438e-07
Gc21_251 0 n42 ns251 0 4.8413698426e-06
Gc21_252 0 n42 ns252 0 8.80982103684e-07
Gc21_253 0 n42 ns253 0 -8.10236164991e-07
Gc21_254 0 n42 ns254 0 2.51543216331e-06
Gc21_255 0 n42 ns255 0 6.82198892097e-07
Gc21_256 0 n42 ns256 0 2.70054115857e-06
Gd21_17 0 n42 ni17 0 -9.64707390169e-06
Gd21_18 0 n42 ni18 0 -2.83614667589e-05
Gd21_19 0 n42 ni19 0 0.000288419473067
Gd21_20 0 n42 ni20 0 0.000628164002486
Gd21_21 0 n42 ni21 0 -0.00101848957804
Gd21_22 0 n42 ni22 0 0.000558945010528
Gd21_23 0 n42 ni23 0 0.000196085987071
Gd21_24 0 n42 ni24 0 -4.3100061764e-05
Gd21_25 0 n42 ni25 0 -3.12519358751e-06
Gd21_26 0 n42 ni26 0 8.31518675384e-05
Gd21_27 0 n42 ni27 0 0.000697977125634
Gd21_28 0 n42 ni28 0 0.00242730950401
Gd21_29 0 n42 ni29 0 -0.00120936735797
Gd21_30 0 n42 ni30 0 0.000274444029911
Gd21_31 0 n42 ni31 0 -1.90454185308e-05
Gd21_32 0 n42 ni32 0 -3.25757267317e-05
Gc22_129 0 n44 ns129 0 -3.06050536826e-05
Gc22_130 0 n44 ns130 0 6.60081195375e-07
Gc22_131 0 n44 ns131 0 -3.91670304776e-06
Gc22_132 0 n44 ns132 0 -7.07286218715e-06
Gc22_133 0 n44 ns133 0 -9.00732037322e-06
Gc22_134 0 n44 ns134 0 -9.24992987795e-07
Gc22_135 0 n44 ns135 0 -1.36981950601e-06
Gc22_136 0 n44 ns136 0 -2.40553908227e-06
Gc22_137 0 n44 ns137 0 -1.71945529931e-05
Gc22_138 0 n44 ns138 0 4.07382377781e-07
Gc22_139 0 n44 ns139 0 -2.2089364016e-06
Gc22_140 0 n44 ns140 0 -5.9138010829e-06
Gc22_141 0 n44 ns141 0 -6.2668396593e-06
Gc22_142 0 n44 ns142 0 -1.42431326888e-07
Gc22_143 0 n44 ns143 0 -7.92191301715e-07
Gc22_144 0 n44 ns144 0 -1.37370821033e-06
Gc22_145 0 n44 ns145 0 3.59291539627e-05
Gc22_146 0 n44 ns146 0 -5.17275241691e-07
Gc22_147 0 n44 ns147 0 4.52266992836e-06
Gc22_148 0 n44 ns148 0 2.59033604094e-06
Gc22_149 0 n44 ns149 0 4.17125174957e-06
Gc22_150 0 n44 ns150 0 6.85511135141e-06
Gc22_151 0 n44 ns151 0 1.21378701607e-06
Gc22_152 0 n44 ns152 0 2.19875271132e-06
Gc22_153 0 n44 ns153 0 -0.000276443662959
Gc22_154 0 n44 ns154 0 6.38875514535e-06
Gc22_155 0 n44 ns155 0 -3.98279121712e-05
Gc22_156 0 n44 ns156 0 -5.63517492063e-05
Gc22_157 0 n44 ns157 0 -4.12273649965e-05
Gc22_158 0 n44 ns158 0 -1.21031662736e-06
Gc22_159 0 n44 ns159 0 -7.84964740317e-06
Gc22_160 0 n44 ns160 0 -2.47619898646e-05
Gc22_161 0 n44 ns161 0 -4.57559205108e-05
Gc22_162 0 n44 ns162 0 7.67095408912e-07
Gc22_163 0 n44 ns163 0 -3.37241918926e-05
Gc22_164 0 n44 ns164 0 -7.9743616577e-05
Gc22_165 0 n44 ns165 0 -8.58979938445e-05
Gc22_166 0 n44 ns166 0 -7.56112191811e-05
Gc22_167 0 n44 ns167 0 7.92636106253e-06
Gc22_168 0 n44 ns168 0 -3.54730129274e-05
Gc22_169 0 n44 ns169 0 0.00192156903433
Gc22_170 0 n44 ns170 0 -3.09374637099e-05
Gc22_171 0 n44 ns171 0 0.000239213753323
Gc22_172 0 n44 ns172 0 0.00071055823856
Gc22_173 0 n44 ns173 0 3.33686949114e-05
Gc22_174 0 n44 ns174 0 -4.00385782472e-06
Gc22_175 0 n44 ns175 0 -0.000134033973809
Gc22_176 0 n44 ns176 0 0.000430244761039
Gc22_177 0 n44 ns177 0 0.000702153706474
Gc22_178 0 n44 ns178 0 -1.60958182142e-05
Gc22_179 0 n44 ns179 0 7.61809351702e-05
Gc22_180 0 n44 ns180 0 0.000111084049443
Gc22_181 0 n44 ns181 0 -5.3667063409e-05
Gc22_182 0 n44 ns182 0 -6.50788150424e-05
Gc22_183 0 n44 ns183 0 1.17854112503e-05
Gc22_184 0 n44 ns184 0 4.17672609415e-05
Gc22_185 0 n44 ns185 0 -0.000169376832916
Gc22_186 0 n44 ns186 0 3.61064851698e-06
Gc22_187 0 n44 ns187 0 -2.36873422387e-05
Gc22_188 0 n44 ns188 0 -5.1580872406e-05
Gc22_189 0 n44 ns189 0 -5.08619738567e-05
Gc22_190 0 n44 ns190 0 -1.71329139902e-05
Gc22_191 0 n44 ns191 0 -6.40293377735e-06
Gc22_192 0 n44 ns192 0 -1.3810386846e-05
Gc22_193 0 n44 ns193 0 9.7323880913e-05
Gc22_194 0 n44 ns194 0 -1.87183261737e-06
Gc22_195 0 n44 ns195 0 1.36542410049e-05
Gc22_196 0 n44 ns196 0 9.18009403794e-06
Gc22_197 0 n44 ns197 0 4.7664335293e-06
Gc22_198 0 n44 ns198 0 7.21042618057e-06
Gc22_199 0 n44 ns199 0 2.47540795848e-06
Gc22_200 0 n44 ns200 0 7.49728276233e-06
Gc22_201 0 n44 ns201 0 -2.44664340862e-07
Gc22_202 0 n44 ns202 0 1.53022803091e-07
Gc22_203 0 n44 ns203 0 -2.87421576414e-07
Gc22_204 0 n44 ns204 0 -3.07995996449e-06
Gc22_205 0 n44 ns205 0 -8.6899931677e-07
Gc22_206 0 n44 ns206 0 3.0667550508e-06
Gc22_207 0 n44 ns207 0 7.73937785179e-08
Gc22_208 0 n44 ns208 0 -4.05074848322e-07
Gc22_209 0 n44 ns209 0 -4.4516484898e-05
Gc22_210 0 n44 ns210 0 1.37551926006e-06
Gc22_211 0 n44 ns211 0 -7.07019150765e-06
Gc22_212 0 n44 ns212 0 -8.3552148196e-06
Gc22_213 0 n44 ns213 0 -6.42900882486e-06
Gc22_214 0 n44 ns214 0 9.65652119655e-06
Gc22_215 0 n44 ns215 0 -1.27291011538e-06
Gc22_216 0 n44 ns216 0 -5.36127815906e-06
Gc22_217 0 n44 ns217 0 -0.00094957645976
Gc22_218 0 n44 ns218 0 2.08885327754e-05
Gc22_219 0 n44 ns219 0 -0.000138802811919
Gc22_220 0 n44 ns220 0 -0.000214130955143
Gc22_221 0 n44 ns221 0 -0.000130656649253
Gc22_222 0 n44 ns222 0 -4.17738721932e-05
Gc22_223 0 n44 ns223 0 -2.16205792165e-05
Gc22_224 0 n44 ns224 0 -8.70011645526e-05
Gc22_225 0 n44 ns225 0 0.00253107630446
Gc22_226 0 n44 ns226 0 -4.3690007843e-05
Gc22_227 0 n44 ns227 0 5.36737371871e-05
Gc22_228 0 n44 ns228 0 0.000227173564971
Gc22_229 0 n44 ns229 0 0.000157374025965
Gc22_230 0 n44 ns230 0 -0.000152362149267
Gc22_231 0 n44 ns231 0 0.000173429951137
Gc22_232 0 n44 ns232 0 -0.000104104854591
Gc22_233 0 n44 ns233 0 0.00200150135913
Gc22_234 0 n44 ns234 0 -3.90851185788e-05
Gc22_235 0 n44 ns235 0 0.000170772526484
Gc22_236 0 n44 ns236 0 0.000491206869421
Gc22_237 0 n44 ns237 0 4.18926906033e-05
Gc22_238 0 n44 ns238 0 -1.7047538038e-05
Gc22_239 0 n44 ns239 0 4.09461375119e-05
Gc22_240 0 n44 ns240 0 9.01416772668e-05
Gc22_241 0 n44 ns241 0 -0.000155117365667
Gc22_242 0 n44 ns242 0 2.60999310966e-06
Gc22_243 0 n44 ns243 0 -2.32484571994e-05
Gc22_244 0 n44 ns244 0 -6.53841012324e-05
Gc22_245 0 n44 ns245 0 -9.18139425139e-05
Gc22_246 0 n44 ns246 0 -5.12667348643e-05
Gc22_247 0 n44 ns247 0 -8.92727097601e-06
Gc22_248 0 n44 ns248 0 -1.18666599177e-05
Gc22_249 0 n44 ns249 0 4.67361772516e-05
Gc22_250 0 n44 ns250 0 -8.39908711039e-07
Gc22_251 0 n44 ns251 0 6.66103360451e-06
Gc22_252 0 n44 ns252 0 -5.51356213722e-06
Gc22_253 0 n44 ns253 0 -7.21231675159e-06
Gc22_254 0 n44 ns254 0 8.62277580491e-07
Gc22_255 0 n44 ns255 0 7.54105666793e-07
Gc22_256 0 n44 ns256 0 3.84090475125e-06
Gd22_17 0 n44 ni17 0 3.09789765259e-05
Gd22_18 0 n44 ni18 0 1.93801761121e-05
Gd22_19 0 n44 ni19 0 -2.69957025158e-05
Gd22_20 0 n44 ni20 0 0.000326244483298
Gd22_21 0 n44 ni21 0 0.000558945010528
Gd22_22 0 n44 ni22 0 -0.00158327171391
Gd22_23 0 n44 ni23 0 -0.000325790285352
Gd22_24 0 n44 ni24 0 0.000209111420328
Gd22_25 0 n44 ni25 0 -9.58020907761e-05
Gd22_26 0 n44 ni26 0 7.17996859018e-06
Gd22_27 0 n44 ni27 0 6.49626601179e-05
Gd22_28 0 n44 ni28 0 0.00114747239867
Gd22_29 0 n44 ni29 0 0.00229255632795
Gd22_30 0 n44 ni30 0 -0.000341002411723
Gd22_31 0 n44 ni31 0 0.000245742976004
Gd22_32 0 n44 ni32 0 -3.71823980704e-05
Gc23_129 0 n46 ns129 0 -1.47916828061e-05
Gc23_130 0 n46 ns130 0 3.12076773426e-07
Gc23_131 0 n46 ns131 0 -1.77396695398e-06
Gc23_132 0 n46 ns132 0 -2.72953712497e-06
Gc23_133 0 n46 ns133 0 -5.5532784192e-06
Gc23_134 0 n46 ns134 0 -1.57461685514e-07
Gc23_135 0 n46 ns135 0 -8.5981085107e-07
Gc23_136 0 n46 ns136 0 -1.13303185558e-06
Gc23_137 0 n46 ns137 0 -1.50620155548e-05
Gc23_138 0 n46 ns138 0 3.19179100052e-07
Gc23_139 0 n46 ns139 0 -1.82797677892e-06
Gc23_140 0 n46 ns140 0 -4.00163507526e-06
Gc23_141 0 n46 ns141 0 -5.62410315084e-06
Gc23_142 0 n46 ns142 0 -6.3835544089e-07
Gc23_143 0 n46 ns143 0 -7.89271096538e-07
Gc23_144 0 n46 ns144 0 -1.10776446439e-06
Gc23_145 0 n46 ns145 0 4.41802438122e-06
Gc23_146 0 n46 ns146 0 -4.89953204648e-08
Gc23_147 0 n46 ns147 0 7.48482092281e-07
Gc23_148 0 n46 ns148 0 -4.04150364066e-06
Gc23_149 0 n46 ns149 0 -3.0161971271e-06
Gc23_150 0 n46 ns150 0 5.65313466912e-08
Gc23_151 0 n46 ns151 0 2.48215745122e-08
Gc23_152 0 n46 ns152 0 4.33779109321e-07
Gc23_153 0 n46 ns153 0 5.17091479984e-05
Gc23_154 0 n46 ns154 0 -8.82283467562e-07
Gc23_155 0 n46 ns155 0 6.80720005299e-06
Gc23_156 0 n46 ns156 0 1.78669389651e-06
Gc23_157 0 n46 ns157 0 4.97113112419e-06
Gc23_158 0 n46 ns158 0 5.34172995064e-06
Gc23_159 0 n46 ns159 0 1.77878004493e-06
Gc23_160 0 n46 ns160 0 3.72902072723e-06
Gc23_161 0 n46 ns161 0 -0.000157891414269
Gc23_162 0 n46 ns162 0 3.308961004e-06
Gc23_163 0 n46 ns163 0 -2.1950177423e-05
Gc23_164 0 n46 ns164 0 -4.96536090927e-05
Gc23_165 0 n46 ns165 0 -5.23795027206e-05
Gc23_166 0 n46 ns166 0 -1.81648417013e-05
Gc23_167 0 n46 ns167 0 -6.29681737742e-06
Gc23_168 0 n46 ns168 0 -1.29235588521e-05
Gc23_169 0 n46 ns169 0 0.000702153706474
Gc23_170 0 n46 ns170 0 -1.60958182142e-05
Gc23_171 0 n46 ns171 0 7.61809351702e-05
Gc23_172 0 n46 ns172 0 0.000111084049443
Gc23_173 0 n46 ns173 0 -5.3667063409e-05
Gc23_174 0 n46 ns174 0 -6.50788150424e-05
Gc23_175 0 n46 ns175 0 1.17854112503e-05
Gc23_176 0 n46 ns176 0 4.17672609415e-05
Gc23_177 0 n46 ns177 0 0.00295191386611
Gc23_178 0 n46 ns178 0 -5.20404027502e-05
Gc23_179 0 n46 ns179 0 0.000297818723023
Gc23_180 0 n46 ns180 0 0.000534889018834
Gc23_181 0 n46 ns181 0 0.000228609822567
Gc23_182 0 n46 ns182 0 -0.000102604166166
Gc23_183 0 n46 ns183 0 -1.26998192699e-05
Gc23_184 0 n46 ns184 0 0.000374685832255
Gc23_185 0 n46 ns185 0 6.47767887685e-05
Gc23_186 0 n46 ns186 0 -1.38228417418e-06
Gc23_187 0 n46 ns187 0 -1.65565387546e-05
Gc23_188 0 n46 ns188 0 -2.32145882801e-05
Gc23_189 0 n46 ns189 0 -7.52061869237e-05
Gc23_190 0 n46 ns190 0 -5.65450869799e-05
Gc23_191 0 n46 ns191 0 4.96671616193e-06
Gc23_192 0 n46 ns192 0 -2.09505595987e-05
Gc23_193 0 n46 ns193 0 -0.000188351896852
Gc23_194 0 n46 ns194 0 4.15046223047e-06
Gc23_195 0 n46 ns195 0 -2.6383195687e-05
Gc23_196 0 n46 ns196 0 -5.11428571693e-05
Gc23_197 0 n46 ns197 0 -5.29693161327e-05
Gc23_198 0 n46 ns198 0 -1.17689088319e-05
Gc23_199 0 n46 ns199 0 -7.03144286372e-06
Gc23_200 0 n46 ns200 0 -1.63246759535e-05
Gc23_201 0 n46 ns201 0 -1.61008523467e-05
Gc23_202 0 n46 ns202 0 3.59827497179e-07
Gc23_203 0 n46 ns203 0 -2.06331921685e-06
Gc23_204 0 n46 ns204 0 -5.98599290458e-06
Gc23_205 0 n46 ns205 0 -5.35095720294e-06
Gc23_206 0 n46 ns206 0 -9.22148049252e-07
Gc23_207 0 n46 ns207 0 -6.45801883397e-07
Gc23_208 0 n46 ns208 0 -1.20270738376e-06
Gc23_209 0 n46 ns209 0 3.18023255019e-05
Gc23_210 0 n46 ns210 0 -5.47762019543e-07
Gc23_211 0 n46 ns211 0 4.35062999712e-06
Gc23_212 0 n46 ns212 0 6.2799285415e-07
Gc23_213 0 n46 ns213 0 1.26896283374e-06
Gc23_214 0 n46 ns214 0 3.33791513969e-06
Gc23_215 0 n46 ns215 0 9.20354319055e-07
Gc23_216 0 n46 ns216 0 2.33677321354e-06
Gc23_217 0 n46 ns217 0 -2.36714626784e-05
Gc23_218 0 n46 ns218 0 8.64957387927e-07
Gc23_219 0 n46 ns219 0 -4.00407741026e-06
Gc23_220 0 n46 ns220 0 -8.68811366534e-06
Gc23_221 0 n46 ns221 0 -6.79321679903e-06
Gc23_222 0 n46 ns222 0 6.98559659355e-06
Gc23_223 0 n46 ns223 0 -7.41187393036e-07
Gc23_224 0 n46 ns224 0 -3.2647921404e-06
Gc23_225 0 n46 ns225 0 -0.000678295146722
Gc23_226 0 n46 ns226 0 1.4650463463e-05
Gc23_227 0 n46 ns227 0 -0.000100265801325
Gc23_228 0 n46 ns228 0 -0.000159252700152
Gc23_229 0 n46 ns229 0 -0.000120664269025
Gc23_230 0 n46 ns230 0 -4.52098909272e-05
Gc23_231 0 n46 ns231 0 -1.76077753778e-05
Gc23_232 0 n46 ns232 0 -6.24332445921e-05
Gc23_233 0 n46 ns233 0 0.00129296325347
Gc23_234 0 n46 ns234 0 -1.83063987927e-05
Gc23_235 0 n46 ns235 0 -2.89758585615e-05
Gc23_236 0 n46 ns236 0 0.000370996653913
Gc23_237 0 n46 ns237 0 -6.20836812017e-05
Gc23_238 0 n46 ns238 0 -5.44813082553e-05
Gc23_239 0 n46 ns239 0 4.50852083397e-05
Gc23_240 0 n46 ns240 0 -6.22659363203e-05
Gc23_241 0 n46 ns241 0 0.00150170228499
Gc23_242 0 n46 ns242 0 -2.77113772417e-05
Gc23_243 0 n46 ns243 0 9.39328674134e-05
Gc23_244 0 n46 ns244 0 0.000365584014813
Gc23_245 0 n46 ns245 0 8.94566061998e-06
Gc23_246 0 n46 ns246 0 -3.01103714361e-05
Gc23_247 0 n46 ns247 0 3.70497460607e-05
Gc23_248 0 n46 ns248 0 3.73395384038e-05
Gc23_249 0 n46 ns249 0 -0.000231555473431
Gc23_250 0 n46 ns250 0 4.57349135246e-06
Gc23_251 0 n46 ns251 0 -3.45426840415e-05
Gc23_252 0 n46 ns252 0 -6.68798370633e-05
Gc23_253 0 n46 ns253 0 -8.92243529918e-05
Gc23_254 0 n46 ns254 0 -3.91627588734e-05
Gc23_255 0 n46 ns255 0 -1.04206879445e-05
Gc23_256 0 n46 ns256 0 -2.00611940406e-05
Gd23_17 0 n46 ni17 0 1.34367946382e-05
Gd23_18 0 n46 ni18 0 1.45647470786e-05
Gd23_19 0 n46 ni19 0 -2.22104834109e-06
Gd23_20 0 n46 ni20 0 -4.30734856707e-05
Gd23_21 0 n46 ni21 0 0.000196085987071
Gd23_22 0 n46 ni22 0 -0.000325790285352
Gd23_23 0 n46 ni23 0 -0.00120854489048
Gd23_24 0 n46 ni24 0 0.000399681550558
Gd23_25 0 n46 ni25 0 0.000229292468736
Gd23_26 0 n46 ni26 0 1.78086122525e-05
Gd23_27 0 n46 ni27 0 -2.78568872112e-05
Gd23_28 0 n46 ni28 0 4.32617636639e-05
Gd23_29 0 n46 ni29 0 0.00085421845383
Gd23_30 0 n46 ni30 0 0.00205758093149
Gd23_31 0 n46 ni31 0 0.000310365219524
Gd23_32 0 n46 ni32 0 0.000327283176686
Gc24_129 0 n48 ns129 0 -1.25620906464e-06
Gc24_130 0 n48 ns130 0 4.08974149788e-08
Gc24_131 0 n48 ns131 0 -1.60982709195e-07
Gc24_132 0 n48 ns132 0 -9.16825760851e-07
Gc24_133 0 n48 ns133 0 -8.07864029922e-07
Gc24_134 0 n48 ns134 0 2.9464859174e-07
Gc24_135 0 n48 ns135 0 -6.87981632435e-08
Gc24_136 0 n48 ns136 0 -1.24079376585e-07
Gc24_137 0 n48 ns137 0 -3.30015529186e-06
Gc24_138 0 n48 ns138 0 8.08517218538e-08
Gc24_139 0 n48 ns139 0 -4.1069396312e-07
Gc24_140 0 n48 ns140 0 -1.43027707199e-06
Gc24_141 0 n48 ns141 0 -1.4633355967e-06
Gc24_142 0 n48 ns142 0 7.52478281486e-08
Gc24_143 0 n48 ns143 0 -1.65319921253e-07
Gc24_144 0 n48 ns144 0 -2.61099207903e-07
Gc24_145 0 n48 ns145 0 -1.0728648796e-05
Gc24_146 0 n48 ns146 0 2.36920505096e-07
Gc24_147 0 n48 ns147 0 -1.37831665325e-06
Gc24_148 0 n48 ns148 0 -4.46597855045e-06
Gc24_149 0 n48 ns149 0 -3.54116510808e-06
Gc24_150 0 n48 ns150 0 -8.31523477796e-07
Gc24_151 0 n48 ns151 0 -3.92367661306e-07
Gc24_152 0 n48 ns152 0 -7.81671188253e-07
Gc24_153 0 n48 ns153 0 -5.38563464307e-06
Gc24_154 0 n48 ns154 0 1.7010665414e-07
Gc24_155 0 n48 ns155 0 -7.84867720737e-07
Gc24_156 0 n48 ns156 0 -6.40379803217e-06
Gc24_157 0 n48 ns157 0 -2.54063903107e-06
Gc24_158 0 n48 ns158 0 -4.99140861372e-07
Gc24_159 0 n48 ns159 0 -8.31991487463e-09
Gc24_160 0 n48 ns160 0 -4.06454994006e-07
Gc24_161 0 n48 ns161 0 4.98858490247e-05
Gc24_162 0 n48 ns162 0 -8.41613722655e-07
Gc24_163 0 n48 ns163 0 6.67519611143e-06
Gc24_164 0 n48 ns164 0 2.85917292361e-06
Gc24_165 0 n48 ns165 0 3.77290856164e-06
Gc24_166 0 n48 ns166 0 6.04942341069e-06
Gc24_167 0 n48 ns167 0 1.51283826448e-06
Gc24_168 0 n48 ns168 0 3.54572171625e-06
Gc24_169 0 n48 ns169 0 -0.000169376832916
Gc24_170 0 n48 ns170 0 3.61064851698e-06
Gc24_171 0 n48 ns171 0 -2.36873422387e-05
Gc24_172 0 n48 ns172 0 -5.1580872406e-05
Gc24_173 0 n48 ns173 0 -5.08619738567e-05
Gc24_174 0 n48 ns174 0 -1.71329139902e-05
Gc24_175 0 n48 ns175 0 -6.40293377735e-06
Gc24_176 0 n48 ns176 0 -1.3810386846e-05
Gc24_177 0 n48 ns177 0 6.47767887685e-05
Gc24_178 0 n48 ns178 0 -1.38228417418e-06
Gc24_179 0 n48 ns179 0 -1.65565387546e-05
Gc24_180 0 n48 ns180 0 -2.32145882801e-05
Gc24_181 0 n48 ns181 0 -7.52061869237e-05
Gc24_182 0 n48 ns182 0 -5.65450869799e-05
Gc24_183 0 n48 ns183 0 4.96671616193e-06
Gc24_184 0 n48 ns184 0 -2.09505595987e-05
Gc24_185 0 n48 ns185 0 0.00243943725984
Gc24_186 0 n48 ns186 0 -4.01013981524e-05
Gc24_187 0 n48 ns187 0 0.000232317258542
Gc24_188 0 n48 ns188 0 0.000554515292865
Gc24_189 0 n48 ns189 0 0.000135199668747
Gc24_190 0 n48 ns190 0 -8.55522334048e-05
Gc24_191 0 n48 ns191 0 -5.36364373481e-05
Gc24_192 0 n48 ns192 0 0.000361828969118
Gc24_193 0 n48 ns193 0 0.000298469502188
Gc24_194 0 n48 ns194 0 -7.28202934984e-06
Gc24_195 0 n48 ns195 0 1.89434520639e-05
Gc24_196 0 n48 ns196 0 1.25806559363e-05
Gc24_197 0 n48 ns197 0 -0.000101821579636
Gc24_198 0 n48 ns198 0 -8.17212896933e-05
Gc24_199 0 n48 ns199 0 4.07977822429e-06
Gc24_200 0 n48 ns200 0 5.26618616598e-06
Gc24_201 0 n48 ns201 0 -7.82317063008e-06
Gc24_202 0 n48 ns202 0 1.78570270538e-07
Gc24_203 0 n48 ns203 0 -1.03790972311e-06
Gc24_204 0 n48 ns204 0 -2.92565101132e-06
Gc24_205 0 n48 ns205 0 -2.24466951774e-06
Gc24_206 0 n48 ns206 0 -3.21863551552e-07
Gc24_207 0 n48 ns207 0 -2.71006712544e-07
Gc24_208 0 n48 ns208 0 -6.06972782175e-07
Gc24_209 0 n48 ns209 0 -1.48485290281e-05
Gc24_210 0 n48 ns210 0 3.36813311676e-07
Gc24_211 0 n48 ns211 0 -1.93117961481e-06
Gc24_212 0 n48 ns212 0 -5.88402822729e-06
Gc24_213 0 n48 ns213 0 -4.7749632929e-06
Gc24_214 0 n48 ns214 0 -8.54236571696e-07
Gc24_215 0 n48 ns215 0 -5.4733159164e-07
Gc24_216 0 n48 ns216 0 -1.12748424439e-06
Gc24_217 0 n48 ns217 0 2.77757243943e-06
Gc24_218 0 n48 ns218 0 8.12671061269e-08
Gc24_219 0 n48 ns219 0 1.3163611215e-07
Gc24_220 0 n48 ns220 0 -3.82868455244e-06
Gc24_221 0 n48 ns221 0 -5.77811286216e-07
Gc24_222 0 n48 ns222 0 2.49301273114e-06
Gc24_223 0 n48 ns223 0 2.52599116937e-07
Gc24_224 0 n48 ns224 0 -1.07311707093e-07
Gc24_225 0 n48 ns225 0 -7.29200407164e-05
Gc24_226 0 n48 ns226 0 2.0573619414e-06
Gc24_227 0 n48 ns227 0 -1.12256766218e-05
Gc24_228 0 n48 ns228 0 -1.22416716916e-05
Gc24_229 0 n48 ns229 0 -6.15492280793e-06
Gc24_230 0 n48 ns230 0 1.10599114214e-05
Gc24_231 0 n48 ns231 0 -1.79804228454e-06
Gc24_232 0 n48 ns232 0 -7.81932768613e-06
Gc24_233 0 n48 ns233 0 -0.000416599261666
Gc24_234 0 n48 ns234 0 8.7272101259e-06
Gc24_235 0 n48 ns235 0 -6.29683440543e-05
Gc24_236 0 n48 ns236 0 -0.000107319559922
Gc24_237 0 n48 ns237 0 -0.000104110516999
Gc24_238 0 n48 ns238 0 -4.45713692311e-05
Gc24_239 0 n48 ns239 0 -1.28187691966e-05
Gc24_240 0 n48 ns240 0 -3.91193847136e-05
Gc24_241 0 n48 ns241 0 0.00124437971124
Gc24_242 0 n48 ns242 0 -1.70907301975e-05
Gc24_243 0 n48 ns243 0 -5.76368441398e-05
Gc24_244 0 n48 ns244 0 0.000203442363139
Gc24_245 0 n48 ns245 0 -9.88018390123e-06
Gc24_246 0 n48 ns246 0 -9.11873638941e-05
Gc24_247 0 n48 ns247 0 8.39017295758e-05
Gc24_248 0 n48 ns248 0 -0.000116067609704
Gc24_249 0 n48 ns249 0 0.00148408529907
Gc24_250 0 n48 ns250 0 -2.7796314362e-05
Gc24_251 0 n48 ns251 0 0.000103661824823
Gc24_252 0 n48 ns252 0 0.000396942021576
Gc24_253 0 n48 ns253 0 -1.59415601016e-05
Gc24_254 0 n48 ns254 0 -2.59341134303e-05
Gc24_255 0 n48 ns255 0 2.40672500713e-05
Gc24_256 0 n48 ns256 0 5.52197315714e-05
Gd24_17 0 n48 ni17 0 1.91103853184e-06
Gd24_18 0 n48 ni18 0 3.81327801596e-06
Gd24_19 0 n48 ni19 0 1.21001062324e-05
Gd24_20 0 n48 ni20 0 1.02280488526e-05
Gd24_21 0 n48 ni21 0 -4.3100061764e-05
Gd24_22 0 n48 ni22 0 0.000209111420328
Gd24_23 0 n48 ni23 0 0.000399681550558
Gd24_24 0 n48 ni24 0 -0.000781678154864
Gd24_25 0 n48 ni25 0 0.000132661865229
Gd24_26 0 n48 ni26 0 9.03634275714e-06
Gd24_27 0 n48 ni27 0 1.6976596658e-05
Gd24_28 0 n48 ni28 0 4.56627397379e-06
Gd24_29 0 n48 ni29 0 9.61544824062e-05
Gd24_30 0 n48 ni30 0 0.00056648777286
Gd24_31 0 n48 ni31 0 0.00249515285216
Gd24_32 0 n48 ni32 0 0.000130833325332
Gc25_129 0 n50 ns129 0 1.67725608497e-06
Gc25_130 0 n50 ns130 0 -1.89545011707e-08
Gc25_131 0 n50 ns131 0 2.08393457017e-07
Gc25_132 0 n50 ns132 0 -3.97220728028e-07
Gc25_133 0 n50 ns133 0 2.66068565959e-08
Gc25_134 0 n50 ns134 0 4.58268492725e-07
Gc25_135 0 n50 ns135 0 7.09971356125e-08
Gc25_136 0 n50 ns136 0 9.4965052511e-08
Gc25_137 0 n50 ns137 0 1.141003238e-10
Gc25_138 0 n50 ns138 0 1.31414501056e-08
Gc25_139 0 n50 ns139 0 1.66909831802e-08
Gc25_140 0 n50 ns140 0 -3.93996171683e-07
Gc25_141 0 n50 ns141 0 -5.95047448575e-07
Gc25_142 0 n50 ns142 0 4.29406188071e-07
Gc25_143 0 n50 ns143 0 -4.8404230285e-08
Gc25_144 0 n50 ns144 0 -2.71601396184e-08
Gc25_145 0 n50 ns145 0 -5.16237636419e-06
Gc25_146 0 n50 ns146 0 1.15175557401e-07
Gc25_147 0 n50 ns147 0 -5.79125061106e-07
Gc25_148 0 n50 ns148 0 -1.38421003863e-06
Gc25_149 0 n50 ns149 0 -2.67882728836e-06
Gc25_150 0 n50 ns150 0 1.36255822705e-07
Gc25_151 0 n50 ns151 0 -3.60297080737e-07
Gc25_152 0 n50 ns152 0 -3.95732490212e-07
Gc25_153 0 n50 ns153 0 -1.29585490452e-05
Gc25_154 0 n50 ns154 0 2.78515819321e-07
Gc25_155 0 n50 ns155 0 -1.59040419369e-06
Gc25_156 0 n50 ns156 0 -4.93828053284e-06
Gc25_157 0 n50 ns157 0 -4.97049521728e-06
Gc25_158 0 n50 ns158 0 -9.34367104711e-07
Gc25_159 0 n50 ns159 0 -5.80137857788e-07
Gc25_160 0 n50 ns160 0 -9.40202246415e-07
Gc25_161 0 n50 ns161 0 3.07314839005e-06
Gc25_162 0 n50 ns162 0 -3.63272599161e-08
Gc25_163 0 n50 ns163 0 8.08308920139e-07
Gc25_164 0 n50 ns164 0 -4.29492203614e-06
Gc25_165 0 n50 ns165 0 -6.0311872348e-06
Gc25_166 0 n50 ns166 0 -3.37206458522e-08
Gc25_167 0 n50 ns167 0 -3.27225691668e-07
Gc25_168 0 n50 ns168 0 3.68825479228e-07
Gc25_169 0 n50 ns169 0 9.7323880913e-05
Gc25_170 0 n50 ns170 0 -1.87183261737e-06
Gc25_171 0 n50 ns171 0 1.36542410049e-05
Gc25_172 0 n50 ns172 0 9.18009403794e-06
Gc25_173 0 n50 ns173 0 4.7664335293e-06
Gc25_174 0 n50 ns174 0 7.21042618057e-06
Gc25_175 0 n50 ns175 0 2.47540795848e-06
Gc25_176 0 n50 ns176 0 7.49728276233e-06
Gc25_177 0 n50 ns177 0 -0.000188351896852
Gc25_178 0 n50 ns178 0 4.15046223047e-06
Gc25_179 0 n50 ns179 0 -2.6383195687e-05
Gc25_180 0 n50 ns180 0 -5.11428571693e-05
Gc25_181 0 n50 ns181 0 -5.29693161327e-05
Gc25_182 0 n50 ns182 0 -1.17689088319e-05
Gc25_183 0 n50 ns183 0 -7.03144286372e-06
Gc25_184 0 n50 ns184 0 -1.63246759535e-05
Gc25_185 0 n50 ns185 0 0.000298469502188
Gc25_186 0 n50 ns186 0 -7.28202934984e-06
Gc25_187 0 n50 ns187 0 1.89434520639e-05
Gc25_188 0 n50 ns188 0 1.25806559363e-05
Gc25_189 0 n50 ns189 0 -0.000101821579636
Gc25_190 0 n50 ns190 0 -8.17212896933e-05
Gc25_191 0 n50 ns191 0 4.07977822429e-06
Gc25_192 0 n50 ns192 0 5.26618616598e-06
Gc25_193 0 n50 ns193 0 0.00482412265773
Gc25_194 0 n50 ns194 0 -9.41745793617e-05
Gc25_195 0 n50 ns195 0 0.000564754755818
Gc25_196 0 n50 ns196 0 0.000948226465641
Gc25_197 0 n50 ns197 0 0.000340236023701
Gc25_198 0 n50 ns198 0 -8.0390557213e-05
Gc25_199 0 n50 ns199 0 1.63250577656e-05
Gc25_200 0 n50 ns200 0 0.000542659269161
Gc25_201 0 n50 ns201 0 -2.20551803116e-06
Gc25_202 0 n50 ns202 0 5.96563651273e-08
Gc25_203 0 n50 ns203 0 -2.67664482802e-07
Gc25_204 0 n50 ns204 0 -8.00903765654e-07
Gc25_205 0 n50 ns205 0 -1.17333923648e-06
Gc25_206 0 n50 ns206 0 3.49972228782e-07
Gc25_207 0 n50 ns207 0 -1.4676534513e-07
Gc25_208 0 n50 ns208 0 -1.98158055057e-07
Gc25_209 0 n50 ns209 0 -1.35875538918e-05
Gc25_210 0 n50 ns210 0 2.87159301283e-07
Gc25_211 0 n50 ns211 0 -1.62356783139e-06
Gc25_212 0 n50 ns212 0 -2.75694565033e-06
Gc25_213 0 n50 ns213 0 -5.24091861324e-06
Gc25_214 0 n50 ns214 0 -1.9611521658e-07
Gc25_215 0 n50 ns215 0 -7.87212734778e-07
Gc25_216 0 n50 ns216 0 -1.03697069322e-06
Gc25_217 0 n50 ns217 0 -2.45849597891e-05
Gc25_218 0 n50 ns218 0 5.33485310171e-07
Gc25_219 0 n50 ns219 0 -3.11165758654e-06
Gc25_220 0 n50 ns220 0 -7.00390833216e-06
Gc25_221 0 n50 ns221 0 -7.95306681656e-06
Gc25_222 0 n50 ns222 0 -1.03985360159e-06
Gc25_223 0 n50 ns223 0 -1.09156872047e-06
Gc25_224 0 n50 ns224 0 -1.89379088407e-06
Gc25_225 0 n50 ns225 0 4.65815313607e-06
Gc25_226 0 n50 ns226 0 4.7114778579e-08
Gc25_227 0 n50 ns227 0 5.83822376398e-07
Gc25_228 0 n50 ns228 0 -2.87510704481e-06
Gc25_229 0 n50 ns229 0 -2.57803982741e-06
Gc25_230 0 n50 ns230 0 3.37730434843e-06
Gc25_231 0 n50 ns231 0 1.68503252042e-08
Gc25_232 0 n50 ns232 0 -1.29739392451e-08
Gc25_233 0 n50 ns233 0 1.33902058401e-05
Gc25_234 0 n50 ns234 0 5.01568964822e-08
Gc25_235 0 n50 ns235 0 1.58673190283e-06
Gc25_236 0 n50 ns236 0 -7.33827661407e-06
Gc25_237 0 n50 ns237 0 -7.87647664545e-06
Gc25_238 0 n50 ns238 0 6.46051916995e-06
Gc25_239 0 n50 ns239 0 5.87190208234e-08
Gc25_240 0 n50 ns240 0 -1.98930176874e-08
Gc25_241 0 n50 ns241 0 -0.000457770310533
Gc25_242 0 n50 ns242 0 9.48035414528e-06
Gc25_243 0 n50 ns243 0 -6.82936761093e-05
Gc25_244 0 n50 ns244 0 -0.000123778383046
Gc25_245 0 n50 ns245 0 -0.000122416962197
Gc25_246 0 n50 ns246 0 -5.23943178946e-05
Gc25_247 0 n50 ns247 0 -1.43754952682e-05
Gc25_248 0 n50 ns248 0 -4.28130746993e-05
Gc25_249 0 n50 ns249 0 0.00187371620734
Gc25_250 0 n50 ns250 0 -3.17497051811e-05
Gc25_251 0 n50 ns251 0 3.07717004616e-05
Gc25_252 0 n50 ns252 0 0.000305336987388
Gc25_253 0 n50 ns253 0 7.70972823382e-06
Gc25_254 0 n50 ns254 0 -0.000112436701004
Gc25_255 0 n50 ns255 0 9.60324222662e-05
Gc25_256 0 n50 ns256 0 -6.15655091428e-05
Gd25_17 0 n50 ni17 0 -8.50607552001e-07
Gd25_18 0 n50 ni18 0 3.55350447338e-07
Gd25_19 0 n50 ni19 0 4.73051916026e-06
Gd25_20 0 n50 ni20 0 1.35884040403e-05
Gd25_21 0 n50 ni21 0 -3.12519358751e-06
Gd25_22 0 n50 ni22 0 -9.58020907761e-05
Gd25_23 0 n50 ni23 0 0.000229292468736
Gd25_24 0 n50 ni24 0 0.000132661865229
Gd25_25 0 n50 ni25 0 -0.00328185608091
Gd25_26 0 n50 ni26 0 2.52556454644e-06
Gd25_27 0 n50 ni27 0 1.24461582371e-05
Gd25_28 0 n50 ni28 0 2.53776202141e-05
Gd25_29 0 n50 ni29 0 6.37593505202e-07
Gd25_30 0 n50 ni30 0 2.54085872691e-06
Gd25_31 0 n50 ni31 0 0.000614880238506
Gd25_32 0 n50 ni32 0 0.00184398665632
Gc26_129 0 n52 ns129 0 0.000310054649495
Gc26_130 0 n52 ns130 0 -7.5790263544e-06
Gc26_131 0 n52 ns131 0 1.94747088505e-05
Gc26_132 0 n52 ns132 0 -1.95408506006e-06
Gc26_133 0 n52 ns133 0 -9.17915853797e-05
Gc26_134 0 n52 ns134 0 -8.37137922697e-05
Gc26_135 0 n52 ns135 0 8.83866439149e-06
Gc26_136 0 n52 ns136 0 1.52706257142e-06
Gc26_137 0 n52 ns137 0 0.00178206886175
Gc26_138 0 n52 ns138 0 -3.40637084719e-05
Gc26_139 0 n52 ns139 0 0.000135569811946
Gc26_140 0 n52 ns140 0 0.000416849249638
Gc26_141 0 n52 ns141 0 2.44606450997e-05
Gc26_142 0 n52 ns142 0 -3.22037957035e-05
Gc26_143 0 n52 ns143 0 4.05626890389e-05
Gc26_144 0 n52 ns144 0 6.66321845711e-05
Gc26_145 0 n52 ns145 0 0.00127287147905
Gc26_146 0 n52 ns146 0 -1.70232403006e-05
Gc26_147 0 n52 ns147 0 -6.09795598043e-05
Gc26_148 0 n52 ns148 0 0.000267415140037
Gc26_149 0 n52 ns149 0 -3.50050203318e-05
Gc26_150 0 n52 ns150 0 -8.29567995603e-05
Gc26_151 0 n52 ns151 0 7.31693981773e-05
Gc26_152 0 n52 ns152 0 -0.000109603359805
Gc26_153 0 n52 ns153 0 -0.000508213037802
Gc26_154 0 n52 ns154 0 1.08195802248e-05
Gc26_155 0 n52 ns155 0 -7.58612447122e-05
Gc26_156 0 n52 ns156 0 -0.000126150320067
Gc26_157 0 n52 ns157 0 -0.00010990400649
Gc26_158 0 n52 ns158 0 -4.52722846055e-05
Gc26_159 0 n52 ns159 0 -1.48603195403e-05
Gc26_160 0 n52 ns160 0 -4.63364501973e-05
Gc26_161 0 n52 ns161 0 -6.17816254036e-05
Gc26_162 0 n52 ns162 0 1.74986330091e-06
Gc26_163 0 n52 ns163 0 -9.40333936283e-06
Gc26_164 0 n52 ns164 0 -1.34449001868e-05
Gc26_165 0 n52 ns165 0 -8.54082041553e-06
Gc26_166 0 n52 ns166 0 8.35419128121e-06
Gc26_167 0 n52 ns167 0 -1.70450106561e-06
Gc26_168 0 n52 ns168 0 -6.49632100499e-06
Gc26_169 0 n52 ns169 0 -2.44664340862e-07
Gc26_170 0 n52 ns170 0 1.53022803091e-07
Gc26_171 0 n52 ns171 0 -2.87421576414e-07
Gc26_172 0 n52 ns172 0 -3.07995996449e-06
Gc26_173 0 n52 ns173 0 -8.6899931677e-07
Gc26_174 0 n52 ns174 0 3.0667550508e-06
Gc26_175 0 n52 ns175 0 7.73937785179e-08
Gc26_176 0 n52 ns176 0 -4.05074848322e-07
Gc26_177 0 n52 ns177 0 -1.61008523467e-05
Gc26_178 0 n52 ns178 0 3.59827497179e-07
Gc26_179 0 n52 ns179 0 -2.06331921685e-06
Gc26_180 0 n52 ns180 0 -5.98599290458e-06
Gc26_181 0 n52 ns181 0 -5.35095720294e-06
Gc26_182 0 n52 ns182 0 -9.22148049252e-07
Gc26_183 0 n52 ns183 0 -6.45801883397e-07
Gc26_184 0 n52 ns184 0 -1.20270738376e-06
Gc26_185 0 n52 ns185 0 -7.82317063008e-06
Gc26_186 0 n52 ns186 0 1.78570270538e-07
Gc26_187 0 n52 ns187 0 -1.03790972311e-06
Gc26_188 0 n52 ns188 0 -2.92565101132e-06
Gc26_189 0 n52 ns189 0 -2.24466951774e-06
Gc26_190 0 n52 ns190 0 -3.21863551552e-07
Gc26_191 0 n52 ns191 0 -2.71006712544e-07
Gc26_192 0 n52 ns192 0 -6.06972782175e-07
Gc26_193 0 n52 ns193 0 -2.20551803116e-06
Gc26_194 0 n52 ns194 0 5.96563651273e-08
Gc26_195 0 n52 ns195 0 -2.67664482802e-07
Gc26_196 0 n52 ns196 0 -8.00903765654e-07
Gc26_197 0 n52 ns197 0 -1.17333923648e-06
Gc26_198 0 n52 ns198 0 3.49972228782e-07
Gc26_199 0 n52 ns199 0 -1.4676534513e-07
Gc26_200 0 n52 ns200 0 -1.98158055057e-07
Gc26_201 0 n52 ns201 0 0.00251193448623
Gc26_202 0 n52 ns202 0 -4.2713771945e-05
Gc26_203 0 n52 ns203 0 0.000257934816309
Gc26_204 0 n52 ns204 0 0.000558729664045
Gc26_205 0 n52 ns205 0 0.000154868370246
Gc26_206 0 n52 ns206 0 -7.58528130613e-05
Gc26_207 0 n52 ns207 0 -4.94905480023e-05
Gc26_208 0 n52 ns208 0 0.000373116379158
Gc26_209 0 n52 ns209 0 5.56821911567e-05
Gc26_210 0 n52 ns210 0 -1.26594036241e-06
Gc26_211 0 n52 ns211 0 -1.68089689763e-05
Gc26_212 0 n52 ns212 0 -1.58843340394e-05
Gc26_213 0 n52 ns213 0 -8.83578894e-05
Gc26_214 0 n52 ns214 0 -6.04027503407e-05
Gc26_215 0 n52 ns215 0 8.95068250094e-07
Gc26_216 0 n52 ns216 0 -1.74118722635e-05
Gc26_217 0 n52 ns217 0 -0.00018827456904
Gc26_218 0 n52 ns218 0 4.13143306466e-06
Gc26_219 0 n52 ns219 0 -2.66019243087e-05
Gc26_220 0 n52 ns220 0 -5.18009944935e-05
Gc26_221 0 n52 ns221 0 -4.77679411483e-05
Gc26_222 0 n52 ns222 0 -1.3384243664e-05
Gc26_223 0 n52 ns223 0 -6.62046115786e-06
Gc26_224 0 n52 ns224 0 -1.56929449014e-05
Gc26_225 0 n52 ns225 0 6.1787282259e-05
Gc26_226 0 n52 ns226 0 -1.09162369067e-06
Gc26_227 0 n52 ns227 0 8.348810839e-06
Gc26_228 0 n52 ns228 0 4.51813876628e-06
Gc26_229 0 n52 ns229 0 5.13013748845e-06
Gc26_230 0 n52 ns230 0 6.42711146867e-06
Gc26_231 0 n52 ns231 0 1.84263697676e-06
Gc26_232 0 n52 ns232 0 4.57907597193e-06
Gc26_233 0 n52 ns233 0 -7.14200261755e-06
Gc26_234 0 n52 ns234 0 2.01916189915e-07
Gc26_235 0 n52 ns235 0 -9.28668116194e-07
Gc26_236 0 n52 ns236 0 -5.57265812495e-06
Gc26_237 0 n52 ns237 0 -3.77867555255e-06
Gc26_238 0 n52 ns238 0 -1.88548786289e-07
Gc26_239 0 n52 ns239 0 -2.62446667277e-07
Gc26_240 0 n52 ns240 0 -5.46261921005e-07
Gc26_241 0 n52 ns241 0 -1.12064892543e-05
Gc26_242 0 n52 ns242 0 2.47598106005e-07
Gc26_243 0 n52 ns243 0 -1.44796052741e-06
Gc26_244 0 n52 ns244 0 -4.51788056499e-06
Gc26_245 0 n52 ns245 0 -3.56374876056e-06
Gc26_246 0 n52 ns246 0 -8.33524767247e-07
Gc26_247 0 n52 ns247 0 -4.0589357044e-07
Gc26_248 0 n52 ns248 0 -8.19269843515e-07
Gc26_249 0 n52 ns249 0 -4.08222680894e-06
Gc26_250 0 n52 ns250 0 9.63011977173e-08
Gc26_251 0 n52 ns251 0 -5.00258096905e-07
Gc26_252 0 n52 ns252 0 -1.34727374393e-06
Gc26_253 0 n52 ns253 0 -1.7440016758e-06
Gc26_254 0 n52 ns254 0 1.11787171816e-07
Gc26_255 0 n52 ns255 0 -2.26493397531e-07
Gc26_256 0 n52 ns256 0 -3.21301083324e-07
Gd26_17 0 n52 ni17 0 0.000139649861222
Gd26_18 0 n52 ni18 0 -2.12815643513e-05
Gd26_19 0 n52 ni19 0 0.00257494590141
Gd26_20 0 n52 ni20 0 0.000665020699165
Gd26_21 0 n52 ni21 0 8.31518675384e-05
Gd26_22 0 n52 ni22 0 7.17996859018e-06
Gd26_23 0 n52 ni23 0 1.78086122525e-05
Gd26_24 0 n52 ni24 0 9.03634275714e-06
Gd26_25 0 n52 ni25 0 2.52556454644e-06
Gd26_26 0 n52 ni26 0 -0.00111370708785
Gd26_27 0 n52 ni27 0 0.000395681513498
Gd26_28 0 n52 ni28 0 0.000229938919943
Gd26_29 0 n52 ni29 0 -5.57271017975e-05
Gd26_30 0 n52 ni30 0 1.05510764412e-05
Gd26_31 0 n52 ni31 0 1.26247628802e-05
Gd26_32 0 n52 ni32 0 4.33959101293e-06
Gc27_129 0 n54 ns129 0 -0.000182158362103
Gc27_130 0 n54 ns130 0 4.02845363093e-06
Gc27_131 0 n54 ns131 0 -2.55371836663e-05
Gc27_132 0 n54 ns132 0 -4.97734747553e-05
Gc27_133 0 n54 ns133 0 -5.17000566399e-05
Gc27_134 0 n54 ns134 0 -1.10632181189e-05
Gc27_135 0 n54 ns135 0 -6.80721247628e-06
Gc27_136 0 n54 ns136 0 -1.58904781004e-05
Gc27_137 0 n54 ns137 0 -0.000267174996208
Gc27_138 0 n54 ns138 0 5.3447858213e-06
Gc27_139 0 n54 ns139 0 -3.94151121682e-05
Gc27_140 0 n54 ns140 0 -7.5982279035e-05
Gc27_141 0 n54 ns141 0 -9.31847931764e-05
Gc27_142 0 n54 ns142 0 -4.10644691591e-05
Gc27_143 0 n54 ns143 0 -1.12262584765e-05
Gc27_144 0 n54 ns144 0 -2.27800045622e-05
Gc27_145 0 n54 ns145 0 0.00166906749824
Gc27_146 0 n54 ns146 0 -3.15684708875e-05
Gc27_147 0 n54 ns147 0 0.000122405720945
Gc27_148 0 n54 ns148 0 0.000417289081472
Gc27_149 0 n54 ns149 0 1.90010912889e-05
Gc27_150 0 n54 ns150 0 -2.18361121753e-05
Gc27_151 0 n54 ns151 0 3.58491100484e-05
Gc27_152 0 n54 ns152 0 5.92064875233e-05
Gc27_153 0 n54 ns153 0 0.00130887914861
Gc27_154 0 n54 ns154 0 -1.8676172166e-05
Gc27_155 0 n54 ns155 0 -3.47104426868e-05
Gc27_156 0 n54 ns156 0 0.000290435613173
Gc27_157 0 n54 ns157 0 -2.68253148113e-05
Gc27_158 0 n54 ns158 0 -7.24735164399e-05
Gc27_159 0 n54 ns159 0 6.49422394252e-05
Gc27_160 0 n54 ns160 0 -8.1551587668e-05
Gc27_161 0 n54 ns161 0 -0.000531780502685
Gc27_162 0 n54 ns162 0 1.13471956681e-05
Gc27_163 0 n54 ns163 0 -7.97480222113e-05
Gc27_164 0 n54 ns164 0 -0.000129903300348
Gc27_165 0 n54 ns165 0 -0.000109889199387
Gc27_166 0 n54 ns166 0 -4.42226622106e-05
Gc27_167 0 n54 ns167 0 -1.4473930927e-05
Gc27_168 0 n54 ns168 0 -5.0179212223e-05
Gc27_169 0 n54 ns169 0 -4.4516484898e-05
Gc27_170 0 n54 ns170 0 1.37551926006e-06
Gc27_171 0 n54 ns171 0 -7.07019150765e-06
Gc27_172 0 n54 ns172 0 -8.3552148196e-06
Gc27_173 0 n54 ns173 0 -6.42900882486e-06
Gc27_174 0 n54 ns174 0 9.65652119656e-06
Gc27_175 0 n54 ns175 0 -1.27291011538e-06
Gc27_176 0 n54 ns176 0 -5.36127815906e-06
Gc27_177 0 n54 ns177 0 3.18023255019e-05
Gc27_178 0 n54 ns178 0 -5.47762019543e-07
Gc27_179 0 n54 ns179 0 4.35062999712e-06
Gc27_180 0 n54 ns180 0 6.2799285415e-07
Gc27_181 0 n54 ns181 0 1.26896283374e-06
Gc27_182 0 n54 ns182 0 3.33791513969e-06
Gc27_183 0 n54 ns183 0 9.20354319055e-07
Gc27_184 0 n54 ns184 0 2.33677321354e-06
Gc27_185 0 n54 ns185 0 -1.48485290281e-05
Gc27_186 0 n54 ns186 0 3.36813311676e-07
Gc27_187 0 n54 ns187 0 -1.93117961481e-06
Gc27_188 0 n54 ns188 0 -5.88402822729e-06
Gc27_189 0 n54 ns189 0 -4.7749632929e-06
Gc27_190 0 n54 ns190 0 -8.54236571696e-07
Gc27_191 0 n54 ns191 0 -5.4733159164e-07
Gc27_192 0 n54 ns192 0 -1.12748424439e-06
Gc27_193 0 n54 ns193 0 -1.35875538918e-05
Gc27_194 0 n54 ns194 0 2.87159301283e-07
Gc27_195 0 n54 ns195 0 -1.62356783139e-06
Gc27_196 0 n54 ns196 0 -2.75694565033e-06
Gc27_197 0 n54 ns197 0 -5.24091861324e-06
Gc27_198 0 n54 ns198 0 -1.9611521658e-07
Gc27_199 0 n54 ns199 0 -7.87212734778e-07
Gc27_200 0 n54 ns200 0 -1.03697069322e-06
Gc27_201 0 n54 ns201 0 5.56821911567e-05
Gc27_202 0 n54 ns202 0 -1.26594036241e-06
Gc27_203 0 n54 ns203 0 -1.68089689763e-05
Gc27_204 0 n54 ns204 0 -1.58843340394e-05
Gc27_205 0 n54 ns205 0 -8.83578894e-05
Gc27_206 0 n54 ns206 0 -6.04027503407e-05
Gc27_207 0 n54 ns207 0 8.95068250094e-07
Gc27_208 0 n54 ns208 0 -1.74118722635e-05
Gc27_209 0 n54 ns209 0 0.00248805566046
Gc27_210 0 n54 ns210 0 -4.1181195092e-05
Gc27_211 0 n54 ns211 0 0.000230244143848
Gc27_212 0 n54 ns212 0 0.00050469732451
Gc27_213 0 n54 ns213 0 0.000161685381596
Gc27_214 0 n54 ns214 0 -9.87546384096e-05
Gc27_215 0 n54 ns215 0 -3.65068970531e-05
Gc27_216 0 n54 ns216 0 0.00034518809125
Gc27_217 0 n54 ns217 0 0.000504424704303
Gc27_218 0 n54 ns218 0 -1.14984754973e-05
Gc27_219 0 n54 ns219 0 4.76295253701e-05
Gc27_220 0 n54 ns220 0 6.5701674109e-05
Gc27_221 0 n54 ns221 0 -5.42387942364e-05
Gc27_222 0 n54 ns222 0 -6.07300266646e-05
Gc27_223 0 n54 ns223 0 1.08664459975e-05
Gc27_224 0 n54 ns224 0 2.18283228276e-05
Gc27_225 0 n54 ns225 0 -0.000163302929946
Gc27_226 0 n54 ns226 0 3.39678208492e-06
Gc27_227 0 n54 ns227 0 -2.26179114945e-05
Gc27_228 0 n54 ns228 0 -5.31492742708e-05
Gc27_229 0 n54 ns229 0 -5.39115647609e-05
Gc27_230 0 n54 ns230 0 -2.01533228426e-05
Gc27_231 0 n54 ns231 0 -6.4025326624e-06
Gc27_232 0 n54 ns232 0 -1.30906550953e-05
Gc27_233 0 n54 ns233 0 4.1355917412e-05
Gc27_234 0 n54 ns234 0 -6.72047735793e-07
Gc27_235 0 n54 ns235 0 5.43291143996e-06
Gc27_236 0 n54 ns236 0 8.68569192634e-07
Gc27_237 0 n54 ns237 0 2.8317596651e-06
Gc27_238 0 n54 ns238 0 5.07424372759e-06
Gc27_239 0 n54 ns239 0 1.34210249701e-06
Gc27_240 0 n54 ns240 0 2.85041012946e-06
Gc27_241 0 n54 ns241 0 1.26588162345e-06
Gc27_242 0 n54 ns242 0 1.97037590375e-08
Gc27_243 0 n54 ns243 0 2.66911264936e-07
Gc27_244 0 n54 ns244 0 -4.72465584684e-06
Gc27_245 0 n54 ns245 0 -3.00456203151e-06
Gc27_246 0 n54 ns246 0 -1.32292346428e-07
Gc27_247 0 n54 ns247 0 -6.04545900448e-09
Gc27_248 0 n54 ns248 0 1.64820160386e-07
Gc27_249 0 n54 ns249 0 -1.41157795285e-05
Gc27_250 0 n54 ns250 0 3.00381887275e-07
Gc27_251 0 n54 ns251 0 -1.71623590345e-06
Gc27_252 0 n54 ns252 0 -3.95139921113e-06
Gc27_253 0 n54 ns253 0 -5.3040850564e-06
Gc27_254 0 n54 ns254 0 -6.30088140268e-07
Gc27_255 0 n54 ns255 0 -7.28929730822e-07
Gc27_256 0 n54 ns256 0 -1.03753106782e-06
Gd27_17 0 n54 ni17 0 0.000222617609962
Gd27_18 0 n54 ni18 0 0.000364881563081
Gd27_19 0 n54 ni19 0 4.47447586163e-05
Gd27_20 0 n54 ni20 0 0.00218462950339
Gd27_21 0 n54 ni21 0 0.000697977125634
Gd27_22 0 n54 ni22 0 6.49626601179e-05
Gd27_23 0 n54 ni23 0 -2.78568872112e-05
Gd27_24 0 n54 ni24 0 1.6976596658e-05
Gd27_25 0 n54 ni25 0 1.24461582371e-05
Gd27_26 0 n54 ni26 0 0.000395681513498
Gd27_27 0 n54 ni27 0 -0.000679194867621
Gd27_28 0 n54 ni28 0 -0.000105819315704
Gd27_29 0 n54 ni29 0 0.000201935722417
Gd27_30 0 n54 ni30 0 -3.31026307353e-05
Gd27_31 0 n54 ni31 0 1.6371865763e-06
Gd27_32 0 n54 ni32 0 1.38176184722e-05
Gc28_129 0 n56 ns129 0 7.733002638e-05
Gc28_130 0 n56 ns130 0 -1.42954198782e-06
Gc28_131 0 n56 ns131 0 1.07058650543e-05
Gc28_132 0 n56 ns132 0 6.19313766866e-06
Gc28_133 0 n56 ns133 0 4.05951133347e-06
Gc28_134 0 n56 ns134 0 6.9131254031e-06
Gc28_135 0 n56 ns135 0 2.07944567914e-06
Gc28_136 0 n56 ns136 0 5.76371935762e-06
Gc28_137 0 n56 ns137 0 3.32870787667e-05
Gc28_138 0 n56 ns138 0 -5.00182165155e-07
Gc28_139 0 n56 ns139 0 4.54448540439e-06
Gc28_140 0 n56 ns140 0 -6.23033590648e-06
Gc28_141 0 n56 ns141 0 -5.70600452125e-06
Gc28_142 0 n56 ns142 0 2.33656965896e-06
Gc28_143 0 n56 ns143 0 6.18588789146e-07
Gc28_144 0 n56 ns144 0 2.48166174707e-06
Gc28_145 0 n56 ns145 0 -0.00017177073103
Gc28_146 0 n56 ns146 0 3.03997583428e-06
Gc28_147 0 n56 ns147 0 -2.5688780132e-05
Gc28_148 0 n56 ns148 0 -6.60011769802e-05
Gc28_149 0 n56 ns149 0 -8.99652185167e-05
Gc28_150 0 n56 ns150 0 -4.82944389287e-05
Gc28_151 0 n56 ns151 0 -9.03026798271e-06
Gc28_152 0 n56 ns152 0 -1.37709351205e-05
Gc28_153 0 n56 ns153 0 0.00156320061994
Gc28_154 0 n56 ns154 0 -2.93045088013e-05
Gc28_155 0 n56 ns155 0 0.000109309459108
Gc28_156 0 n56 ns156 0 0.000391708020177
Gc28_157 0 n56 ns157 0 8.39797280059e-06
Gc28_158 0 n56 ns158 0 -2.70096610872e-05
Gc28_159 0 n56 ns159 0 3.25200382389e-05
Gc28_160 0 n56 ns160 0 5.36158478825e-05
Gc28_161 0 n56 ns161 0 0.00199390528219
Gc28_162 0 n56 ns162 0 -3.21546787817e-05
Gc28_163 0 n56 ns163 0 3.61632466142e-06
Gc28_164 0 n56 ns164 0 0.000264246952066
Gc28_165 0 n56 ns165 0 6.72188830779e-05
Gc28_166 0 n56 ns166 0 -0.000119199496022
Gc28_167 0 n56 ns167 0 0.000126839976001
Gc28_168 0 n56 ns168 0 -0.000104421539545
Gc28_169 0 n56 ns169 0 -0.00094957645976
Gc28_170 0 n56 ns170 0 2.08885327754e-05
Gc28_171 0 n56 ns171 0 -0.000138802811919
Gc28_172 0 n56 ns172 0 -0.000214130955143
Gc28_173 0 n56 ns173 0 -0.000130656649253
Gc28_174 0 n56 ns174 0 -4.17738721932e-05
Gc28_175 0 n56 ns175 0 -2.16205792165e-05
Gc28_176 0 n56 ns176 0 -8.70011645526e-05
Gc28_177 0 n56 ns177 0 -2.36714626784e-05
Gc28_178 0 n56 ns178 0 8.64957387927e-07
Gc28_179 0 n56 ns179 0 -4.00407741026e-06
Gc28_180 0 n56 ns180 0 -8.68811366533e-06
Gc28_181 0 n56 ns181 0 -6.79321679903e-06
Gc28_182 0 n56 ns182 0 6.98559659355e-06
Gc28_183 0 n56 ns183 0 -7.41187393036e-07
Gc28_184 0 n56 ns184 0 -3.2647921404e-06
Gc28_185 0 n56 ns185 0 2.77757243943e-06
Gc28_186 0 n56 ns186 0 8.12671061269e-08
Gc28_187 0 n56 ns187 0 1.3163611215e-07
Gc28_188 0 n56 ns188 0 -3.82868455244e-06
Gc28_189 0 n56 ns189 0 -5.77811286216e-07
Gc28_190 0 n56 ns190 0 2.49301273114e-06
Gc28_191 0 n56 ns191 0 2.52599116937e-07
Gc28_192 0 n56 ns192 0 -1.07311707093e-07
Gc28_193 0 n56 ns193 0 -2.45849597891e-05
Gc28_194 0 n56 ns194 0 5.33485310171e-07
Gc28_195 0 n56 ns195 0 -3.11165758654e-06
Gc28_196 0 n56 ns196 0 -7.00390833216e-06
Gc28_197 0 n56 ns197 0 -7.95306681656e-06
Gc28_198 0 n56 ns198 0 -1.03985360159e-06
Gc28_199 0 n56 ns199 0 -1.09156872047e-06
Gc28_200 0 n56 ns200 0 -1.89379088407e-06
Gc28_201 0 n56 ns201 0 -0.00018827456904
Gc28_202 0 n56 ns202 0 4.13143306466e-06
Gc28_203 0 n56 ns203 0 -2.66019243087e-05
Gc28_204 0 n56 ns204 0 -5.18009944935e-05
Gc28_205 0 n56 ns205 0 -4.77679411483e-05
Gc28_206 0 n56 ns206 0 -1.3384243664e-05
Gc28_207 0 n56 ns207 0 -6.62046115786e-06
Gc28_208 0 n56 ns208 0 -1.56929449014e-05
Gc28_209 0 n56 ns209 0 0.000504424704303
Gc28_210 0 n56 ns210 0 -1.14984754973e-05
Gc28_211 0 n56 ns211 0 4.76295253701e-05
Gc28_212 0 n56 ns212 0 6.5701674109e-05
Gc28_213 0 n56 ns213 0 -5.42387942364e-05
Gc28_214 0 n56 ns214 0 -6.07300266646e-05
Gc28_215 0 n56 ns215 0 1.08664459975e-05
Gc28_216 0 n56 ns216 0 2.18283228276e-05
Gc28_217 0 n56 ns217 0 0.00204196224529
Gc28_218 0 n56 ns218 0 -3.30176948129e-05
Gc28_219 0 n56 ns219 0 0.000225458410692
Gc28_220 0 n56 ns220 0 0.000588901108749
Gc28_221 0 n56 ns221 0 7.96862212591e-05
Gc28_222 0 n56 ns222 0 -4.9191433724e-05
Gc28_223 0 n56 ns223 0 -9.60232991003e-05
Gc28_224 0 n56 ns224 0 0.00039066116816
Gc28_225 0 n56 ns225 0 0.000285895561059
Gc28_226 0 n56 ns226 0 -6.69512671712e-06
Gc28_227 0 n56 ns227 0 1.56806688204e-05
Gc28_228 0 n56 ns228 0 5.10737983647e-06
Gc28_229 0 n56 ns229 0 -6.94760053029e-05
Gc28_230 0 n56 ns230 0 -7.00510814387e-05
Gc28_231 0 n56 ns231 0 9.3122775697e-06
Gc28_232 0 n56 ns232 0 1.06394160587e-07
Gc28_233 0 n56 ns233 0 -0.000220325407771
Gc28_234 0 n56 ns234 0 5.04732577646e-06
Gc28_235 0 n56 ns235 0 -3.18589915483e-05
Gc28_236 0 n56 ns236 0 -4.7531801923e-05
Gc28_237 0 n56 ns237 0 -4.08581896209e-05
Gc28_238 0 n56 ns238 0 -4.00906268301e-06
Gc28_239 0 n56 ns239 0 -6.82328725228e-06
Gc28_240 0 n56 ns240 0 -1.99142879207e-05
Gc28_241 0 n56 ns241 0 4.11707815558e-05
Gc28_242 0 n56 ns242 0 -6.34907008116e-07
Gc28_243 0 n56 ns243 0 5.2283705931e-06
Gc28_244 0 n56 ns244 0 2.25341054598e-06
Gc28_245 0 n56 ns245 0 4.85328957022e-06
Gc28_246 0 n56 ns246 0 6.32853351275e-06
Gc28_247 0 n56 ns247 0 1.44768687659e-06
Gc28_248 0 n56 ns248 0 2.70655127281e-06
Gc28_249 0 n56 ns249 0 -1.04323121728e-05
Gc28_250 0 n56 ns250 0 2.65625266703e-07
Gc28_251 0 n56 ns251 0 -1.2887555747e-06
Gc28_252 0 n56 ns252 0 -5.49192986133e-06
Gc28_253 0 n56 ns253 0 -5.18261684693e-06
Gc28_254 0 n56 ns254 0 -1.16653793939e-07
Gc28_255 0 n56 ns255 0 -5.19051296579e-07
Gc28_256 0 n56 ns256 0 -8.02298559639e-07
Gd28_17 0 n56 ni17 0 -7.31066984986e-05
Gd28_18 0 n56 ni18 0 -2.12523804366e-05
Gd28_19 0 n56 ni19 0 0.000262585654946
Gd28_20 0 n56 ni20 0 0.000133009848401
Gd28_21 0 n56 ni21 0 0.00242730950401
Gd28_22 0 n56 ni22 0 0.00114747239867
Gd28_23 0 n56 ni23 0 4.32617636639e-05
Gd28_24 0 n56 ni24 0 4.56627397379e-06
Gd28_25 0 n56 ni25 0 2.53776202141e-05
Gd28_26 0 n56 ni26 0 0.000229938919943
Gd28_27 0 n56 ni27 0 -0.000105819315704
Gd28_28 0 n56 ni28 0 -0.00117887152163
Gd28_29 0 n56 ni29 0 0.00015478569166
Gd28_30 0 n56 ni30 0 0.000267411405598
Gd28_31 0 n56 ni31 0 -3.16853273065e-05
Gd28_32 0 n56 ni32 0 1.27444282105e-05
Gc29_129 0 n58 ns129 0 4.9081659875e-06
Gc29_130 0 n58 ns130 0 -7.3050743847e-08
Gc29_131 0 n58 ns131 0 1.0356195598e-06
Gc29_132 0 n58 ns132 0 -4.51008781946e-06
Gc29_133 0 n58 ns133 0 -5.52285259528e-06
Gc29_134 0 n58 ns134 0 -1.29066089474e-07
Gc29_135 0 n58 ns135 0 -2.06717282931e-07
Gc29_136 0 n58 ns136 0 5.30744237983e-07
Gc29_137 0 n58 ns137 0 3.79524285912e-05
Gc29_138 0 n58 ns138 0 -7.1416073835e-07
Gc29_139 0 n58 ns139 0 5.43240328863e-06
Gc29_140 0 n58 ns140 0 1.10493777751e-06
Gc29_141 0 n58 ns141 0 -1.3867833371e-08
Gc29_142 0 n58 ns142 0 2.55301134937e-06
Gc29_143 0 n58 ns143 0 8.72325500788e-07
Gc29_144 0 n58 ns144 0 3.07434730433e-06
Gc29_145 0 n58 ns145 0 3.84017844558e-05
Gc29_146 0 n58 ns146 0 -6.21160805768e-07
Gc29_147 0 n58 ns147 0 5.29937603072e-06
Gc29_148 0 n58 ns148 0 -7.1009321353e-06
Gc29_149 0 n58 ns149 0 -5.09336172222e-06
Gc29_150 0 n58 ns150 0 1.553232906e-06
Gc29_151 0 n58 ns151 0 8.77393960938e-07
Gc29_152 0 n58 ns152 0 3.03333521248e-06
Gc29_153 0 n58 ns153 0 -0.000170186034785
Gc29_154 0 n58 ns154 0 3.03358613983e-06
Gc29_155 0 n58 ns155 0 -2.58088438595e-05
Gc29_156 0 n58 ns156 0 -6.8780230585e-05
Gc29_157 0 n58 ns157 0 -8.72485474163e-05
Gc29_158 0 n58 ns158 0 -4.85698399507e-05
Gc29_159 0 n58 ns159 0 -8.30723890537e-06
Gc29_160 0 n58 ns160 0 -1.40684582433e-05
Gc29_161 0 n58 ns161 0 0.00285122941534
Gc29_162 0 n58 ns162 0 -5.76952618647e-05
Gc29_163 0 n58 ns163 0 0.000287364733151
Gc29_164 0 n58 ns164 0 0.000666227611578
Gc29_165 0 n58 ns165 0 0.000107110229529
Gc29_166 0 n58 ns166 0 -1.04027360321e-05
Gc29_167 0 n58 ns167 0 5.52341999835e-05
Gc29_168 0 n58 ns168 0 0.000167912032143
Gc29_169 0 n58 ns169 0 0.00253107630446
Gc29_170 0 n58 ns170 0 -4.3690007843e-05
Gc29_171 0 n58 ns171 0 5.36737371871e-05
Gc29_172 0 n58 ns172 0 0.000227173564971
Gc29_173 0 n58 ns173 0 0.000157374025965
Gc29_174 0 n58 ns174 0 -0.000152362149267
Gc29_175 0 n58 ns175 0 0.000173429951137
Gc29_176 0 n58 ns176 0 -0.000104104854591
Gc29_177 0 n58 ns177 0 -0.000678295146722
Gc29_178 0 n58 ns178 0 1.4650463463e-05
Gc29_179 0 n58 ns179 0 -0.000100265801325
Gc29_180 0 n58 ns180 0 -0.000159252700152
Gc29_181 0 n58 ns181 0 -0.000120664269025
Gc29_182 0 n58 ns182 0 -4.52098909272e-05
Gc29_183 0 n58 ns183 0 -1.76077753778e-05
Gc29_184 0 n58 ns184 0 -6.24332445921e-05
Gc29_185 0 n58 ns185 0 -7.29200407164e-05
Gc29_186 0 n58 ns186 0 2.0573619414e-06
Gc29_187 0 n58 ns187 0 -1.12256766218e-05
Gc29_188 0 n58 ns188 0 -1.22416716916e-05
Gc29_189 0 n58 ns189 0 -6.15492280793e-06
Gc29_190 0 n58 ns190 0 1.10599114214e-05
Gc29_191 0 n58 ns191 0 -1.79804228454e-06
Gc29_192 0 n58 ns192 0 -7.81932768613e-06
Gc29_193 0 n58 ns193 0 4.65815313607e-06
Gc29_194 0 n58 ns194 0 4.7114778579e-08
Gc29_195 0 n58 ns195 0 5.83822376398e-07
Gc29_196 0 n58 ns196 0 -2.87510704481e-06
Gc29_197 0 n58 ns197 0 -2.57803982741e-06
Gc29_198 0 n58 ns198 0 3.37730434843e-06
Gc29_199 0 n58 ns199 0 1.68503252042e-08
Gc29_200 0 n58 ns200 0 -1.29739392451e-08
Gc29_201 0 n58 ns201 0 6.1787282259e-05
Gc29_202 0 n58 ns202 0 -1.09162369067e-06
Gc29_203 0 n58 ns203 0 8.348810839e-06
Gc29_204 0 n58 ns204 0 4.51813876628e-06
Gc29_205 0 n58 ns205 0 5.13013748845e-06
Gc29_206 0 n58 ns206 0 6.42711146867e-06
Gc29_207 0 n58 ns207 0 1.84263697676e-06
Gc29_208 0 n58 ns208 0 4.57907597193e-06
Gc29_209 0 n58 ns209 0 -0.000163302929946
Gc29_210 0 n58 ns210 0 3.39678208492e-06
Gc29_211 0 n58 ns211 0 -2.26179114945e-05
Gc29_212 0 n58 ns212 0 -5.31492742708e-05
Gc29_213 0 n58 ns213 0 -5.39115647609e-05
Gc29_214 0 n58 ns214 0 -2.01533228426e-05
Gc29_215 0 n58 ns215 0 -6.4025326624e-06
Gc29_216 0 n58 ns216 0 -1.30906550953e-05
Gc29_217 0 n58 ns217 0 0.000285895561059
Gc29_218 0 n58 ns218 0 -6.69512671712e-06
Gc29_219 0 n58 ns219 0 1.56806688204e-05
Gc29_220 0 n58 ns220 0 5.10737983647e-06
Gc29_221 0 n58 ns221 0 -6.94760053029e-05
Gc29_222 0 n58 ns222 0 -7.00510814387e-05
Gc29_223 0 n58 ns223 0 9.3122775697e-06
Gc29_224 0 n58 ns224 0 1.06394160588e-07
Gc29_225 0 n58 ns225 0 0.00129804057179
Gc29_226 0 n58 ns226 0 -1.74853113586e-05
Gc29_227 0 n58 ns227 0 0.000155244449296
Gc29_228 0 n58 ns228 0 0.000596464713705
Gc29_229 0 n58 ns229 0 -2.56112035058e-05
Gc29_230 0 n58 ns230 0 -8.04123118626e-06
Gc29_231 0 n58 ns231 0 -0.000147089944813
Gc29_232 0 n58 ns232 0 0.000374202178872
Gc29_233 0 n58 ns233 0 -0.000357714451997
Gc29_234 0 n58 ns234 0 8.05045672245e-06
Gc29_235 0 n58 ns235 0 -7.91019302198e-05
Gc29_236 0 n58 ns236 0 -0.000132600918628
Gc29_237 0 n58 ns237 0 -0.000103234520753
Gc29_238 0 n58 ns238 0 -7.02326857493e-05
Gc29_239 0 n58 ns239 0 1.19498718424e-06
Gc29_240 0 n58 ns240 0 -6.29281111419e-05
Gc29_241 0 n58 ns241 0 -0.000302760809671
Gc29_242 0 n58 ns242 0 6.90189005423e-06
Gc29_243 0 n58 ns243 0 -4.31927928537e-05
Gc29_244 0 n58 ns244 0 -6.30382486985e-05
Gc29_245 0 n58 ns245 0 -4.77107280627e-05
Gc29_246 0 n58 ns246 0 -4.39313221041e-06
Gc29_247 0 n58 ns247 0 -8.92273823042e-06
Gc29_248 0 n58 ns248 0 -2.63972193447e-05
Gc29_249 0 n58 ns249 0 2.51431649309e-05
Gc29_250 0 n58 ns250 0 -2.82059674326e-07
Gc29_251 0 n58 ns251 0 3.11587113905e-06
Gc29_252 0 n58 ns252 0 1.22051915095e-06
Gc29_253 0 n58 ns253 0 2.13802733064e-06
Gc29_254 0 n58 ns254 0 6.9233845622e-06
Gc29_255 0 n58 ns255 0 7.65762054461e-07
Gc29_256 0 n58 ns256 0 1.34843742501e-06
Gd29_17 0 n58 ni17 0 -4.53758675177e-06
Gd29_18 0 n58 ni18 0 -3.67400193527e-05
Gd29_19 0 n58 ni19 0 -2.66429824284e-05
Gd29_20 0 n58 ni20 0 0.000266384621423
Gd29_21 0 n58 ni21 0 -0.00120936735797
Gd29_22 0 n58 ni22 0 0.00229255632795
Gd29_23 0 n58 ni23 0 0.00085421845383
Gd29_24 0 n58 ni24 0 9.61544824062e-05
Gd29_25 0 n58 ni25 0 6.37593505202e-07
Gd29_26 0 n58 ni26 0 -5.57271017975e-05
Gd29_27 0 n58 ni27 0 0.000201935722417
Gd29_28 0 n58 ni28 0 0.00015478569166
Gd29_29 0 n58 ni29 0 -0.000972505527827
Gd29_30 0 n58 ni30 0 0.000912475190511
Gd29_31 0 n58 ni31 0 0.000351968411453
Gd29_32 0 n58 ni32 0 -1.68166488884e-05
Gc30_129 0 n60 ns129 0 -1.69827161015e-05
Gc30_130 0 n60 ns130 0 3.59693814167e-07
Gc30_131 0 n60 ns131 0 -2.06151375346e-06
Gc30_132 0 n60 ns132 0 -4.41115606647e-06
Gc30_133 0 n60 ns133 0 -6.33549784162e-06
Gc30_134 0 n60 ns134 0 -6.60134767694e-07
Gc30_135 0 n60 ns135 0 -8.87678411229e-07
Gc30_136 0 n60 ns136 0 -1.27264896543e-06
Gc30_137 0 n60 ns137 0 -1.33355424201e-05
Gc30_138 0 n60 ns138 0 2.91817450727e-07
Gc30_139 0 n60 ns139 0 -1.60742569852e-06
Gc30_140 0 n60 ns140 0 -5.08720653946e-06
Gc30_141 0 n60 ns141 0 -5.64978307588e-06
Gc30_142 0 n60 ns142 0 -8.36443791649e-07
Gc30_143 0 n60 ns143 0 -6.7268816613e-07
Gc30_144 0 n60 ns144 0 -9.47913571328e-07
Gc30_145 0 n60 ns145 0 2.60666358716e-05
Gc30_146 0 n60 ns146 0 -4.51887875034e-07
Gc30_147 0 n60 ns147 0 3.58886350753e-06
Gc30_148 0 n60 ns148 0 -1.08883575176e-06
Gc30_149 0 n60 ns149 0 4.3894775372e-07
Gc30_150 0 n60 ns150 0 2.0404767572e-06
Gc30_151 0 n60 ns151 0 7.75710499288e-07
Gc30_152 0 n60 ns152 0 2.03417517817e-06
Gc30_153 0 n60 ns153 0 1.06417417816e-05
Gc30_154 0 n60 ns154 0 4.49536344769e-08
Gc30_155 0 n60 ns155 0 8.87549088776e-07
Gc30_156 0 n60 ns156 0 -7.92784942294e-06
Gc30_157 0 n60 ns157 0 -2.86039764916e-06
Gc30_158 0 n60 ns158 0 3.62068457176e-06
Gc30_159 0 n60 ns159 0 4.89944621164e-07
Gc30_160 0 n60 ns160 0 2.27252652544e-07
Gc30_161 0 n60 ns161 0 -0.000173215164082
Gc30_162 0 n60 ns162 0 3.18960499216e-06
Gc30_163 0 n60 ns163 0 -2.6785850694e-05
Gc30_164 0 n60 ns164 0 -6.44675872247e-05
Gc30_165 0 n60 ns165 0 -8.34645613861e-05
Gc30_166 0 n60 ns166 0 -4.36229344444e-05
Gc30_167 0 n60 ns167 0 -7.80898851309e-06
Gc30_168 0 n60 ns168 0 -1.59229212503e-05
Gc30_169 0 n60 ns169 0 0.00200150135913
Gc30_170 0 n60 ns170 0 -3.90851185788e-05
Gc30_171 0 n60 ns171 0 0.000170772526484
Gc30_172 0 n60 ns172 0 0.000491206869421
Gc30_173 0 n60 ns173 0 4.18926906033e-05
Gc30_174 0 n60 ns174 0 -1.7047538038e-05
Gc30_175 0 n60 ns175 0 4.09461375119e-05
Gc30_176 0 n60 ns176 0 9.01416772668e-05
Gc30_177 0 n60 ns177 0 0.00129296325347
Gc30_178 0 n60 ns178 0 -1.83063987927e-05
Gc30_179 0 n60 ns179 0 -2.89758585615e-05
Gc30_180 0 n60 ns180 0 0.000370996653914
Gc30_181 0 n60 ns181 0 -6.20836812017e-05
Gc30_182 0 n60 ns182 0 -5.44813082553e-05
Gc30_183 0 n60 ns183 0 4.50852083397e-05
Gc30_184 0 n60 ns184 0 -6.22659363203e-05
Gc30_185 0 n60 ns185 0 -0.000416599261666
Gc30_186 0 n60 ns186 0 8.7272101259e-06
Gc30_187 0 n60 ns187 0 -6.29683440543e-05
Gc30_188 0 n60 ns188 0 -0.000107319559922
Gc30_189 0 n60 ns189 0 -0.000104110516999
Gc30_190 0 n60 ns190 0 -4.45713692311e-05
Gc30_191 0 n60 ns191 0 -1.28187691966e-05
Gc30_192 0 n60 ns192 0 -3.91193847136e-05
Gc30_193 0 n60 ns193 0 1.339020584e-05
Gc30_194 0 n60 ns194 0 5.01568964822e-08
Gc30_195 0 n60 ns195 0 1.58673190283e-06
Gc30_196 0 n60 ns196 0 -7.33827661407e-06
Gc30_197 0 n60 ns197 0 -7.87647664545e-06
Gc30_198 0 n60 ns198 0 6.46051916995e-06
Gc30_199 0 n60 ns199 0 5.87190208233e-08
Gc30_200 0 n60 ns200 0 -1.98930176876e-08
Gc30_201 0 n60 ns201 0 -7.14200261755e-06
Gc30_202 0 n60 ns202 0 2.01916189915e-07
Gc30_203 0 n60 ns203 0 -9.28668116194e-07
Gc30_204 0 n60 ns204 0 -5.57265812495e-06
Gc30_205 0 n60 ns205 0 -3.77867555255e-06
Gc30_206 0 n60 ns206 0 -1.8854878629e-07
Gc30_207 0 n60 ns207 0 -2.62446667277e-07
Gc30_208 0 n60 ns208 0 -5.46261921005e-07
Gc30_209 0 n60 ns209 0 4.1355917412e-05
Gc30_210 0 n60 ns210 0 -6.72047735793e-07
Gc30_211 0 n60 ns211 0 5.43291143996e-06
Gc30_212 0 n60 ns212 0 8.68569192634e-07
Gc30_213 0 n60 ns213 0 2.8317596651e-06
Gc30_214 0 n60 ns214 0 5.07424372759e-06
Gc30_215 0 n60 ns215 0 1.34210249701e-06
Gc30_216 0 n60 ns216 0 2.85041012946e-06
Gc30_217 0 n60 ns217 0 -0.000220325407771
Gc30_218 0 n60 ns218 0 5.04732577646e-06
Gc30_219 0 n60 ns219 0 -3.18589915483e-05
Gc30_220 0 n60 ns220 0 -4.7531801923e-05
Gc30_221 0 n60 ns221 0 -4.08581896209e-05
Gc30_222 0 n60 ns222 0 -4.00906268301e-06
Gc30_223 0 n60 ns223 0 -6.82328725228e-06
Gc30_224 0 n60 ns224 0 -1.99142879207e-05
Gc30_225 0 n60 ns225 0 -0.000357714451997
Gc30_226 0 n60 ns226 0 8.05045672245e-06
Gc30_227 0 n60 ns227 0 -7.91019302198e-05
Gc30_228 0 n60 ns228 0 -0.000132600918628
Gc30_229 0 n60 ns229 0 -0.000103234520753
Gc30_230 0 n60 ns230 0 -7.02326857493e-05
Gc30_231 0 n60 ns231 0 1.19498718424e-06
Gc30_232 0 n60 ns232 0 -6.29281111419e-05
Gc30_233 0 n60 ns233 0 0.00269430294726
Gc30_234 0 n60 ns234 0 -4.61613315894e-05
Gc30_235 0 n60 ns235 0 0.000259563004476
Gc30_236 0 n60 ns236 0 0.000487606116303
Gc30_237 0 n60 ns237 0 0.000194865372243
Gc30_238 0 n60 ns238 0 -0.000113832156712
Gc30_239 0 n60 ns239 0 -2.20507191043e-05
Gc30_240 0 n60 ns240 0 0.000356742992797
Gc30_241 0 n60 ns241 0 0.000239247547721
Gc30_242 0 n60 ns242 0 -5.55237512768e-06
Gc30_243 0 n60 ns243 0 1.06463253619e-05
Gc30_244 0 n60 ns244 0 1.8193197296e-05
Gc30_245 0 n60 ns245 0 -7.94921768874e-05
Gc30_246 0 n60 ns246 0 -6.3314655019e-05
Gc30_247 0 n60 ns247 0 3.63692919042e-06
Gc30_248 0 n60 ns248 0 7.41152804842e-07
Gc30_249 0 n60 ns249 0 -0.000155689908071
Gc30_250 0 n60 ns250 0 3.37922151203e-06
Gc30_251 0 n60 ns251 0 -2.18984569127e-05
Gc30_252 0 n60 ns252 0 -4.70665637267e-05
Gc30_253 0 n60 ns253 0 -4.75150528505e-05
Gc30_254 0 n60 ns254 0 -1.41703497349e-05
Gc30_255 0 n60 ns255 0 -6.02373260463e-06
Gc30_256 0 n60 ns256 0 -1.28758344114e-05
Gd30_17 0 n60 ni17 0 1.63795167917e-05
Gd30_18 0 n60 ni18 0 1.38752198232e-05
Gd30_19 0 n60 ni19 0 -2.21435560549e-05
Gd30_20 0 n60 ni20 0 6.88572029591e-06
Gd30_21 0 n60 ni21 0 0.000274444029911
Gd30_22 0 n60 ni22 0 -0.000341002411723
Gd30_23 0 n60 ni23 0 0.00205758093149
Gd30_24 0 n60 ni24 0 0.00056648777286
Gd30_25 0 n60 ni25 0 2.54085872691e-06
Gd30_26 0 n60 ni26 0 1.05510764412e-05
Gd30_27 0 n60 ni27 0 -3.31026307353e-05
Gd30_28 0 n60 ni28 0 0.000267411405598
Gd30_29 0 n60 ni29 0 0.000912475190511
Gd30_30 0 n60 ni30 0 -0.000892361184715
Gd30_31 0 n60 ni31 0 0.000175135010191
Gd30_32 0 n60 ni32 0 0.000194916344004
Gc31_129 0 n62 ns129 0 -4.40896228817e-06
Gc31_130 0 n62 ns130 0 1.01540444749e-07
Gc31_131 0 n62 ns131 0 -5.04656543256e-07
Gc31_132 0 n62 ns132 0 -1.45244153256e-06
Gc31_133 0 n62 ns133 0 -2.28280679221e-06
Gc31_134 0 n62 ns134 0 1.22043923387e-07
Gc31_135 0 n62 ns135 0 -2.88582963005e-07
Gc31_136 0 n62 ns136 0 -3.41532995247e-07
Gc31_137 0 n62 ns137 0 -6.21514766582e-06
Gc31_138 0 n62 ns138 0 1.36817946084e-07
Gc31_139 0 n62 ns139 0 -7.33781561121e-07
Gc31_140 0 n62 ns140 0 -2.38815207263e-06
Gc31_141 0 n62 ns141 0 -2.83567387845e-06
Gc31_142 0 n62 ns142 0 -2.699612921e-07
Gc31_143 0 n62 ns143 0 -3.37327672664e-07
Gc31_144 0 n62 ns144 0 -4.44846641079e-07
Gc31_145 0 n62 ns145 0 -7.87620638845e-06
Gc31_146 0 n62 ns146 0 1.79741965036e-07
Gc31_147 0 n62 ns147 0 -9.4776889781e-07
Gc31_148 0 n62 ns148 0 -5.50734435248e-06
Gc31_149 0 n62 ns149 0 -3.96035923335e-06
Gc31_150 0 n62 ns150 0 -1.14493889138e-06
Gc31_151 0 n62 ns151 0 -2.98283274329e-07
Gc31_152 0 n62 ns152 0 -4.90177944627e-07
Gc31_153 0 n62 ns153 0 2.41720982126e-05
Gc31_154 0 n62 ns154 0 -4.07348547403e-07
Gc31_155 0 n62 ns155 0 3.21228125022e-06
Gc31_156 0 n62 ns156 0 -2.60139744367e-06
Gc31_157 0 n62 ns157 0 1.30438576621e-06
Gc31_158 0 n62 ns158 0 1.48443556621e-06
Gc31_159 0 n62 ns159 0 9.30459771362e-07
Gc31_160 0 n62 ns160 0 1.89943721576e-06
Gc31_161 0 n62 ns161 0 3.18982930675e-05
Gc31_162 0 n62 ns162 0 -4.60668994107e-07
Gc31_163 0 n62 ns163 0 4.2504089657e-06
Gc31_164 0 n62 ns164 0 -6.23127892136e-06
Gc31_165 0 n62 ns165 0 -4.47765563216e-06
Gc31_166 0 n62 ns166 0 2.56348621427e-06
Gc31_167 0 n62 ns167 0 7.30172313007e-07
Gc31_168 0 n62 ns168 0 2.30131295973e-06
Gc31_169 0 n62 ns169 0 -0.000155117365667
Gc31_170 0 n62 ns170 0 2.60999310966e-06
Gc31_171 0 n62 ns171 0 -2.32484571994e-05
Gc31_172 0 n62 ns172 0 -6.53841012324e-05
Gc31_173 0 n62 ns173 0 -9.18139425139e-05
Gc31_174 0 n62 ns174 0 -5.12667348643e-05
Gc31_175 0 n62 ns175 0 -8.92727097601e-06
Gc31_176 0 n62 ns176 0 -1.18666599177e-05
Gc31_177 0 n62 ns177 0 0.00150170228499
Gc31_178 0 n62 ns178 0 -2.77113772417e-05
Gc31_179 0 n62 ns179 0 9.39328674134e-05
Gc31_180 0 n62 ns180 0 0.000365584014813
Gc31_181 0 n62 ns181 0 8.94566061998e-06
Gc31_182 0 n62 ns182 0 -3.01103714361e-05
Gc31_183 0 n62 ns183 0 3.70497460607e-05
Gc31_184 0 n62 ns184 0 3.73395384038e-05
Gc31_185 0 n62 ns185 0 0.00124437971124
Gc31_186 0 n62 ns186 0 -1.70907301975e-05
Gc31_187 0 n62 ns187 0 -5.76368441398e-05
Gc31_188 0 n62 ns188 0 0.000203442363139
Gc31_189 0 n62 ns189 0 -9.8801839012e-06
Gc31_190 0 n62 ns190 0 -9.11873638941e-05
Gc31_191 0 n62 ns191 0 8.39017295758e-05
Gc31_192 0 n62 ns192 0 -0.000116067609704
Gc31_193 0 n62 ns193 0 -0.000457770310533
Gc31_194 0 n62 ns194 0 9.48035414528e-06
Gc31_195 0 n62 ns195 0 -6.82936761093e-05
Gc31_196 0 n62 ns196 0 -0.000123778383046
Gc31_197 0 n62 ns197 0 -0.000122416962197
Gc31_198 0 n62 ns198 0 -5.23943178946e-05
Gc31_199 0 n62 ns199 0 -1.43754952682e-05
Gc31_200 0 n62 ns200 0 -4.28130746993e-05
Gc31_201 0 n62 ns201 0 -1.12064892543e-05
Gc31_202 0 n62 ns202 0 2.47598106005e-07
Gc31_203 0 n62 ns203 0 -1.44796052741e-06
Gc31_204 0 n62 ns204 0 -4.51788056499e-06
Gc31_205 0 n62 ns205 0 -3.56374876056e-06
Gc31_206 0 n62 ns206 0 -8.33524767247e-07
Gc31_207 0 n62 ns207 0 -4.0589357044e-07
Gc31_208 0 n62 ns208 0 -8.19269843515e-07
Gc31_209 0 n62 ns209 0 1.26588162345e-06
Gc31_210 0 n62 ns210 0 1.97037590375e-08
Gc31_211 0 n62 ns211 0 2.66911264936e-07
Gc31_212 0 n62 ns212 0 -4.72465584684e-06
Gc31_213 0 n62 ns213 0 -3.00456203151e-06
Gc31_214 0 n62 ns214 0 -1.32292346428e-07
Gc31_215 0 n62 ns215 0 -6.04545900447e-09
Gc31_216 0 n62 ns216 0 1.64820160386e-07
Gc31_217 0 n62 ns217 0 4.11707815558e-05
Gc31_218 0 n62 ns218 0 -6.34907008116e-07
Gc31_219 0 n62 ns219 0 5.2283705931e-06
Gc31_220 0 n62 ns220 0 2.25341054598e-06
Gc31_221 0 n62 ns221 0 4.85328957022e-06
Gc31_222 0 n62 ns222 0 6.32853351275e-06
Gc31_223 0 n62 ns223 0 1.44768687659e-06
Gc31_224 0 n62 ns224 0 2.70655127281e-06
Gc31_225 0 n62 ns225 0 -0.000302760809671
Gc31_226 0 n62 ns226 0 6.90189005423e-06
Gc31_227 0 n62 ns227 0 -4.31927928537e-05
Gc31_228 0 n62 ns228 0 -6.30382486985e-05
Gc31_229 0 n62 ns229 0 -4.77107280627e-05
Gc31_230 0 n62 ns230 0 -4.39313221041e-06
Gc31_231 0 n62 ns231 0 -8.92273823042e-06
Gc31_232 0 n62 ns232 0 -2.63972193447e-05
Gc31_233 0 n62 ns233 0 0.000239247547721
Gc31_234 0 n62 ns234 0 -5.55237512768e-06
Gc31_235 0 n62 ns235 0 1.06463253619e-05
Gc31_236 0 n62 ns236 0 1.8193197296e-05
Gc31_237 0 n62 ns237 0 -7.94921768874e-05
Gc31_238 0 n62 ns238 0 -6.3314655019e-05
Gc31_239 0 n62 ns239 0 3.63692919042e-06
Gc31_240 0 n62 ns240 0 7.41152804841e-07
Gc31_241 0 n62 ns241 0 0.00270627018522
Gc31_242 0 n62 ns242 0 -4.64843012389e-05
Gc31_243 0 n62 ns243 0 0.000280434358888
Gc31_244 0 n62 ns244 0 0.000620125251387
Gc31_245 0 n62 ns245 0 0.000162434482363
Gc31_246 0 n62 ns246 0 -7.35723697972e-05
Gc31_247 0 n62 ns247 0 -5.18939151453e-05
Gc31_248 0 n62 ns248 0 0.000395701082466
Gc31_249 0 n62 ns249 0 0.00022721151411
Gc31_250 0 n62 ns250 0 -5.17718445994e-06
Gc31_251 0 n62 ns251 0 8.34330108285e-06
Gc31_252 0 n62 ns252 0 1.60413911386e-05
Gc31_253 0 n62 ns253 0 -7.78581589153e-05
Gc31_254 0 n62 ns254 0 -5.9534358962e-05
Gc31_255 0 n62 ns255 0 4.23420870589e-06
Gc31_256 0 n62 ns256 0 -2.08005604369e-06
Gd31_17 0 n62 ni17 0 4.33983755983e-06
Gd31_18 0 n62 ni18 0 6.35537833744e-06
Gd31_19 0 n62 ni19 0 9.71314523216e-06
Gd31_20 0 n62 ni20 0 -1.84350154855e-05
Gd31_21 0 n62 ni21 0 -1.90454185308e-05
Gd31_22 0 n62 ni22 0 0.000245742976004
Gd31_23 0 n62 ni23 0 0.000310365219524
Gd31_24 0 n62 ni24 0 0.00249515285216
Gd31_25 0 n62 ni25 0 0.000614880238506
Gd31_26 0 n62 ni26 0 1.26247628802e-05
Gd31_27 0 n62 ni27 0 1.6371865763e-06
Gd31_28 0 n62 ni28 0 -3.16853273065e-05
Gd31_29 0 n62 ni29 0 0.000351968411453
Gd31_30 0 n62 ni30 0 0.000175135010191
Gd31_31 0 n62 ni31 0 -0.00124868464243
Gd31_32 0 n62 ni32 0 0.000196918382157
Gc32_129 0 n64 ns129 0 5.47928584667e-08
Gc32_130 0 n64 ns130 0 1.23386166374e-08
Gc32_131 0 n64 ns131 0 1.87981375548e-08
Gc32_132 0 n64 ns132 0 -4.08227354013e-07
Gc32_133 0 n64 ns133 0 -5.29882634366e-07
Gc32_134 0 n64 ns134 0 4.24206541947e-07
Gc32_135 0 n64 ns135 0 -3.83760312087e-08
Gc32_136 0 n64 ns136 0 -2.36854284737e-08
Gc32_137 0 n64 ns137 0 -1.57066795593e-06
Gc32_138 0 n64 ns138 0 4.35766279547e-08
Gc32_139 0 n64 ns139 0 -1.70641176063e-07
Gc32_140 0 n64 ns140 0 -5.68180280887e-07
Gc32_141 0 n64 ns141 0 -1.11537023788e-06
Gc32_142 0 n64 ns142 0 3.34263086421e-07
Gc32_143 0 n64 ns143 0 -1.40862230092e-07
Gc32_144 0 n64 ns144 0 -1.36606983246e-07
Gc32_145 0 n64 ns145 0 -7.00660133042e-06
Gc32_146 0 n64 ns146 0 1.5167016135e-07
Gc32_147 0 n64 ns147 0 -8.20297489284e-07
Gc32_148 0 n64 ns148 0 -2.35232568451e-06
Gc32_149 0 n64 ns149 0 -3.1640734489e-06
Gc32_150 0 n64 ns150 0 -2.66343538937e-07
Gc32_151 0 n64 ns151 0 -4.00116692533e-07
Gc32_152 0 n64 ns152 0 -5.02843839907e-07
Gc32_153 0 n64 ns153 0 -1.00470253424e-05
Gc32_154 0 n64 ns154 0 2.26299914288e-07
Gc32_155 0 n64 ns155 0 -1.23212275319e-06
Gc32_156 0 n64 ns156 0 -5.53469931986e-06
Gc32_157 0 n64 ns157 0 -4.41550244487e-06
Gc32_158 0 n64 ns158 0 -1.05923420368e-06
Gc32_159 0 n64 ns159 0 -4.07754826767e-07
Gc32_160 0 n64 ns160 0 -6.7638426384e-07
Gc32_161 0 n64 ns161 0 3.35154064557e-05
Gc32_162 0 n64 ns162 0 -6.2324267438e-07
Gc32_163 0 n64 ns163 0 4.8413698426e-06
Gc32_164 0 n64 ns164 0 8.80982103685e-07
Gc32_165 0 n64 ns165 0 -8.10236164992e-07
Gc32_166 0 n64 ns166 0 2.51543216331e-06
Gc32_167 0 n64 ns167 0 6.82198892097e-07
Gc32_168 0 n64 ns168 0 2.70054115857e-06
Gc32_169 0 n64 ns169 0 4.67361772516e-05
Gc32_170 0 n64 ns170 0 -8.39908711039e-07
Gc32_171 0 n64 ns171 0 6.66103360451e-06
Gc32_172 0 n64 ns172 0 -5.51356213722e-06
Gc32_173 0 n64 ns173 0 -7.21231675159e-06
Gc32_174 0 n64 ns174 0 8.62277580491e-07
Gc32_175 0 n64 ns175 0 7.54105666793e-07
Gc32_176 0 n64 ns176 0 3.84090475125e-06
Gc32_177 0 n64 ns177 0 -0.000231555473431
Gc32_178 0 n64 ns178 0 4.57349135246e-06
Gc32_179 0 n64 ns179 0 -3.45426840415e-05
Gc32_180 0 n64 ns180 0 -6.68798370633e-05
Gc32_181 0 n64 ns181 0 -8.92243529918e-05
Gc32_182 0 n64 ns182 0 -3.91627588734e-05
Gc32_183 0 n64 ns183 0 -1.04206879445e-05
Gc32_184 0 n64 ns184 0 -2.00611940406e-05
Gc32_185 0 n64 ns185 0 0.00148408529907
Gc32_186 0 n64 ns186 0 -2.7796314362e-05
Gc32_187 0 n64 ns187 0 0.000103661824823
Gc32_188 0 n64 ns188 0 0.000396942021576
Gc32_189 0 n64 ns189 0 -1.59415601016e-05
Gc32_190 0 n64 ns190 0 -2.59341134303e-05
Gc32_191 0 n64 ns191 0 2.40672500713e-05
Gc32_192 0 n64 ns192 0 5.52197315714e-05
Gc32_193 0 n64 ns193 0 0.00187371620734
Gc32_194 0 n64 ns194 0 -3.17497051811e-05
Gc32_195 0 n64 ns195 0 3.07717004615e-05
Gc32_196 0 n64 ns196 0 0.000305336987388
Gc32_197 0 n64 ns197 0 7.70972823382e-06
Gc32_198 0 n64 ns198 0 -0.000112436701004
Gc32_199 0 n64 ns199 0 9.60324222662e-05
Gc32_200 0 n64 ns200 0 -6.15655091428e-05
Gc32_201 0 n64 ns201 0 -4.08222680894e-06
Gc32_202 0 n64 ns202 0 9.63011977173e-08
Gc32_203 0 n64 ns203 0 -5.00258096905e-07
Gc32_204 0 n64 ns204 0 -1.34727374393e-06
Gc32_205 0 n64 ns205 0 -1.7440016758e-06
Gc32_206 0 n64 ns206 0 1.11787171816e-07
Gc32_207 0 n64 ns207 0 -2.26493397531e-07
Gc32_208 0 n64 ns208 0 -3.21301083324e-07
Gc32_209 0 n64 ns209 0 -1.41157795285e-05
Gc32_210 0 n64 ns210 0 3.00381887275e-07
Gc32_211 0 n64 ns211 0 -1.71623590345e-06
Gc32_212 0 n64 ns212 0 -3.95139921113e-06
Gc32_213 0 n64 ns213 0 -5.3040850564e-06
Gc32_214 0 n64 ns214 0 -6.30088140268e-07
Gc32_215 0 n64 ns215 0 -7.28929730822e-07
Gc32_216 0 n64 ns216 0 -1.03753106782e-06
Gc32_217 0 n64 ns217 0 -1.04323121728e-05
Gc32_218 0 n64 ns218 0 2.65625266703e-07
Gc32_219 0 n64 ns219 0 -1.2887555747e-06
Gc32_220 0 n64 ns220 0 -5.49192986133e-06
Gc32_221 0 n64 ns221 0 -5.18261684693e-06
Gc32_222 0 n64 ns222 0 -1.16653793939e-07
Gc32_223 0 n64 ns223 0 -5.19051296579e-07
Gc32_224 0 n64 ns224 0 -8.02298559639e-07
Gc32_225 0 n64 ns225 0 2.51431649309e-05
Gc32_226 0 n64 ns226 0 -2.82059674326e-07
Gc32_227 0 n64 ns227 0 3.11587113905e-06
Gc32_228 0 n64 ns228 0 1.22051915095e-06
Gc32_229 0 n64 ns229 0 2.13802733064e-06
Gc32_230 0 n64 ns230 0 6.9233845622e-06
Gc32_231 0 n64 ns231 0 7.65762054461e-07
Gc32_232 0 n64 ns232 0 1.34843742501e-06
Gc32_233 0 n64 ns233 0 -0.000155689908071
Gc32_234 0 n64 ns234 0 3.37922151203e-06
Gc32_235 0 n64 ns235 0 -2.18984569127e-05
Gc32_236 0 n64 ns236 0 -4.70665637267e-05
Gc32_237 0 n64 ns237 0 -4.75150528505e-05
Gc32_238 0 n64 ns238 0 -1.41703497349e-05
Gc32_239 0 n64 ns239 0 -6.02373260463e-06
Gc32_240 0 n64 ns240 0 -1.28758344114e-05
Gc32_241 0 n64 ns241 0 0.00022721151411
Gc32_242 0 n64 ns242 0 -5.17718445994e-06
Gc32_243 0 n64 ns243 0 8.34330108285e-06
Gc32_244 0 n64 ns244 0 1.60413911386e-05
Gc32_245 0 n64 ns245 0 -7.78581589153e-05
Gc32_246 0 n64 ns246 0 -5.9534358962e-05
Gc32_247 0 n64 ns247 0 4.23420870589e-06
Gc32_248 0 n64 ns248 0 -2.08005604369e-06
Gc32_249 0 n64 ns249 0 0.00243993572499
Gc32_250 0 n64 ns250 0 -4.03758899864e-05
Gc32_251 0 n64 ns251 0 0.000229365982974
Gc32_252 0 n64 ns252 0 0.000545535065575
Gc32_253 0 n64 ns253 0 0.000118046928444
Gc32_254 0 n64 ns254 0 -9.61741256901e-05
Gc32_255 0 n64 ns255 0 -5.1386239511e-05
Gc32_256 0 n64 ns256 0 0.000354297930429
Gd32_17 0 n64 ni17 0 3.63182731526e-07
Gd32_18 0 n64 ni18 0 1.65374822263e-06
Gd32_19 0 n64 ni19 0 6.86507352528e-06
Gd32_20 0 n64 ni20 0 1.1690764446e-05
Gd32_21 0 n64 ni21 0 -3.25757267317e-05
Gd32_22 0 n64 ni22 0 -3.71823980704e-05
Gd32_23 0 n64 ni23 0 0.000327283176686
Gd32_24 0 n64 ni24 0 0.000130833325332
Gd32_25 0 n64 ni25 0 0.00184398665632
Gd32_26 0 n64 ni26 0 4.33959101293e-06
Gd32_27 0 n64 ni27 0 1.38176184722e-05
Gd32_28 0 n64 ni28 0 1.27444282105e-05
Gd32_29 0 n64 ni29 0 -1.68166488884e-05
Gd32_30 0 n64 ni30 0 0.000194916344004
Gd32_31 0 n64 ni31 0 0.000196918382157
Gd32_32 0 n64 ni32 0 -0.000722006019578
.ends m16lines_port_fws
