* BEGIN ANSOFT HEADER
* node 1    trace_p_0_T1
* node 2    trace_n_0_T1
* node 3    trace_p_1_T1
* node 4    trace_n_1_T1
* node 5    trace_p_0_T2
* node 6    trace_n_0_T2
* node 7    trace_p_1_T2
* node 8    trace_n_1_T2
*   Format: HSPICE
*   Topckt: m4lines_HFSS_fws
*     Date: Wed Jun 03 22:25:34 2020
*    Notes: Frequency range: 1e+08 to 7e+10 Hz, 700 points
*         : Maximum number of poles: 10000
*         : S-Matrix fitting error tolerance: 0.001
*         : Causality check tolerance: auto
*         : Passivity enforcement: on (by iterated fitting)
*         : Causality enforcement: off
*         : Fitting method: FastFit
*         : Matrix fitting: By entire matrix (required by FastFit)
*         : Ensure Z-parameter accuracy: on
*         : Relative error control: off
*         : Common ground option: on
*         : Final fitting error: 0.002983
*         : Final model order: 296
* END ANSOFT HEADER

.subckt m4lines_HFSS_fws 1 2 3 4 5 6 7 8
Vam1 1 n2 dc 0
Rport1 n2 0 50 noise=0
Vam2 2 n4 dc 0
Rport2 n4 0 50 noise=0
Vam3 3 n6 dc 0
Rport3 n6 0 50 noise=0
Vam4 4 n8 dc 0
Rport4 n8 0 50 noise=0
Vam5 5 n10 dc 0
Rport5 n10 0 50 noise=0
Vam6 6 n12 dc 0
Rport6 n12 0 50 noise=0
Vam7 7 n14 dc 0
Rport7 n14 0 50 noise=0
Vam8 8 n16 dc 0
Rport8 n16 0 50 noise=0

Fi1 0 ni1 Vam1 50
Gi1 0 ni1 1 0 1
Rt1 ni1 0 1 noise=0
Fi2 0 ni2 Vam2 50
Gi2 0 ni2 2 0 1
Rt2 ni2 0 1 noise=0
Fi3 0 ni3 Vam3 50
Gi3 0 ni3 3 0 1
Rt3 ni3 0 1 noise=0
Fi4 0 ni4 Vam4 50
Gi4 0 ni4 4 0 1
Rt4 ni4 0 1 noise=0
Fi5 0 ni5 Vam5 50
Gi5 0 ni5 5 0 1
Rt5 ni5 0 1 noise=0
Fi6 0 ni6 Vam6 50
Gi6 0 ni6 6 0 1
Rt6 ni6 0 1 noise=0
Fi7 0 ni7 Vam7 50
Gi7 0 ni7 7 0 1
Rt7 ni7 0 1 noise=0
Fi8 0 ni8 Vam8 50
Gi8 0 ni8 8 0 1
Rt8 ni8 0 1 noise=0

Ca1 ns1 0 1e-12
Ra1 ns1 0 1.00629317801 noise=0
Ca2 ns2 0 1e-12
Ca3 ns3 0 1e-12
Ra2 ns2 0 3.23514518726 noise=0
Ra3 ns3 0 3.23514518726 noise=0
Ga2 ns2 0 ns3 0 -0.496444529287
Ga3 ns3 0 ns2 0 0.496444529287
Ca4 ns4 0 1e-12
Ca5 ns5 0 1e-12
Ra4 ns4 0 99.2967616202 noise=0
Ra5 ns5 0 99.2967616202 noise=0
Ga4 ns4 0 ns5 0 -0.503988242707
Ga5 ns5 0 ns4 0 0.503988242707
Ca6 ns6 0 1e-12
Ca7 ns7 0 1e-12
Ra6 ns6 0 46.6813218836 noise=0
Ra7 ns7 0 46.6813218836 noise=0
Ga6 ns6 0 ns7 0 -0.489302368603
Ga7 ns7 0 ns6 0 0.489302368603
Ca8 ns8 0 1e-12
Ca9 ns9 0 1e-12
Ra8 ns8 0 34.9646419918 noise=0
Ra9 ns9 0 34.9646419918 noise=0
Ga8 ns8 0 ns9 0 -0.465240916059
Ga9 ns9 0 ns8 0 0.465240916059
Ca10 ns10 0 1e-12
Ca11 ns11 0 1e-12
Ra10 ns10 0 30.2486203037 noise=0
Ra11 ns11 0 30.2486203037 noise=0
Ga10 ns10 0 ns11 0 -0.433297630249
Ga11 ns11 0 ns10 0 0.433297630249
Ca12 ns12 0 1e-12
Ca13 ns13 0 1e-12
Ra12 ns12 0 20.2165502189 noise=0
Ra13 ns13 0 20.2165502189 noise=0
Ga12 ns12 0 ns13 0 -0.415689448636
Ga13 ns13 0 ns12 0 0.415689448636
Ca14 ns14 0 1e-12
Ca15 ns15 0 1e-12
Ra14 ns14 0 40.8940460192 noise=0
Ra15 ns15 0 40.8940460192 noise=0
Ga14 ns14 0 ns15 0 -0.385147744818
Ga15 ns15 0 ns14 0 0.385147744818
Ca16 ns16 0 1e-12
Ca17 ns17 0 1e-12
Ra16 ns16 0 19.9117226261 noise=0
Ra17 ns17 0 19.9117226261 noise=0
Ga16 ns16 0 ns17 0 -0.346186931449
Ga17 ns17 0 ns16 0 0.346186931449
Ca18 ns18 0 1e-12
Ca19 ns19 0 1e-12
Ra18 ns18 0 22.383359742 noise=0
Ra19 ns19 0 22.383359742 noise=0
Ga18 ns18 0 ns19 0 -0.317452973336
Ga19 ns19 0 ns18 0 0.317452973336
Ca20 ns20 0 1e-12
Ca21 ns21 0 1e-12
Ra20 ns20 0 38.0479358576 noise=0
Ra21 ns21 0 38.0479358576 noise=0
Ga20 ns20 0 ns21 0 -0.29186865188
Ga21 ns21 0 ns20 0 0.29186865188
Ca22 ns22 0 1e-12
Ca23 ns23 0 1e-12
Ra22 ns22 0 12.4189583497 noise=0
Ra23 ns23 0 12.4189583497 noise=0
Ga22 ns22 0 ns23 0 -0.258059325384
Ga23 ns23 0 ns22 0 0.258059325384
Ca24 ns24 0 1e-12
Ca25 ns25 0 1e-12
Ra24 ns24 0 23.0324462867 noise=0
Ra25 ns25 0 23.0324462867 noise=0
Ga24 ns24 0 ns25 0 -0.212645067874
Ga25 ns25 0 ns24 0 0.212645067874
Ca26 ns26 0 1e-12
Ca27 ns27 0 1e-12
Ra26 ns26 0 34.7188374441 noise=0
Ra27 ns27 0 34.7188374441 noise=0
Ga26 ns26 0 ns27 0 -0.19740480044
Ga27 ns27 0 ns26 0 0.19740480044
Ca28 ns28 0 1e-12
Ca29 ns29 0 1e-12
Ra28 ns28 0 13.2633244371 noise=0
Ra29 ns29 0 13.2633244371 noise=0
Ga28 ns28 0 ns29 0 -0.121026208723
Ga29 ns29 0 ns28 0 0.121026208723
Ca30 ns30 0 1e-12
Ca31 ns31 0 1e-12
Ra30 ns30 0 18.9661932554 noise=0
Ra31 ns31 0 18.9661932554 noise=0
Ga30 ns30 0 ns31 0 -0.10544020576
Ga31 ns31 0 ns30 0 0.10544020576
Ca32 ns32 0 1e-12
Ca33 ns33 0 1e-12
Ra32 ns32 0 32.7496561073 noise=0
Ra33 ns33 0 32.7496561073 noise=0
Ga32 ns32 0 ns33 0 -0.100351912105
Ga33 ns33 0 ns32 0 0.100351912105
Ca34 ns34 0 1e-12
Ra34 ns34 0 24.8522946037 noise=0
Ca35 ns35 0 1e-12
Ca36 ns36 0 1e-12
Ra35 ns35 0 27.1312266605 noise=0
Ra36 ns36 0 27.1312266605 noise=0
Ga35 ns35 0 ns36 0 -0.0077220911993
Ga36 ns36 0 ns35 0 0.0077220911993
Ca37 ns37 0 1e-12
Ra37 ns37 0 1255.41863382 noise=0
Ca38 ns38 0 1e-12
Ra38 ns38 0 1.00629317801 noise=0
Ca39 ns39 0 1e-12
Ca40 ns40 0 1e-12
Ra39 ns39 0 3.23514518726 noise=0
Ra40 ns40 0 3.23514518726 noise=0
Ga39 ns39 0 ns40 0 -0.496444529287
Ga40 ns40 0 ns39 0 0.496444529287
Ca41 ns41 0 1e-12
Ca42 ns42 0 1e-12
Ra41 ns41 0 99.2967616202 noise=0
Ra42 ns42 0 99.2967616202 noise=0
Ga41 ns41 0 ns42 0 -0.503988242707
Ga42 ns42 0 ns41 0 0.503988242707
Ca43 ns43 0 1e-12
Ca44 ns44 0 1e-12
Ra43 ns43 0 46.6813218836 noise=0
Ra44 ns44 0 46.6813218836 noise=0
Ga43 ns43 0 ns44 0 -0.489302368603
Ga44 ns44 0 ns43 0 0.489302368603
Ca45 ns45 0 1e-12
Ca46 ns46 0 1e-12
Ra45 ns45 0 34.9646419918 noise=0
Ra46 ns46 0 34.9646419918 noise=0
Ga45 ns45 0 ns46 0 -0.465240916059
Ga46 ns46 0 ns45 0 0.465240916059
Ca47 ns47 0 1e-12
Ca48 ns48 0 1e-12
Ra47 ns47 0 30.2486203037 noise=0
Ra48 ns48 0 30.2486203037 noise=0
Ga47 ns47 0 ns48 0 -0.433297630249
Ga48 ns48 0 ns47 0 0.433297630249
Ca49 ns49 0 1e-12
Ca50 ns50 0 1e-12
Ra49 ns49 0 20.2165502189 noise=0
Ra50 ns50 0 20.2165502189 noise=0
Ga49 ns49 0 ns50 0 -0.415689448636
Ga50 ns50 0 ns49 0 0.415689448636
Ca51 ns51 0 1e-12
Ca52 ns52 0 1e-12
Ra51 ns51 0 40.8940460192 noise=0
Ra52 ns52 0 40.8940460192 noise=0
Ga51 ns51 0 ns52 0 -0.385147744818
Ga52 ns52 0 ns51 0 0.385147744818
Ca53 ns53 0 1e-12
Ca54 ns54 0 1e-12
Ra53 ns53 0 19.9117226261 noise=0
Ra54 ns54 0 19.9117226261 noise=0
Ga53 ns53 0 ns54 0 -0.346186931449
Ga54 ns54 0 ns53 0 0.346186931449
Ca55 ns55 0 1e-12
Ca56 ns56 0 1e-12
Ra55 ns55 0 22.383359742 noise=0
Ra56 ns56 0 22.383359742 noise=0
Ga55 ns55 0 ns56 0 -0.317452973336
Ga56 ns56 0 ns55 0 0.317452973336
Ca57 ns57 0 1e-12
Ca58 ns58 0 1e-12
Ra57 ns57 0 38.0479358576 noise=0
Ra58 ns58 0 38.0479358576 noise=0
Ga57 ns57 0 ns58 0 -0.29186865188
Ga58 ns58 0 ns57 0 0.29186865188
Ca59 ns59 0 1e-12
Ca60 ns60 0 1e-12
Ra59 ns59 0 12.4189583497 noise=0
Ra60 ns60 0 12.4189583497 noise=0
Ga59 ns59 0 ns60 0 -0.258059325384
Ga60 ns60 0 ns59 0 0.258059325384
Ca61 ns61 0 1e-12
Ca62 ns62 0 1e-12
Ra61 ns61 0 23.0324462867 noise=0
Ra62 ns62 0 23.0324462867 noise=0
Ga61 ns61 0 ns62 0 -0.212645067874
Ga62 ns62 0 ns61 0 0.212645067874
Ca63 ns63 0 1e-12
Ca64 ns64 0 1e-12
Ra63 ns63 0 34.7188374441 noise=0
Ra64 ns64 0 34.7188374441 noise=0
Ga63 ns63 0 ns64 0 -0.19740480044
Ga64 ns64 0 ns63 0 0.19740480044
Ca65 ns65 0 1e-12
Ca66 ns66 0 1e-12
Ra65 ns65 0 13.2633244371 noise=0
Ra66 ns66 0 13.2633244371 noise=0
Ga65 ns65 0 ns66 0 -0.121026208723
Ga66 ns66 0 ns65 0 0.121026208723
Ca67 ns67 0 1e-12
Ca68 ns68 0 1e-12
Ra67 ns67 0 18.9661932554 noise=0
Ra68 ns68 0 18.9661932554 noise=0
Ga67 ns67 0 ns68 0 -0.10544020576
Ga68 ns68 0 ns67 0 0.10544020576
Ca69 ns69 0 1e-12
Ca70 ns70 0 1e-12
Ra69 ns69 0 32.7496561073 noise=0
Ra70 ns70 0 32.7496561073 noise=0
Ga69 ns69 0 ns70 0 -0.100351912105
Ga70 ns70 0 ns69 0 0.100351912105
Ca71 ns71 0 1e-12
Ra71 ns71 0 24.8522946037 noise=0
Ca72 ns72 0 1e-12
Ca73 ns73 0 1e-12
Ra72 ns72 0 27.1312266605 noise=0
Ra73 ns73 0 27.1312266605 noise=0
Ga72 ns72 0 ns73 0 -0.0077220911993
Ga73 ns73 0 ns72 0 0.0077220911993
Ca74 ns74 0 1e-12
Ra74 ns74 0 1255.41863382 noise=0
Ca75 ns75 0 1e-12
Ra75 ns75 0 1.00629317801 noise=0
Ca76 ns76 0 1e-12
Ca77 ns77 0 1e-12
Ra76 ns76 0 3.23514518726 noise=0
Ra77 ns77 0 3.23514518726 noise=0
Ga76 ns76 0 ns77 0 -0.496444529287
Ga77 ns77 0 ns76 0 0.496444529287
Ca78 ns78 0 1e-12
Ca79 ns79 0 1e-12
Ra78 ns78 0 99.2967616202 noise=0
Ra79 ns79 0 99.2967616202 noise=0
Ga78 ns78 0 ns79 0 -0.503988242707
Ga79 ns79 0 ns78 0 0.503988242707
Ca80 ns80 0 1e-12
Ca81 ns81 0 1e-12
Ra80 ns80 0 46.6813218836 noise=0
Ra81 ns81 0 46.6813218836 noise=0
Ga80 ns80 0 ns81 0 -0.489302368603
Ga81 ns81 0 ns80 0 0.489302368603
Ca82 ns82 0 1e-12
Ca83 ns83 0 1e-12
Ra82 ns82 0 34.9646419918 noise=0
Ra83 ns83 0 34.9646419918 noise=0
Ga82 ns82 0 ns83 0 -0.465240916059
Ga83 ns83 0 ns82 0 0.465240916059
Ca84 ns84 0 1e-12
Ca85 ns85 0 1e-12
Ra84 ns84 0 30.2486203037 noise=0
Ra85 ns85 0 30.2486203037 noise=0
Ga84 ns84 0 ns85 0 -0.433297630249
Ga85 ns85 0 ns84 0 0.433297630249
Ca86 ns86 0 1e-12
Ca87 ns87 0 1e-12
Ra86 ns86 0 20.2165502189 noise=0
Ra87 ns87 0 20.2165502189 noise=0
Ga86 ns86 0 ns87 0 -0.415689448636
Ga87 ns87 0 ns86 0 0.415689448636
Ca88 ns88 0 1e-12
Ca89 ns89 0 1e-12
Ra88 ns88 0 40.8940460192 noise=0
Ra89 ns89 0 40.8940460192 noise=0
Ga88 ns88 0 ns89 0 -0.385147744818
Ga89 ns89 0 ns88 0 0.385147744818
Ca90 ns90 0 1e-12
Ca91 ns91 0 1e-12
Ra90 ns90 0 19.9117226261 noise=0
Ra91 ns91 0 19.9117226261 noise=0
Ga90 ns90 0 ns91 0 -0.346186931449
Ga91 ns91 0 ns90 0 0.346186931449
Ca92 ns92 0 1e-12
Ca93 ns93 0 1e-12
Ra92 ns92 0 22.383359742 noise=0
Ra93 ns93 0 22.383359742 noise=0
Ga92 ns92 0 ns93 0 -0.317452973336
Ga93 ns93 0 ns92 0 0.317452973336
Ca94 ns94 0 1e-12
Ca95 ns95 0 1e-12
Ra94 ns94 0 38.0479358576 noise=0
Ra95 ns95 0 38.0479358576 noise=0
Ga94 ns94 0 ns95 0 -0.29186865188
Ga95 ns95 0 ns94 0 0.29186865188
Ca96 ns96 0 1e-12
Ca97 ns97 0 1e-12
Ra96 ns96 0 12.4189583497 noise=0
Ra97 ns97 0 12.4189583497 noise=0
Ga96 ns96 0 ns97 0 -0.258059325384
Ga97 ns97 0 ns96 0 0.258059325384
Ca98 ns98 0 1e-12
Ca99 ns99 0 1e-12
Ra98 ns98 0 23.0324462867 noise=0
Ra99 ns99 0 23.0324462867 noise=0
Ga98 ns98 0 ns99 0 -0.212645067874
Ga99 ns99 0 ns98 0 0.212645067874
Ca100 ns100 0 1e-12
Ca101 ns101 0 1e-12
Ra100 ns100 0 34.7188374441 noise=0
Ra101 ns101 0 34.7188374441 noise=0
Ga100 ns100 0 ns101 0 -0.19740480044
Ga101 ns101 0 ns100 0 0.19740480044
Ca102 ns102 0 1e-12
Ca103 ns103 0 1e-12
Ra102 ns102 0 13.2633244371 noise=0
Ra103 ns103 0 13.2633244371 noise=0
Ga102 ns102 0 ns103 0 -0.121026208723
Ga103 ns103 0 ns102 0 0.121026208723
Ca104 ns104 0 1e-12
Ca105 ns105 0 1e-12
Ra104 ns104 0 18.9661932554 noise=0
Ra105 ns105 0 18.9661932554 noise=0
Ga104 ns104 0 ns105 0 -0.10544020576
Ga105 ns105 0 ns104 0 0.10544020576
Ca106 ns106 0 1e-12
Ca107 ns107 0 1e-12
Ra106 ns106 0 32.7496561073 noise=0
Ra107 ns107 0 32.7496561073 noise=0
Ga106 ns106 0 ns107 0 -0.100351912105
Ga107 ns107 0 ns106 0 0.100351912105
Ca108 ns108 0 1e-12
Ra108 ns108 0 24.8522946037 noise=0
Ca109 ns109 0 1e-12
Ca110 ns110 0 1e-12
Ra109 ns109 0 27.1312266605 noise=0
Ra110 ns110 0 27.1312266605 noise=0
Ga109 ns109 0 ns110 0 -0.0077220911993
Ga110 ns110 0 ns109 0 0.0077220911993
Ca111 ns111 0 1e-12
Ra111 ns111 0 1255.41863382 noise=0
Ca112 ns112 0 1e-12
Ra112 ns112 0 1.00629317801 noise=0
Ca113 ns113 0 1e-12
Ca114 ns114 0 1e-12
Ra113 ns113 0 3.23514518726 noise=0
Ra114 ns114 0 3.23514518726 noise=0
Ga113 ns113 0 ns114 0 -0.496444529287
Ga114 ns114 0 ns113 0 0.496444529287
Ca115 ns115 0 1e-12
Ca116 ns116 0 1e-12
Ra115 ns115 0 99.2967616202 noise=0
Ra116 ns116 0 99.2967616202 noise=0
Ga115 ns115 0 ns116 0 -0.503988242707
Ga116 ns116 0 ns115 0 0.503988242707
Ca117 ns117 0 1e-12
Ca118 ns118 0 1e-12
Ra117 ns117 0 46.6813218836 noise=0
Ra118 ns118 0 46.6813218836 noise=0
Ga117 ns117 0 ns118 0 -0.489302368603
Ga118 ns118 0 ns117 0 0.489302368603
Ca119 ns119 0 1e-12
Ca120 ns120 0 1e-12
Ra119 ns119 0 34.9646419918 noise=0
Ra120 ns120 0 34.9646419918 noise=0
Ga119 ns119 0 ns120 0 -0.465240916059
Ga120 ns120 0 ns119 0 0.465240916059
Ca121 ns121 0 1e-12
Ca122 ns122 0 1e-12
Ra121 ns121 0 30.2486203037 noise=0
Ra122 ns122 0 30.2486203037 noise=0
Ga121 ns121 0 ns122 0 -0.433297630249
Ga122 ns122 0 ns121 0 0.433297630249
Ca123 ns123 0 1e-12
Ca124 ns124 0 1e-12
Ra123 ns123 0 20.2165502189 noise=0
Ra124 ns124 0 20.2165502189 noise=0
Ga123 ns123 0 ns124 0 -0.415689448636
Ga124 ns124 0 ns123 0 0.415689448636
Ca125 ns125 0 1e-12
Ca126 ns126 0 1e-12
Ra125 ns125 0 40.8940460192 noise=0
Ra126 ns126 0 40.8940460192 noise=0
Ga125 ns125 0 ns126 0 -0.385147744818
Ga126 ns126 0 ns125 0 0.385147744818
Ca127 ns127 0 1e-12
Ca128 ns128 0 1e-12
Ra127 ns127 0 19.9117226261 noise=0
Ra128 ns128 0 19.9117226261 noise=0
Ga127 ns127 0 ns128 0 -0.346186931449
Ga128 ns128 0 ns127 0 0.346186931449
Ca129 ns129 0 1e-12
Ca130 ns130 0 1e-12
Ra129 ns129 0 22.383359742 noise=0
Ra130 ns130 0 22.383359742 noise=0
Ga129 ns129 0 ns130 0 -0.317452973336
Ga130 ns130 0 ns129 0 0.317452973336
Ca131 ns131 0 1e-12
Ca132 ns132 0 1e-12
Ra131 ns131 0 38.0479358576 noise=0
Ra132 ns132 0 38.0479358576 noise=0
Ga131 ns131 0 ns132 0 -0.29186865188
Ga132 ns132 0 ns131 0 0.29186865188
Ca133 ns133 0 1e-12
Ca134 ns134 0 1e-12
Ra133 ns133 0 12.4189583497 noise=0
Ra134 ns134 0 12.4189583497 noise=0
Ga133 ns133 0 ns134 0 -0.258059325384
Ga134 ns134 0 ns133 0 0.258059325384
Ca135 ns135 0 1e-12
Ca136 ns136 0 1e-12
Ra135 ns135 0 23.0324462867 noise=0
Ra136 ns136 0 23.0324462867 noise=0
Ga135 ns135 0 ns136 0 -0.212645067874
Ga136 ns136 0 ns135 0 0.212645067874
Ca137 ns137 0 1e-12
Ca138 ns138 0 1e-12
Ra137 ns137 0 34.7188374441 noise=0
Ra138 ns138 0 34.7188374441 noise=0
Ga137 ns137 0 ns138 0 -0.19740480044
Ga138 ns138 0 ns137 0 0.19740480044
Ca139 ns139 0 1e-12
Ca140 ns140 0 1e-12
Ra139 ns139 0 13.2633244371 noise=0
Ra140 ns140 0 13.2633244371 noise=0
Ga139 ns139 0 ns140 0 -0.121026208723
Ga140 ns140 0 ns139 0 0.121026208723
Ca141 ns141 0 1e-12
Ca142 ns142 0 1e-12
Ra141 ns141 0 18.9661932554 noise=0
Ra142 ns142 0 18.9661932554 noise=0
Ga141 ns141 0 ns142 0 -0.10544020576
Ga142 ns142 0 ns141 0 0.10544020576
Ca143 ns143 0 1e-12
Ca144 ns144 0 1e-12
Ra143 ns143 0 32.7496561073 noise=0
Ra144 ns144 0 32.7496561073 noise=0
Ga143 ns143 0 ns144 0 -0.100351912105
Ga144 ns144 0 ns143 0 0.100351912105
Ca145 ns145 0 1e-12
Ra145 ns145 0 24.8522946037 noise=0
Ca146 ns146 0 1e-12
Ca147 ns147 0 1e-12
Ra146 ns146 0 27.1312266605 noise=0
Ra147 ns147 0 27.1312266605 noise=0
Ga146 ns146 0 ns147 0 -0.0077220911993
Ga147 ns147 0 ns146 0 0.0077220911993
Ca148 ns148 0 1e-12
Ra148 ns148 0 1255.41863382 noise=0
Ca149 ns149 0 1e-12
Ra149 ns149 0 1.00629317801 noise=0
Ca150 ns150 0 1e-12
Ca151 ns151 0 1e-12
Ra150 ns150 0 3.23514518726 noise=0
Ra151 ns151 0 3.23514518726 noise=0
Ga150 ns150 0 ns151 0 -0.496444529287
Ga151 ns151 0 ns150 0 0.496444529287
Ca152 ns152 0 1e-12
Ca153 ns153 0 1e-12
Ra152 ns152 0 99.2967616202 noise=0
Ra153 ns153 0 99.2967616202 noise=0
Ga152 ns152 0 ns153 0 -0.503988242707
Ga153 ns153 0 ns152 0 0.503988242707
Ca154 ns154 0 1e-12
Ca155 ns155 0 1e-12
Ra154 ns154 0 46.6813218836 noise=0
Ra155 ns155 0 46.6813218836 noise=0
Ga154 ns154 0 ns155 0 -0.489302368603
Ga155 ns155 0 ns154 0 0.489302368603
Ca156 ns156 0 1e-12
Ca157 ns157 0 1e-12
Ra156 ns156 0 34.9646419918 noise=0
Ra157 ns157 0 34.9646419918 noise=0
Ga156 ns156 0 ns157 0 -0.465240916059
Ga157 ns157 0 ns156 0 0.465240916059
Ca158 ns158 0 1e-12
Ca159 ns159 0 1e-12
Ra158 ns158 0 30.2486203037 noise=0
Ra159 ns159 0 30.2486203037 noise=0
Ga158 ns158 0 ns159 0 -0.433297630249
Ga159 ns159 0 ns158 0 0.433297630249
Ca160 ns160 0 1e-12
Ca161 ns161 0 1e-12
Ra160 ns160 0 20.2165502189 noise=0
Ra161 ns161 0 20.2165502189 noise=0
Ga160 ns160 0 ns161 0 -0.415689448636
Ga161 ns161 0 ns160 0 0.415689448636
Ca162 ns162 0 1e-12
Ca163 ns163 0 1e-12
Ra162 ns162 0 40.8940460192 noise=0
Ra163 ns163 0 40.8940460192 noise=0
Ga162 ns162 0 ns163 0 -0.385147744818
Ga163 ns163 0 ns162 0 0.385147744818
Ca164 ns164 0 1e-12
Ca165 ns165 0 1e-12
Ra164 ns164 0 19.9117226261 noise=0
Ra165 ns165 0 19.9117226261 noise=0
Ga164 ns164 0 ns165 0 -0.346186931449
Ga165 ns165 0 ns164 0 0.346186931449
Ca166 ns166 0 1e-12
Ca167 ns167 0 1e-12
Ra166 ns166 0 22.383359742 noise=0
Ra167 ns167 0 22.383359742 noise=0
Ga166 ns166 0 ns167 0 -0.317452973336
Ga167 ns167 0 ns166 0 0.317452973336
Ca168 ns168 0 1e-12
Ca169 ns169 0 1e-12
Ra168 ns168 0 38.0479358576 noise=0
Ra169 ns169 0 38.0479358576 noise=0
Ga168 ns168 0 ns169 0 -0.29186865188
Ga169 ns169 0 ns168 0 0.29186865188
Ca170 ns170 0 1e-12
Ca171 ns171 0 1e-12
Ra170 ns170 0 12.4189583497 noise=0
Ra171 ns171 0 12.4189583497 noise=0
Ga170 ns170 0 ns171 0 -0.258059325384
Ga171 ns171 0 ns170 0 0.258059325384
Ca172 ns172 0 1e-12
Ca173 ns173 0 1e-12
Ra172 ns172 0 23.0324462867 noise=0
Ra173 ns173 0 23.0324462867 noise=0
Ga172 ns172 0 ns173 0 -0.212645067874
Ga173 ns173 0 ns172 0 0.212645067874
Ca174 ns174 0 1e-12
Ca175 ns175 0 1e-12
Ra174 ns174 0 34.7188374441 noise=0
Ra175 ns175 0 34.7188374441 noise=0
Ga174 ns174 0 ns175 0 -0.19740480044
Ga175 ns175 0 ns174 0 0.19740480044
Ca176 ns176 0 1e-12
Ca177 ns177 0 1e-12
Ra176 ns176 0 13.2633244371 noise=0
Ra177 ns177 0 13.2633244371 noise=0
Ga176 ns176 0 ns177 0 -0.121026208723
Ga177 ns177 0 ns176 0 0.121026208723
Ca178 ns178 0 1e-12
Ca179 ns179 0 1e-12
Ra178 ns178 0 18.9661932554 noise=0
Ra179 ns179 0 18.9661932554 noise=0
Ga178 ns178 0 ns179 0 -0.10544020576
Ga179 ns179 0 ns178 0 0.10544020576
Ca180 ns180 0 1e-12
Ca181 ns181 0 1e-12
Ra180 ns180 0 32.7496561073 noise=0
Ra181 ns181 0 32.7496561073 noise=0
Ga180 ns180 0 ns181 0 -0.100351912105
Ga181 ns181 0 ns180 0 0.100351912105
Ca182 ns182 0 1e-12
Ra182 ns182 0 24.8522946037 noise=0
Ca183 ns183 0 1e-12
Ca184 ns184 0 1e-12
Ra183 ns183 0 27.1312266605 noise=0
Ra184 ns184 0 27.1312266605 noise=0
Ga183 ns183 0 ns184 0 -0.0077220911993
Ga184 ns184 0 ns183 0 0.0077220911993
Ca185 ns185 0 1e-12
Ra185 ns185 0 1255.41863382 noise=0
Ca186 ns186 0 1e-12
Ra186 ns186 0 1.00629317801 noise=0
Ca187 ns187 0 1e-12
Ca188 ns188 0 1e-12
Ra187 ns187 0 3.23514518726 noise=0
Ra188 ns188 0 3.23514518726 noise=0
Ga187 ns187 0 ns188 0 -0.496444529287
Ga188 ns188 0 ns187 0 0.496444529287
Ca189 ns189 0 1e-12
Ca190 ns190 0 1e-12
Ra189 ns189 0 99.2967616202 noise=0
Ra190 ns190 0 99.2967616202 noise=0
Ga189 ns189 0 ns190 0 -0.503988242707
Ga190 ns190 0 ns189 0 0.503988242707
Ca191 ns191 0 1e-12
Ca192 ns192 0 1e-12
Ra191 ns191 0 46.6813218836 noise=0
Ra192 ns192 0 46.6813218836 noise=0
Ga191 ns191 0 ns192 0 -0.489302368603
Ga192 ns192 0 ns191 0 0.489302368603
Ca193 ns193 0 1e-12
Ca194 ns194 0 1e-12
Ra193 ns193 0 34.9646419918 noise=0
Ra194 ns194 0 34.9646419918 noise=0
Ga193 ns193 0 ns194 0 -0.465240916059
Ga194 ns194 0 ns193 0 0.465240916059
Ca195 ns195 0 1e-12
Ca196 ns196 0 1e-12
Ra195 ns195 0 30.2486203037 noise=0
Ra196 ns196 0 30.2486203037 noise=0
Ga195 ns195 0 ns196 0 -0.433297630249
Ga196 ns196 0 ns195 0 0.433297630249
Ca197 ns197 0 1e-12
Ca198 ns198 0 1e-12
Ra197 ns197 0 20.2165502189 noise=0
Ra198 ns198 0 20.2165502189 noise=0
Ga197 ns197 0 ns198 0 -0.415689448636
Ga198 ns198 0 ns197 0 0.415689448636
Ca199 ns199 0 1e-12
Ca200 ns200 0 1e-12
Ra199 ns199 0 40.8940460192 noise=0
Ra200 ns200 0 40.8940460192 noise=0
Ga199 ns199 0 ns200 0 -0.385147744818
Ga200 ns200 0 ns199 0 0.385147744818
Ca201 ns201 0 1e-12
Ca202 ns202 0 1e-12
Ra201 ns201 0 19.9117226261 noise=0
Ra202 ns202 0 19.9117226261 noise=0
Ga201 ns201 0 ns202 0 -0.346186931449
Ga202 ns202 0 ns201 0 0.346186931449
Ca203 ns203 0 1e-12
Ca204 ns204 0 1e-12
Ra203 ns203 0 22.383359742 noise=0
Ra204 ns204 0 22.383359742 noise=0
Ga203 ns203 0 ns204 0 -0.317452973336
Ga204 ns204 0 ns203 0 0.317452973336
Ca205 ns205 0 1e-12
Ca206 ns206 0 1e-12
Ra205 ns205 0 38.0479358576 noise=0
Ra206 ns206 0 38.0479358576 noise=0
Ga205 ns205 0 ns206 0 -0.29186865188
Ga206 ns206 0 ns205 0 0.29186865188
Ca207 ns207 0 1e-12
Ca208 ns208 0 1e-12
Ra207 ns207 0 12.4189583497 noise=0
Ra208 ns208 0 12.4189583497 noise=0
Ga207 ns207 0 ns208 0 -0.258059325384
Ga208 ns208 0 ns207 0 0.258059325384
Ca209 ns209 0 1e-12
Ca210 ns210 0 1e-12
Ra209 ns209 0 23.0324462867 noise=0
Ra210 ns210 0 23.0324462867 noise=0
Ga209 ns209 0 ns210 0 -0.212645067874
Ga210 ns210 0 ns209 0 0.212645067874
Ca211 ns211 0 1e-12
Ca212 ns212 0 1e-12
Ra211 ns211 0 34.7188374441 noise=0
Ra212 ns212 0 34.7188374441 noise=0
Ga211 ns211 0 ns212 0 -0.19740480044
Ga212 ns212 0 ns211 0 0.19740480044
Ca213 ns213 0 1e-12
Ca214 ns214 0 1e-12
Ra213 ns213 0 13.2633244371 noise=0
Ra214 ns214 0 13.2633244371 noise=0
Ga213 ns213 0 ns214 0 -0.121026208723
Ga214 ns214 0 ns213 0 0.121026208723
Ca215 ns215 0 1e-12
Ca216 ns216 0 1e-12
Ra215 ns215 0 18.9661932554 noise=0
Ra216 ns216 0 18.9661932554 noise=0
Ga215 ns215 0 ns216 0 -0.10544020576
Ga216 ns216 0 ns215 0 0.10544020576
Ca217 ns217 0 1e-12
Ca218 ns218 0 1e-12
Ra217 ns217 0 32.7496561073 noise=0
Ra218 ns218 0 32.7496561073 noise=0
Ga217 ns217 0 ns218 0 -0.100351912105
Ga218 ns218 0 ns217 0 0.100351912105
Ca219 ns219 0 1e-12
Ra219 ns219 0 24.8522946037 noise=0
Ca220 ns220 0 1e-12
Ca221 ns221 0 1e-12
Ra220 ns220 0 27.1312266605 noise=0
Ra221 ns221 0 27.1312266605 noise=0
Ga220 ns220 0 ns221 0 -0.0077220911993
Ga221 ns221 0 ns220 0 0.0077220911993
Ca222 ns222 0 1e-12
Ra222 ns222 0 1255.41863382 noise=0
Ca223 ns223 0 1e-12
Ra223 ns223 0 1.00629317801 noise=0
Ca224 ns224 0 1e-12
Ca225 ns225 0 1e-12
Ra224 ns224 0 3.23514518726 noise=0
Ra225 ns225 0 3.23514518726 noise=0
Ga224 ns224 0 ns225 0 -0.496444529287
Ga225 ns225 0 ns224 0 0.496444529287
Ca226 ns226 0 1e-12
Ca227 ns227 0 1e-12
Ra226 ns226 0 99.2967616202 noise=0
Ra227 ns227 0 99.2967616202 noise=0
Ga226 ns226 0 ns227 0 -0.503988242707
Ga227 ns227 0 ns226 0 0.503988242707
Ca228 ns228 0 1e-12
Ca229 ns229 0 1e-12
Ra228 ns228 0 46.6813218836 noise=0
Ra229 ns229 0 46.6813218836 noise=0
Ga228 ns228 0 ns229 0 -0.489302368603
Ga229 ns229 0 ns228 0 0.489302368603
Ca230 ns230 0 1e-12
Ca231 ns231 0 1e-12
Ra230 ns230 0 34.9646419918 noise=0
Ra231 ns231 0 34.9646419918 noise=0
Ga230 ns230 0 ns231 0 -0.465240916059
Ga231 ns231 0 ns230 0 0.465240916059
Ca232 ns232 0 1e-12
Ca233 ns233 0 1e-12
Ra232 ns232 0 30.2486203037 noise=0
Ra233 ns233 0 30.2486203037 noise=0
Ga232 ns232 0 ns233 0 -0.433297630249
Ga233 ns233 0 ns232 0 0.433297630249
Ca234 ns234 0 1e-12
Ca235 ns235 0 1e-12
Ra234 ns234 0 20.2165502189 noise=0
Ra235 ns235 0 20.2165502189 noise=0
Ga234 ns234 0 ns235 0 -0.415689448636
Ga235 ns235 0 ns234 0 0.415689448636
Ca236 ns236 0 1e-12
Ca237 ns237 0 1e-12
Ra236 ns236 0 40.8940460192 noise=0
Ra237 ns237 0 40.8940460192 noise=0
Ga236 ns236 0 ns237 0 -0.385147744818
Ga237 ns237 0 ns236 0 0.385147744818
Ca238 ns238 0 1e-12
Ca239 ns239 0 1e-12
Ra238 ns238 0 19.9117226261 noise=0
Ra239 ns239 0 19.9117226261 noise=0
Ga238 ns238 0 ns239 0 -0.346186931449
Ga239 ns239 0 ns238 0 0.346186931449
Ca240 ns240 0 1e-12
Ca241 ns241 0 1e-12
Ra240 ns240 0 22.383359742 noise=0
Ra241 ns241 0 22.383359742 noise=0
Ga240 ns240 0 ns241 0 -0.317452973336
Ga241 ns241 0 ns240 0 0.317452973336
Ca242 ns242 0 1e-12
Ca243 ns243 0 1e-12
Ra242 ns242 0 38.0479358576 noise=0
Ra243 ns243 0 38.0479358576 noise=0
Ga242 ns242 0 ns243 0 -0.29186865188
Ga243 ns243 0 ns242 0 0.29186865188
Ca244 ns244 0 1e-12
Ca245 ns245 0 1e-12
Ra244 ns244 0 12.4189583497 noise=0
Ra245 ns245 0 12.4189583497 noise=0
Ga244 ns244 0 ns245 0 -0.258059325384
Ga245 ns245 0 ns244 0 0.258059325384
Ca246 ns246 0 1e-12
Ca247 ns247 0 1e-12
Ra246 ns246 0 23.0324462867 noise=0
Ra247 ns247 0 23.0324462867 noise=0
Ga246 ns246 0 ns247 0 -0.212645067874
Ga247 ns247 0 ns246 0 0.212645067874
Ca248 ns248 0 1e-12
Ca249 ns249 0 1e-12
Ra248 ns248 0 34.7188374441 noise=0
Ra249 ns249 0 34.7188374441 noise=0
Ga248 ns248 0 ns249 0 -0.19740480044
Ga249 ns249 0 ns248 0 0.19740480044
Ca250 ns250 0 1e-12
Ca251 ns251 0 1e-12
Ra250 ns250 0 13.2633244371 noise=0
Ra251 ns251 0 13.2633244371 noise=0
Ga250 ns250 0 ns251 0 -0.121026208723
Ga251 ns251 0 ns250 0 0.121026208723
Ca252 ns252 0 1e-12
Ca253 ns253 0 1e-12
Ra252 ns252 0 18.9661932554 noise=0
Ra253 ns253 0 18.9661932554 noise=0
Ga252 ns252 0 ns253 0 -0.10544020576
Ga253 ns253 0 ns252 0 0.10544020576
Ca254 ns254 0 1e-12
Ca255 ns255 0 1e-12
Ra254 ns254 0 32.7496561073 noise=0
Ra255 ns255 0 32.7496561073 noise=0
Ga254 ns254 0 ns255 0 -0.100351912105
Ga255 ns255 0 ns254 0 0.100351912105
Ca256 ns256 0 1e-12
Ra256 ns256 0 24.8522946037 noise=0
Ca257 ns257 0 1e-12
Ca258 ns258 0 1e-12
Ra257 ns257 0 27.1312266605 noise=0
Ra258 ns258 0 27.1312266605 noise=0
Ga257 ns257 0 ns258 0 -0.0077220911993
Ga258 ns258 0 ns257 0 0.0077220911993
Ca259 ns259 0 1e-12
Ra259 ns259 0 1255.41863382 noise=0
Ca260 ns260 0 1e-12
Ra260 ns260 0 1.00629317801 noise=0
Ca261 ns261 0 1e-12
Ca262 ns262 0 1e-12
Ra261 ns261 0 3.23514518726 noise=0
Ra262 ns262 0 3.23514518726 noise=0
Ga261 ns261 0 ns262 0 -0.496444529287
Ga262 ns262 0 ns261 0 0.496444529287
Ca263 ns263 0 1e-12
Ca264 ns264 0 1e-12
Ra263 ns263 0 99.2967616202 noise=0
Ra264 ns264 0 99.2967616202 noise=0
Ga263 ns263 0 ns264 0 -0.503988242707
Ga264 ns264 0 ns263 0 0.503988242707
Ca265 ns265 0 1e-12
Ca266 ns266 0 1e-12
Ra265 ns265 0 46.6813218836 noise=0
Ra266 ns266 0 46.6813218836 noise=0
Ga265 ns265 0 ns266 0 -0.489302368603
Ga266 ns266 0 ns265 0 0.489302368603
Ca267 ns267 0 1e-12
Ca268 ns268 0 1e-12
Ra267 ns267 0 34.9646419918 noise=0
Ra268 ns268 0 34.9646419918 noise=0
Ga267 ns267 0 ns268 0 -0.465240916059
Ga268 ns268 0 ns267 0 0.465240916059
Ca269 ns269 0 1e-12
Ca270 ns270 0 1e-12
Ra269 ns269 0 30.2486203037 noise=0
Ra270 ns270 0 30.2486203037 noise=0
Ga269 ns269 0 ns270 0 -0.433297630249
Ga270 ns270 0 ns269 0 0.433297630249
Ca271 ns271 0 1e-12
Ca272 ns272 0 1e-12
Ra271 ns271 0 20.2165502189 noise=0
Ra272 ns272 0 20.2165502189 noise=0
Ga271 ns271 0 ns272 0 -0.415689448636
Ga272 ns272 0 ns271 0 0.415689448636
Ca273 ns273 0 1e-12
Ca274 ns274 0 1e-12
Ra273 ns273 0 40.8940460192 noise=0
Ra274 ns274 0 40.8940460192 noise=0
Ga273 ns273 0 ns274 0 -0.385147744818
Ga274 ns274 0 ns273 0 0.385147744818
Ca275 ns275 0 1e-12
Ca276 ns276 0 1e-12
Ra275 ns275 0 19.9117226261 noise=0
Ra276 ns276 0 19.9117226261 noise=0
Ga275 ns275 0 ns276 0 -0.346186931449
Ga276 ns276 0 ns275 0 0.346186931449
Ca277 ns277 0 1e-12
Ca278 ns278 0 1e-12
Ra277 ns277 0 22.383359742 noise=0
Ra278 ns278 0 22.383359742 noise=0
Ga277 ns277 0 ns278 0 -0.317452973336
Ga278 ns278 0 ns277 0 0.317452973336
Ca279 ns279 0 1e-12
Ca280 ns280 0 1e-12
Ra279 ns279 0 38.0479358576 noise=0
Ra280 ns280 0 38.0479358576 noise=0
Ga279 ns279 0 ns280 0 -0.29186865188
Ga280 ns280 0 ns279 0 0.29186865188
Ca281 ns281 0 1e-12
Ca282 ns282 0 1e-12
Ra281 ns281 0 12.4189583497 noise=0
Ra282 ns282 0 12.4189583497 noise=0
Ga281 ns281 0 ns282 0 -0.258059325384
Ga282 ns282 0 ns281 0 0.258059325384
Ca283 ns283 0 1e-12
Ca284 ns284 0 1e-12
Ra283 ns283 0 23.0324462867 noise=0
Ra284 ns284 0 23.0324462867 noise=0
Ga283 ns283 0 ns284 0 -0.212645067874
Ga284 ns284 0 ns283 0 0.212645067874
Ca285 ns285 0 1e-12
Ca286 ns286 0 1e-12
Ra285 ns285 0 34.7188374441 noise=0
Ra286 ns286 0 34.7188374441 noise=0
Ga285 ns285 0 ns286 0 -0.19740480044
Ga286 ns286 0 ns285 0 0.19740480044
Ca287 ns287 0 1e-12
Ca288 ns288 0 1e-12
Ra287 ns287 0 13.2633244371 noise=0
Ra288 ns288 0 13.2633244371 noise=0
Ga287 ns287 0 ns288 0 -0.121026208723
Ga288 ns288 0 ns287 0 0.121026208723
Ca289 ns289 0 1e-12
Ca290 ns290 0 1e-12
Ra289 ns289 0 18.9661932554 noise=0
Ra290 ns290 0 18.9661932554 noise=0
Ga289 ns289 0 ns290 0 -0.10544020576
Ga290 ns290 0 ns289 0 0.10544020576
Ca291 ns291 0 1e-12
Ca292 ns292 0 1e-12
Ra291 ns291 0 32.7496561073 noise=0
Ra292 ns292 0 32.7496561073 noise=0
Ga291 ns291 0 ns292 0 -0.100351912105
Ga292 ns292 0 ns291 0 0.100351912105
Ca293 ns293 0 1e-12
Ra293 ns293 0 24.8522946037 noise=0
Ca294 ns294 0 1e-12
Ca295 ns295 0 1e-12
Ra294 ns294 0 27.1312266605 noise=0
Ra295 ns295 0 27.1312266605 noise=0
Ga294 ns294 0 ns295 0 -0.0077220911993
Ga295 ns295 0 ns294 0 0.0077220911993
Ca296 ns296 0 1e-12
Ra296 ns296 0 1255.41863382 noise=0

Gb1_1 ns1 0 ni1 0 -0.993746178399
Gb2_1 ns2 0 ni1 0 0.206357749572
Gb3_1 ns3 0 ni1 0 0.560418939038
Gb4_1 ns4 0 ni1 0 -0.0439373586586
Gb5_1 ns5 0 ni1 0 -0.503311512913
Gb6_1 ns6 0 ni1 0 0.484702471978
Gb7_1 ns7 0 ni1 0 0.126489377174
Gb8_1 ns8 0 ni1 0 -0.154502502487
Gb9_1 ns9 0 ni1 0 0.45750117795
Gb10_1 ns10 0 ni1 0 0.239858010195
Gb11_1 ns11 0 ni1 0 0.417519489808
Gb12_1 ns12 0 ni1 0 0.364442397777
Gb13_1 ns13 0 ni1 0 -0.378209055662
Gb14_1 ns14 0 ni1 0 -0.290550143198
Gb15_1 ns15 0 ni1 0 0.36825298363
Gb16_1 ns16 0 ni1 0 0.138172492565
Gb17_1 ns17 0 ni1 0 0.333427821107
Gb18_1 ns18 0 ni1 0 -0.284467134658
Gb19_1 ns19 0 ni1 0 0.279062335386
Gb20_1 ns20 0 ni1 0 -0.0902629370133
Gb21_1 ns21 0 ni1 0 0.286107255774
Gb22_1 ns22 0 ni1 0 0.28041018527
Gb23_1 ns23 0 ni1 0 0.00889138929927
Gb24_1 ns24 0 ni1 0 0.186356489801
Gb25_1 ns25 0 ni1 0 -0.172171530087
Gb26_1 ns26 0 ni1 0 -0.0714391928051
Gb27_1 ns27 0 ni1 0 0.191183839252
Gb28_1 ns28 0 ni1 0 0.106816939055
Gb29_1 ns29 0 ni1 0 0.09820473861
Gb30_1 ns30 0 ni1 0 -0.114955578665
Gb31_1 ns31 0 ni1 0 0.0336965571042
Gb32_1 ns32 0 ni1 0 -0.0933250056251
Gb33_1 ns33 0 ni1 0 0.0536285339485
Gb34_1 ns34 0 ni1 0 -0.0402377332133
Gb35_1 ns35 0 ni1 0 0.00827411543063
Gb36_1 ns36 0 ni1 0 -0.0367422440678
Gb37_1 ns37 0 ni1 0 0.000796547042602
Gb38_2 ns38 0 ni2 0 -0.993746178399
Gb39_2 ns39 0 ni2 0 0.206357749572
Gb40_2 ns40 0 ni2 0 0.560418939038
Gb41_2 ns41 0 ni2 0 -0.0439373586586
Gb42_2 ns42 0 ni2 0 -0.503311512913
Gb43_2 ns43 0 ni2 0 0.484702471978
Gb44_2 ns44 0 ni2 0 0.126489377174
Gb45_2 ns45 0 ni2 0 -0.154502502487
Gb46_2 ns46 0 ni2 0 0.45750117795
Gb47_2 ns47 0 ni2 0 0.239858010195
Gb48_2 ns48 0 ni2 0 0.417519489808
Gb49_2 ns49 0 ni2 0 0.364442397777
Gb50_2 ns50 0 ni2 0 -0.378209055662
Gb51_2 ns51 0 ni2 0 -0.290550143198
Gb52_2 ns52 0 ni2 0 0.36825298363
Gb53_2 ns53 0 ni2 0 0.138172492565
Gb54_2 ns54 0 ni2 0 0.333427821107
Gb55_2 ns55 0 ni2 0 -0.284467134658
Gb56_2 ns56 0 ni2 0 0.279062335386
Gb57_2 ns57 0 ni2 0 -0.0902629370133
Gb58_2 ns58 0 ni2 0 0.286107255774
Gb59_2 ns59 0 ni2 0 0.28041018527
Gb60_2 ns60 0 ni2 0 0.00889138929927
Gb61_2 ns61 0 ni2 0 0.186356489801
Gb62_2 ns62 0 ni2 0 -0.172171530087
Gb63_2 ns63 0 ni2 0 -0.0714391928051
Gb64_2 ns64 0 ni2 0 0.191183839252
Gb65_2 ns65 0 ni2 0 0.106816939055
Gb66_2 ns66 0 ni2 0 0.09820473861
Gb67_2 ns67 0 ni2 0 -0.114955578665
Gb68_2 ns68 0 ni2 0 0.0336965571042
Gb69_2 ns69 0 ni2 0 -0.0933250056251
Gb70_2 ns70 0 ni2 0 0.0536285339485
Gb71_2 ns71 0 ni2 0 -0.0402377332133
Gb72_2 ns72 0 ni2 0 0.00827411543063
Gb73_2 ns73 0 ni2 0 -0.0367422440678
Gb74_2 ns74 0 ni2 0 0.000796547042602
Gb75_3 ns75 0 ni3 0 -0.993746178399
Gb76_3 ns76 0 ni3 0 0.206357749572
Gb77_3 ns77 0 ni3 0 0.560418939038
Gb78_3 ns78 0 ni3 0 -0.0439373586586
Gb79_3 ns79 0 ni3 0 -0.503311512913
Gb80_3 ns80 0 ni3 0 0.484702471978
Gb81_3 ns81 0 ni3 0 0.126489377174
Gb82_3 ns82 0 ni3 0 -0.154502502487
Gb83_3 ns83 0 ni3 0 0.45750117795
Gb84_3 ns84 0 ni3 0 0.239858010195
Gb85_3 ns85 0 ni3 0 0.417519489808
Gb86_3 ns86 0 ni3 0 0.364442397777
Gb87_3 ns87 0 ni3 0 -0.378209055662
Gb88_3 ns88 0 ni3 0 -0.290550143198
Gb89_3 ns89 0 ni3 0 0.36825298363
Gb90_3 ns90 0 ni3 0 0.138172492565
Gb91_3 ns91 0 ni3 0 0.333427821107
Gb92_3 ns92 0 ni3 0 -0.284467134658
Gb93_3 ns93 0 ni3 0 0.279062335386
Gb94_3 ns94 0 ni3 0 -0.0902629370133
Gb95_3 ns95 0 ni3 0 0.286107255774
Gb96_3 ns96 0 ni3 0 0.28041018527
Gb97_3 ns97 0 ni3 0 0.00889138929927
Gb98_3 ns98 0 ni3 0 0.186356489801
Gb99_3 ns99 0 ni3 0 -0.172171530087
Gb100_3 ns100 0 ni3 0 -0.0714391928051
Gb101_3 ns101 0 ni3 0 0.191183839252
Gb102_3 ns102 0 ni3 0 0.106816939055
Gb103_3 ns103 0 ni3 0 0.09820473861
Gb104_3 ns104 0 ni3 0 -0.114955578665
Gb105_3 ns105 0 ni3 0 0.0336965571042
Gb106_3 ns106 0 ni3 0 -0.0933250056251
Gb107_3 ns107 0 ni3 0 0.0536285339485
Gb108_3 ns108 0 ni3 0 -0.0402377332133
Gb109_3 ns109 0 ni3 0 0.00827411543063
Gb110_3 ns110 0 ni3 0 -0.0367422440678
Gb111_3 ns111 0 ni3 0 0.000796547042602
Gb112_4 ns112 0 ni4 0 -0.993746178399
Gb113_4 ns113 0 ni4 0 0.206357749572
Gb114_4 ns114 0 ni4 0 0.560418939038
Gb115_4 ns115 0 ni4 0 -0.0439373586586
Gb116_4 ns116 0 ni4 0 -0.503311512913
Gb117_4 ns117 0 ni4 0 0.484702471978
Gb118_4 ns118 0 ni4 0 0.126489377174
Gb119_4 ns119 0 ni4 0 -0.154502502487
Gb120_4 ns120 0 ni4 0 0.45750117795
Gb121_4 ns121 0 ni4 0 0.239858010195
Gb122_4 ns122 0 ni4 0 0.417519489808
Gb123_4 ns123 0 ni4 0 0.364442397777
Gb124_4 ns124 0 ni4 0 -0.378209055662
Gb125_4 ns125 0 ni4 0 -0.290550143198
Gb126_4 ns126 0 ni4 0 0.36825298363
Gb127_4 ns127 0 ni4 0 0.138172492565
Gb128_4 ns128 0 ni4 0 0.333427821107
Gb129_4 ns129 0 ni4 0 -0.284467134658
Gb130_4 ns130 0 ni4 0 0.279062335386
Gb131_4 ns131 0 ni4 0 -0.0902629370133
Gb132_4 ns132 0 ni4 0 0.286107255774
Gb133_4 ns133 0 ni4 0 0.28041018527
Gb134_4 ns134 0 ni4 0 0.00889138929927
Gb135_4 ns135 0 ni4 0 0.186356489801
Gb136_4 ns136 0 ni4 0 -0.172171530087
Gb137_4 ns137 0 ni4 0 -0.0714391928051
Gb138_4 ns138 0 ni4 0 0.191183839252
Gb139_4 ns139 0 ni4 0 0.106816939055
Gb140_4 ns140 0 ni4 0 0.09820473861
Gb141_4 ns141 0 ni4 0 -0.114955578665
Gb142_4 ns142 0 ni4 0 0.0336965571042
Gb143_4 ns143 0 ni4 0 -0.0933250056251
Gb144_4 ns144 0 ni4 0 0.0536285339485
Gb145_4 ns145 0 ni4 0 -0.0402377332133
Gb146_4 ns146 0 ni4 0 0.00827411543063
Gb147_4 ns147 0 ni4 0 -0.0367422440678
Gb148_4 ns148 0 ni4 0 0.000796547042602
Gb149_5 ns149 0 ni5 0 -0.993746178399
Gb150_5 ns150 0 ni5 0 0.206357749572
Gb151_5 ns151 0 ni5 0 0.560418939038
Gb152_5 ns152 0 ni5 0 -0.0439373586586
Gb153_5 ns153 0 ni5 0 -0.503311512913
Gb154_5 ns154 0 ni5 0 0.484702471978
Gb155_5 ns155 0 ni5 0 0.126489377174
Gb156_5 ns156 0 ni5 0 -0.154502502487
Gb157_5 ns157 0 ni5 0 0.45750117795
Gb158_5 ns158 0 ni5 0 0.239858010195
Gb159_5 ns159 0 ni5 0 0.417519489808
Gb160_5 ns160 0 ni5 0 0.364442397777
Gb161_5 ns161 0 ni5 0 -0.378209055662
Gb162_5 ns162 0 ni5 0 -0.290550143198
Gb163_5 ns163 0 ni5 0 0.36825298363
Gb164_5 ns164 0 ni5 0 0.138172492565
Gb165_5 ns165 0 ni5 0 0.333427821107
Gb166_5 ns166 0 ni5 0 -0.284467134658
Gb167_5 ns167 0 ni5 0 0.279062335386
Gb168_5 ns168 0 ni5 0 -0.0902629370133
Gb169_5 ns169 0 ni5 0 0.286107255774
Gb170_5 ns170 0 ni5 0 0.28041018527
Gb171_5 ns171 0 ni5 0 0.00889138929927
Gb172_5 ns172 0 ni5 0 0.186356489801
Gb173_5 ns173 0 ni5 0 -0.172171530087
Gb174_5 ns174 0 ni5 0 -0.0714391928051
Gb175_5 ns175 0 ni5 0 0.191183839252
Gb176_5 ns176 0 ni5 0 0.106816939055
Gb177_5 ns177 0 ni5 0 0.09820473861
Gb178_5 ns178 0 ni5 0 -0.114955578665
Gb179_5 ns179 0 ni5 0 0.0336965571042
Gb180_5 ns180 0 ni5 0 -0.0933250056251
Gb181_5 ns181 0 ni5 0 0.0536285339485
Gb182_5 ns182 0 ni5 0 -0.0402377332133
Gb183_5 ns183 0 ni5 0 0.00827411543063
Gb184_5 ns184 0 ni5 0 -0.0367422440678
Gb185_5 ns185 0 ni5 0 0.000796547042602
Gb186_6 ns186 0 ni6 0 -0.993746178399
Gb187_6 ns187 0 ni6 0 0.206357749572
Gb188_6 ns188 0 ni6 0 0.560418939038
Gb189_6 ns189 0 ni6 0 -0.0439373586586
Gb190_6 ns190 0 ni6 0 -0.503311512913
Gb191_6 ns191 0 ni6 0 0.484702471978
Gb192_6 ns192 0 ni6 0 0.126489377174
Gb193_6 ns193 0 ni6 0 -0.154502502487
Gb194_6 ns194 0 ni6 0 0.45750117795
Gb195_6 ns195 0 ni6 0 0.239858010195
Gb196_6 ns196 0 ni6 0 0.417519489808
Gb197_6 ns197 0 ni6 0 0.364442397777
Gb198_6 ns198 0 ni6 0 -0.378209055662
Gb199_6 ns199 0 ni6 0 -0.290550143198
Gb200_6 ns200 0 ni6 0 0.36825298363
Gb201_6 ns201 0 ni6 0 0.138172492565
Gb202_6 ns202 0 ni6 0 0.333427821107
Gb203_6 ns203 0 ni6 0 -0.284467134658
Gb204_6 ns204 0 ni6 0 0.279062335386
Gb205_6 ns205 0 ni6 0 -0.0902629370133
Gb206_6 ns206 0 ni6 0 0.286107255774
Gb207_6 ns207 0 ni6 0 0.28041018527
Gb208_6 ns208 0 ni6 0 0.00889138929927
Gb209_6 ns209 0 ni6 0 0.186356489801
Gb210_6 ns210 0 ni6 0 -0.172171530087
Gb211_6 ns211 0 ni6 0 -0.0714391928051
Gb212_6 ns212 0 ni6 0 0.191183839252
Gb213_6 ns213 0 ni6 0 0.106816939055
Gb214_6 ns214 0 ni6 0 0.09820473861
Gb215_6 ns215 0 ni6 0 -0.114955578665
Gb216_6 ns216 0 ni6 0 0.0336965571042
Gb217_6 ns217 0 ni6 0 -0.0933250056251
Gb218_6 ns218 0 ni6 0 0.0536285339485
Gb219_6 ns219 0 ni6 0 -0.0402377332133
Gb220_6 ns220 0 ni6 0 0.00827411543063
Gb221_6 ns221 0 ni6 0 -0.0367422440678
Gb222_6 ns222 0 ni6 0 0.000796547042602
Gb223_7 ns223 0 ni7 0 -0.993746178399
Gb224_7 ns224 0 ni7 0 0.206357749572
Gb225_7 ns225 0 ni7 0 0.560418939038
Gb226_7 ns226 0 ni7 0 -0.0439373586586
Gb227_7 ns227 0 ni7 0 -0.503311512913
Gb228_7 ns228 0 ni7 0 0.484702471978
Gb229_7 ns229 0 ni7 0 0.126489377174
Gb230_7 ns230 0 ni7 0 -0.154502502487
Gb231_7 ns231 0 ni7 0 0.45750117795
Gb232_7 ns232 0 ni7 0 0.239858010195
Gb233_7 ns233 0 ni7 0 0.417519489808
Gb234_7 ns234 0 ni7 0 0.364442397777
Gb235_7 ns235 0 ni7 0 -0.378209055662
Gb236_7 ns236 0 ni7 0 -0.290550143198
Gb237_7 ns237 0 ni7 0 0.36825298363
Gb238_7 ns238 0 ni7 0 0.138172492565
Gb239_7 ns239 0 ni7 0 0.333427821107
Gb240_7 ns240 0 ni7 0 -0.284467134658
Gb241_7 ns241 0 ni7 0 0.279062335386
Gb242_7 ns242 0 ni7 0 -0.0902629370133
Gb243_7 ns243 0 ni7 0 0.286107255774
Gb244_7 ns244 0 ni7 0 0.28041018527
Gb245_7 ns245 0 ni7 0 0.00889138929927
Gb246_7 ns246 0 ni7 0 0.186356489801
Gb247_7 ns247 0 ni7 0 -0.172171530087
Gb248_7 ns248 0 ni7 0 -0.0714391928051
Gb249_7 ns249 0 ni7 0 0.191183839252
Gb250_7 ns250 0 ni7 0 0.106816939055
Gb251_7 ns251 0 ni7 0 0.09820473861
Gb252_7 ns252 0 ni7 0 -0.114955578665
Gb253_7 ns253 0 ni7 0 0.0336965571042
Gb254_7 ns254 0 ni7 0 -0.0933250056251
Gb255_7 ns255 0 ni7 0 0.0536285339485
Gb256_7 ns256 0 ni7 0 -0.0402377332133
Gb257_7 ns257 0 ni7 0 0.00827411543063
Gb258_7 ns258 0 ni7 0 -0.0367422440678
Gb259_7 ns259 0 ni7 0 0.000796547042602
Gb260_8 ns260 0 ni8 0 -0.993746178399
Gb261_8 ns261 0 ni8 0 0.206357749572
Gb262_8 ns262 0 ni8 0 0.560418939038
Gb263_8 ns263 0 ni8 0 -0.0439373586586
Gb264_8 ns264 0 ni8 0 -0.503311512913
Gb265_8 ns265 0 ni8 0 0.484702471978
Gb266_8 ns266 0 ni8 0 0.126489377174
Gb267_8 ns267 0 ni8 0 -0.154502502487
Gb268_8 ns268 0 ni8 0 0.45750117795
Gb269_8 ns269 0 ni8 0 0.239858010195
Gb270_8 ns270 0 ni8 0 0.417519489808
Gb271_8 ns271 0 ni8 0 0.364442397777
Gb272_8 ns272 0 ni8 0 -0.378209055662
Gb273_8 ns273 0 ni8 0 -0.290550143198
Gb274_8 ns274 0 ni8 0 0.36825298363
Gb275_8 ns275 0 ni8 0 0.138172492565
Gb276_8 ns276 0 ni8 0 0.333427821107
Gb277_8 ns277 0 ni8 0 -0.284467134658
Gb278_8 ns278 0 ni8 0 0.279062335386
Gb279_8 ns279 0 ni8 0 -0.0902629370133
Gb280_8 ns280 0 ni8 0 0.286107255774
Gb281_8 ns281 0 ni8 0 0.28041018527
Gb282_8 ns282 0 ni8 0 0.00889138929927
Gb283_8 ns283 0 ni8 0 0.186356489801
Gb284_8 ns284 0 ni8 0 -0.172171530087
Gb285_8 ns285 0 ni8 0 -0.0714391928051
Gb286_8 ns286 0 ni8 0 0.191183839252
Gb287_8 ns287 0 ni8 0 0.106816939055
Gb288_8 ns288 0 ni8 0 0.09820473861
Gb289_8 ns289 0 ni8 0 -0.114955578665
Gb290_8 ns290 0 ni8 0 0.0336965571042
Gb291_8 ns291 0 ni8 0 -0.0933250056251
Gb292_8 ns292 0 ni8 0 0.0536285339485
Gb293_8 ns293 0 ni8 0 -0.0402377332133
Gb294_8 ns294 0 ni8 0 0.00827411543063
Gb295_8 ns295 0 ni8 0 -0.0367422440678
Gb296_8 ns296 0 ni8 0 0.000796547042602

Gc1_1 0 n2 ns1 0 0.0108132308795
Gc1_2 0 n2 ns2 0 0.000717611845537
Gc1_3 0 n2 ns3 0 -0.00107372007532
Gc1_4 0 n2 ns4 0 1.3977760174e-06
Gc1_5 0 n2 ns5 0 5.47531978417e-06
Gc1_6 0 n2 ns6 0 0.00011839545812
Gc1_7 0 n2 ns7 0 3.14147048651e-05
Gc1_8 0 n2 ns8 0 -0.000421077801281
Gc1_9 0 n2 ns9 0 7.18097129447e-06
Gc1_10 0 n2 ns10 0 0.000540632090045
Gc1_11 0 n2 ns11 0 -0.000207074360606
Gc1_12 0 n2 ns12 0 0.000782657861359
Gc1_13 0 n2 ns13 0 -0.000311701936873
Gc1_14 0 n2 ns14 0 -0.000204052541882
Gc1_15 0 n2 ns15 0 0.000284880988559
Gc1_16 0 n2 ns16 0 0.000659377884754
Gc1_17 0 n2 ns17 0 -0.00150383602312
Gc1_18 0 n2 ns18 0 -0.00126206325369
Gc1_19 0 n2 ns19 0 0.00075695560162
Gc1_20 0 n2 ns20 0 -0.000143538828107
Gc1_21 0 n2 ns21 0 0.000712263736893
Gc1_22 0 n2 ns22 0 -0.00540660772468
Gc1_23 0 n2 ns23 0 -0.000245273126604
Gc1_24 0 n2 ns24 0 0.00304092260917
Gc1_25 0 n2 ns25 0 -0.000425900367094
Gc1_26 0 n2 ns26 0 -0.000226963061855
Gc1_27 0 n2 ns27 0 0.00159595629012
Gc1_28 0 n2 ns28 0 -0.00673461122134
Gc1_29 0 n2 ns29 0 -0.00789327691041
Gc1_30 0 n2 ns30 0 -0.0128067887866
Gc1_31 0 n2 ns31 0 -0.00145306504782
Gc1_32 0 n2 ns32 0 -0.00196516263974
Gc1_33 0 n2 ns33 0 0.00144545260449
Gc1_34 0 n2 ns34 0 -0.0148455517468
Gc1_35 0 n2 ns35 0 -0.00271620430015
Gc1_36 0 n2 ns36 0 0.00322013550412
Gc1_37 0 n2 ns37 0 9.32850383681e-06
Gc1_38 0 n2 ns38 0 0.0116505548497
Gc1_39 0 n2 ns39 0 -0.000522633064726
Gc1_40 0 n2 ns40 0 -0.00132294932984
Gc1_41 0 n2 ns41 0 -6.14374348827e-06
Gc1_42 0 n2 ns42 0 -6.30832570773e-06
Gc1_43 0 n2 ns43 0 0.000236048250519
Gc1_44 0 n2 ns44 0 -2.18714591071e-05
Gc1_45 0 n2 ns45 0 -0.000448940664989
Gc1_46 0 n2 ns46 0 -1.01766369729e-05
Gc1_47 0 n2 ns47 0 0.000309149910116
Gc1_48 0 n2 ns48 0 -7.59937533176e-05
Gc1_49 0 n2 ns49 0 0.00056817461172
Gc1_50 0 n2 ns50 0 -0.000120727821715
Gc1_51 0 n2 ns51 0 -0.000294973227016
Gc1_52 0 n2 ns52 0 0.000371605917286
Gc1_53 0 n2 ns53 0 8.13308355622e-05
Gc1_54 0 n2 ns54 0 -0.000847474871517
Gc1_55 0 n2 ns55 0 -0.00107558651048
Gc1_56 0 n2 ns56 0 0.000398966734269
Gc1_57 0 n2 ns57 0 -0.000197138930309
Gc1_58 0 n2 ns58 0 0.000881420102543
Gc1_59 0 n2 ns59 0 -0.00249943822312
Gc1_60 0 n2 ns60 0 0.000554126067756
Gc1_61 0 n2 ns61 0 0.00240782011619
Gc1_62 0 n2 ns62 0 -0.000234193818335
Gc1_63 0 n2 ns63 0 -0.000279113463334
Gc1_64 0 n2 ns64 0 0.00177331483978
Gc1_65 0 n2 ns65 0 -0.00278495836661
Gc1_66 0 n2 ns66 0 -0.00190494484905
Gc1_67 0 n2 ns67 0 -0.00766326406645
Gc1_68 0 n2 ns68 0 0.000173062519506
Gc1_69 0 n2 ns69 0 -0.00264086815815
Gc1_70 0 n2 ns70 0 0.00152998383586
Gc1_71 0 n2 ns71 0 -0.0187820376083
Gc1_72 0 n2 ns72 0 -0.00375878490179
Gc1_73 0 n2 ns73 0 0.00686912516919
Gc1_74 0 n2 ns74 0 5.19400911711e-06
Gc1_75 0 n2 ns75 0 0.00217646968611
Gc1_76 0 n2 ns76 0 -0.000914690151819
Gc1_77 0 n2 ns77 0 -0.000452826446091
Gc1_78 0 n2 ns78 0 -1.15241559807e-05
Gc1_79 0 n2 ns79 0 -3.3703214496e-06
Gc1_80 0 n2 ns80 0 0.000193134008985
Gc1_81 0 n2 ns81 0 -9.50392072803e-05
Gc1_82 0 n2 ns82 0 -0.000134244061742
Gc1_83 0 n2 ns83 0 0.000587456746533
Gc1_84 0 n2 ns84 0 -0.000172263728834
Gc1_85 0 n2 ns85 0 0.00046805061971
Gc1_86 0 n2 ns86 0 -0.00207330506334
Gc1_87 0 n2 ns87 0 0.000356072832515
Gc1_88 0 n2 ns88 0 -0.000299620779005
Gc1_89 0 n2 ns89 0 0.00032488215145
Gc1_90 0 n2 ns90 0 -0.000810879502454
Gc1_91 0 n2 ns91 0 0.000686466030814
Gc1_92 0 n2 ns92 0 0.0014375784017
Gc1_93 0 n2 ns93 0 -0.00128096975705
Gc1_94 0 n2 ns94 0 -0.00026856665544
Gc1_95 0 n2 ns95 0 0.000753425763238
Gc1_96 0 n2 ns96 0 0.0035846317741
Gc1_97 0 n2 ns97 0 0.00269292085487
Gc1_98 0 n2 ns98 0 -0.00214069966692
Gc1_99 0 n2 ns99 0 0.0010259092373
Gc1_100 0 n2 ns100 0 -0.000401528397749
Gc1_101 0 n2 ns101 0 0.00141552100929
Gc1_102 0 n2 ns102 0 0.00495880178816
Gc1_103 0 n2 ns103 0 0.00981629834417
Gc1_104 0 n2 ns104 0 0.011179177519
Gc1_105 0 n2 ns105 0 0.00163721909556
Gc1_106 0 n2 ns106 0 -0.0024464837132
Gc1_107 0 n2 ns107 0 0.00182177425986
Gc1_108 0 n2 ns108 0 -0.012312208844
Gc1_109 0 n2 ns109 0 -0.00842663221506
Gc1_110 0 n2 ns110 0 0.0121258713882
Gc1_111 0 n2 ns111 0 1.10240968532e-06
Gc1_112 0 n2 ns112 0 0.00847015168118
Gc1_113 0 n2 ns113 0 -0.000945692155226
Gc1_114 0 n2 ns114 0 -0.000156415016991
Gc1_115 0 n2 ns115 0 -3.03632373508e-05
Gc1_116 0 n2 ns116 0 -1.1932288084e-05
Gc1_117 0 n2 ns117 0 0.00042361062159
Gc1_118 0 n2 ns118 0 -5.74635571025e-05
Gc1_119 0 n2 ns119 0 -0.000386445823665
Gc1_120 0 n2 ns120 0 0.000343565600839
Gc1_121 0 n2 ns121 0 -0.000178826535942
Gc1_122 0 n2 ns122 0 0.000564148283153
Gc1_123 0 n2 ns123 0 -0.00131703294619
Gc1_124 0 n2 ns124 0 -0.000788183498029
Gc1_125 0 n2 ns125 0 -0.000322514422287
Gc1_126 0 n2 ns126 0 0.000401992584575
Gc1_127 0 n2 ns127 0 -4.49266950833e-05
Gc1_128 0 n2 ns128 0 0.000471290777668
Gc1_129 0 n2 ns129 0 0.00129397130655
Gc1_130 0 n2 ns130 0 -0.000235411796042
Gc1_131 0 n2 ns131 0 -0.000219880817969
Gc1_132 0 n2 ns132 0 0.000900548523287
Gc1_133 0 n2 ns133 0 0.0013601923931
Gc1_134 0 n2 ns134 0 0.00103277771807
Gc1_135 0 n2 ns135 0 -0.00184579945016
Gc1_136 0 n2 ns136 0 0.000224234569384
Gc1_137 0 n2 ns137 0 -0.00040786786881
Gc1_138 0 n2 ns138 0 0.00153129149041
Gc1_139 0 n2 ns139 0 0.00387717708835
Gc1_140 0 n2 ns140 0 0.00593218891172
Gc1_141 0 n2 ns141 0 0.0100558491385
Gc1_142 0 n2 ns142 0 0.00164799846318
Gc1_143 0 n2 ns143 0 -0.00301940763953
Gc1_144 0 n2 ns144 0 0.00196009222925
Gc1_145 0 n2 ns145 0 -0.00197886546087
Gc1_146 0 n2 ns146 0 -0.0113338492581
Gc1_147 0 n2 ns147 0 0.00224891796606
Gc1_148 0 n2 ns148 0 4.36079514826e-06
Gc1_149 0 n2 ns149 0 -0.000137579306668
Gc1_150 0 n2 ns150 0 -0.00131688852125
Gc1_151 0 n2 ns151 0 -0.00102576899881
Gc1_152 0 n2 ns152 0 -3.52957991937e-06
Gc1_153 0 n2 ns153 0 -2.05807588648e-05
Gc1_154 0 n2 ns154 0 6.89510108628e-05
Gc1_155 0 n2 ns155 0 0.000261083353747
Gc1_156 0 n2 ns156 0 -0.000570040339822
Gc1_157 0 n2 ns157 0 -0.000212332644995
Gc1_158 0 n2 ns158 0 -0.000160822558169
Gc1_159 0 n2 ns159 0 0.000237007526086
Gc1_160 0 n2 ns160 0 -0.00281942068156
Gc1_161 0 n2 ns161 0 0.000631987780667
Gc1_162 0 n2 ns162 0 0.000255810921592
Gc1_163 0 n2 ns163 0 -0.00032453425551
Gc1_164 0 n2 ns164 0 -0.00075149099453
Gc1_165 0 n2 ns165 0 0.000681891710517
Gc1_166 0 n2 ns166 0 -0.00284915402945
Gc1_167 0 n2 ns167 0 0.00105681769981
Gc1_168 0 n2 ns168 0 -0.000238168216271
Gc1_169 0 n2 ns169 0 0.000809147978602
Gc1_170 0 n2 ns170 0 -0.00459328756148
Gc1_171 0 n2 ns171 0 0.00873010483169
Gc1_172 0 n2 ns172 0 -0.00313547523081
Gc1_173 0 n2 ns173 0 0.000920313719598
Gc1_174 0 n2 ns174 0 0.000188696255121
Gc1_175 0 n2 ns175 0 -0.00156698126586
Gc1_176 0 n2 ns176 0 0.0109925809252
Gc1_177 0 n2 ns177 0 0.0246304680392
Gc1_178 0 n2 ns178 0 -0.00808679815659
Gc1_179 0 n2 ns179 0 0.00937920158165
Gc1_180 0 n2 ns180 0 -0.00212424101495
Gc1_181 0 n2 ns181 0 0.000711642366691
Gc1_182 0 n2 ns182 0 0.0575919941857
Gc1_183 0 n2 ns183 0 -0.00719689701924
Gc1_184 0 n2 ns184 0 -0.0356754948849
Gc1_185 0 n2 ns185 0 2.10961235039e-05
Gc1_186 0 n2 ns186 0 0.00307828984129
Gc1_187 0 n2 ns187 0 -0.000978633064165
Gc1_188 0 n2 ns188 0 0.000686667790227
Gc1_189 0 n2 ns189 0 -2.09924007053e-05
Gc1_190 0 n2 ns190 0 -2.16809901946e-06
Gc1_191 0 n2 ns191 0 0.000435801497816
Gc1_192 0 n2 ns192 0 -0.000143547058374
Gc1_193 0 n2 ns193 0 -0.00064747556274
Gc1_194 0 n2 ns194 0 0.000754299843954
Gc1_195 0 n2 ns195 0 -0.0006837308661
Gc1_196 0 n2 ns196 0 0.000313575462497
Gc1_197 0 n2 ns197 0 0.00135305506405
Gc1_198 0 n2 ns198 0 0.000342380565087
Gc1_199 0 n2 ns199 0 0.000267149396601
Gc1_200 0 n2 ns200 0 -0.000383475567622
Gc1_201 0 n2 ns201 0 0.000445476707242
Gc1_202 0 n2 ns202 0 -0.000996329305835
Gc1_203 0 n2 ns203 0 -0.00072565871553
Gc1_204 0 n2 ns204 0 0.000938988786169
Gc1_205 0 n2 ns205 0 -0.000149479519802
Gc1_206 0 n2 ns206 0 0.00092643667816
Gc1_207 0 n2 ns207 0 0.0112996385347
Gc1_208 0 n2 ns208 0 -0.00591408836196
Gc1_209 0 n2 ns209 0 -0.00186677247397
Gc1_210 0 n2 ns210 0 -0.000109721259747
Gc1_211 0 n2 ns211 0 0.000362921228162
Gc1_212 0 n2 ns212 0 -0.0017118633977
Gc1_213 0 n2 ns213 0 -0.00252591785694
Gc1_214 0 n2 ns214 0 -0.0301118096404
Gc1_215 0 n2 ns215 0 -0.00432126014592
Gc1_216 0 n2 ns216 0 -0.0108536224374
Gc1_217 0 n2 ns217 0 -0.00311158215914
Gc1_218 0 n2 ns218 0 0.00225422806264
Gc1_219 0 n2 ns219 0 -0.0149352911923
Gc1_220 0 n2 ns220 0 0.0127056778017
Gc1_221 0 n2 ns221 0 0.0181232303182
Gc1_222 0 n2 ns222 0 -1.22184931046e-05
Gc1_223 0 n2 ns223 0 -0.00219636688213
Gc1_224 0 n2 ns224 0 0.000886758447146
Gc1_225 0 n2 ns225 0 1.08742803413e-05
Gc1_226 0 n2 ns226 0 2.08387025353e-05
Gc1_227 0 n2 ns227 0 2.39386821189e-05
Gc1_228 0 n2 ns228 0 -0.000170759887379
Gc1_229 0 n2 ns229 0 -0.000156196908494
Gc1_230 0 n2 ns230 0 -3.56763554456e-06
Gc1_231 0 n2 ns231 0 -0.000122465960937
Gc1_232 0 n2 ns232 0 0.000508298306901
Gc1_233 0 n2 ns233 0 -0.000402918273733
Gc1_234 0 n2 ns234 0 0.00096153848505
Gc1_235 0 n2 ns235 0 -0.000648406294999
Gc1_236 0 n2 ns236 0 0.000322566050447
Gc1_237 0 n2 ns237 0 -0.000316233934587
Gc1_238 0 n2 ns238 0 0.000900819500557
Gc1_239 0 n2 ns239 0 0.00105568812387
Gc1_240 0 n2 ns240 0 0.00237159810378
Gc1_241 0 n2 ns241 0 -0.000915009072509
Gc1_242 0 n2 ns242 0 -0.000175080526351
Gc1_243 0 n2 ns243 0 0.000700317446172
Gc1_244 0 n2 ns244 0 -0.00619986619197
Gc1_245 0 n2 ns245 0 0.000345448937945
Gc1_246 0 n2 ns246 0 0.00273647142708
Gc1_247 0 n2 ns247 0 -0.000677324696456
Gc1_248 0 n2 ns248 0 0.000427347193269
Gc1_249 0 n2 ns249 0 -0.00126808616227
Gc1_250 0 n2 ns250 0 -0.0026271807494
Gc1_251 0 n2 ns251 0 0.0103353077776
Gc1_252 0 n2 ns252 0 0.00765272001825
Gc1_253 0 n2 ns253 0 0.00328242433718
Gc1_254 0 n2 ns254 0 -0.00215360501472
Gc1_255 0 n2 ns255 0 0.00175095929366
Gc1_256 0 n2 ns256 0 0.00225573823005
Gc1_257 0 n2 ns257 0 0.00875848202247
Gc1_258 0 n2 ns258 0 -0.00327727788168
Gc1_259 0 n2 ns259 0 -4.89663825961e-06
Gc1_260 0 n2 ns260 0 0.000930893746659
Gc1_261 0 n2 ns261 0 0.000390272179202
Gc1_262 0 n2 ns262 0 0.000346896718907
Gc1_263 0 n2 ns263 0 1.0583588573e-05
Gc1_264 0 n2 ns264 0 1.21332859692e-05
Gc1_265 0 n2 ns265 0 1.80528931606e-05
Gc1_266 0 n2 ns266 0 -0.000211783086318
Gc1_267 0 n2 ns267 0 7.44025815848e-05
Gc1_268 0 n2 ns268 0 0.000241499088942
Gc1_269 0 n2 ns269 0 0.000305806801438
Gc1_270 0 n2 ns270 0 -0.00018641089189
Gc1_271 0 n2 ns271 0 0.00135886257962
Gc1_272 0 n2 ns272 0 -0.000512160288199
Gc1_273 0 n2 ns273 0 0.000324970833482
Gc1_274 0 n2 ns274 0 -0.000372851039728
Gc1_275 0 n2 ns275 0 0.000388750962136
Gc1_276 0 n2 ns276 0 0.000799795663274
Gc1_277 0 n2 ns277 0 0.00173043508161
Gc1_278 0 n2 ns278 0 -0.000183480388234
Gc1_279 0 n2 ns279 0 -0.00017276650256
Gc1_280 0 n2 ns280 0 0.000871929272792
Gc1_281 0 n2 ns281 0 -0.0020444394013
Gc1_282 0 n2 ns282 0 -0.00315159750284
Gc1_283 0 n2 ns283 0 0.00172590810416
Gc1_284 0 n2 ns284 0 -0.000523118108892
Gc1_285 0 n2 ns285 0 0.000458699653148
Gc1_286 0 n2 ns286 0 -0.00156143591291
Gc1_287 0 n2 ns287 0 -0.0030162221473
Gc1_288 0 n2 ns288 0 -0.000192384369104
Gc1_289 0 n2 ns289 0 0.00555290996903
Gc1_290 0 n2 ns290 0 -0.000854843646492
Gc1_291 0 n2 ns291 0 -0.00269912151936
Gc1_292 0 n2 ns292 0 0.00219540696782
Gc1_293 0 n2 ns293 0 0.00230353527392
Gc1_294 0 n2 ns294 0 0.0109005213505
Gc1_295 0 n2 ns295 0 -0.00210730246039
Gc1_296 0 n2 ns296 0 -5.65751252177e-06
Gd1_1 0 n2 ni1 0 -0.00278231931624
Gd1_2 0 n2 ni2 0 -0.00254088312022
Gd1_3 0 n2 ni3 0 -0.000857933704477
Gd1_4 0 n2 ni4 0 -0.00378329763468
Gd1_5 0 n2 ni5 0 0.000552791705623
Gd1_6 0 n2 ni6 0 -0.000405899256147
Gd1_7 0 n2 ni7 0 0.000546119776655
Gd1_8 0 n2 ni8 0 -0.000549183165396
Gc2_1 0 n4 ns1 0 0.0116505548413
Gc2_2 0 n4 ns2 0 -0.000522633063315
Gc2_3 0 n4 ns3 0 -0.0013229493301
Gc2_4 0 n4 ns4 0 -6.14374340974e-06
Gc2_5 0 n4 ns5 0 -6.30832564827e-06
Gc2_6 0 n4 ns6 0 0.000236048250203
Gc2_7 0 n4 ns7 0 -2.18714589773e-05
Gc2_8 0 n4 ns8 0 -0.000448940664824
Gc2_9 0 n4 ns9 0 -1.01766367282e-05
Gc2_10 0 n4 ns10 0 0.000309149910638
Gc2_11 0 n4 ns11 0 -7.59937536346e-05
Gc2_12 0 n4 ns12 0 0.000568174610831
Gc2_13 0 n4 ns13 0 -0.000120727820252
Gc2_14 0 n4 ns14 0 -0.000294973226978
Gc2_15 0 n4 ns15 0 0.000371605917198
Gc2_16 0 n4 ns16 0 8.13308337935e-05
Gc2_17 0 n4 ns17 0 -0.000847474874555
Gc2_18 0 n4 ns18 0 -0.0010755865125
Gc2_19 0 n4 ns19 0 0.000398966731939
Gc2_20 0 n4 ns20 0 -0.000197138930717
Gc2_21 0 n4 ns21 0 0.000881420102826
Gc2_22 0 n4 ns22 0 -0.00249943821556
Gc2_23 0 n4 ns23 0 0.000554126071664
Gc2_24 0 n4 ns24 0 0.00240782011584
Gc2_25 0 n4 ns25 0 -0.000234193820648
Gc2_26 0 n4 ns26 0 -0.000279113463049
Gc2_27 0 n4 ns27 0 0.00177331483912
Gc2_28 0 n4 ns28 0 -0.00278495835038
Gc2_29 0 n4 ns29 0 -0.00190494486789
Gc2_30 0 n4 ns30 0 -0.00766326406276
Gc2_31 0 n4 ns31 0 0.000173062499672
Gc2_32 0 n4 ns32 0 -0.00264086815935
Gc2_33 0 n4 ns33 0 0.00152998383875
Gc2_34 0 n4 ns34 0 -0.0187820375794
Gc2_35 0 n4 ns35 0 -0.00375878490639
Gc2_36 0 n4 ns36 0 0.00686912514473
Gc2_37 0 n4 ns37 0 5.19400954392e-06
Gc2_38 0 n4 ns38 0 0.00625054372057
Gc2_39 0 n4 ns39 0 0.0005431399143
Gc2_40 0 n4 ns40 0 -0.00124822165685
Gc2_41 0 n4 ns41 0 1.66958832304e-05
Gc2_42 0 n4 ns42 0 5.34202429075e-06
Gc2_43 0 n4 ns43 0 9.55740333542e-05
Gc2_44 0 n4 ns44 0 1.78360396165e-05
Gc2_45 0 n4 ns45 0 -0.000313837406935
Gc2_46 0 n4 ns46 0 0.000125305287262
Gc2_47 0 n4 ns47 0 0.000323499446097
Gc2_48 0 n4 ns48 0 -0.000161768544805
Gc2_49 0 n4 ns49 0 0.000153846819142
Gc2_50 0 n4 ns50 0 0.000522403255015
Gc2_51 0 n4 ns51 0 -0.000383794250368
Gc2_52 0 n4 ns52 0 0.000444263585014
Gc2_53 0 n4 ns53 0 -0.000157323008477
Gc2_54 0 n4 ns54 0 -0.000915072575424
Gc2_55 0 n4 ns55 0 -0.000813931369428
Gc2_56 0 n4 ns56 0 7.39706481955e-05
Gc2_57 0 n4 ns57 0 -0.000260456810427
Gc2_58 0 n4 ns58 0 0.0010464459367
Gc2_59 0 n4 ns59 0 -0.00259005008495
Gc2_60 0 n4 ns60 0 0.00103617172229
Gc2_61 0 n4 ns61 0 0.00171121112377
Gc2_62 0 n4 ns62 0 -9.35122890862e-05
Gc2_63 0 n4 ns63 0 -0.000393367680972
Gc2_64 0 n4 ns64 0 0.00196908694669
Gc2_65 0 n4 ns65 0 -0.00339287155517
Gc2_66 0 n4 ns66 0 -0.00349699118912
Gc2_67 0 n4 ns67 0 -0.00593479963724
Gc2_68 0 n4 ns68 0 -0.00089395120201
Gc2_69 0 n4 ns69 0 -0.00304780449005
Gc2_70 0 n4 ns70 0 0.00198668432661
Gc2_71 0 n4 ns71 0 -0.0145165924003
Gc2_72 0 n4 ns72 0 -0.00759268208289
Gc2_73 0 n4 ns73 0 0.00475786764574
Gc2_74 0 n4 ns74 0 1.04565049628e-05
Gc2_75 0 n4 ns75 0 0.00847331945783
Gc2_76 0 n4 ns76 0 -0.00093677920452
Gc2_77 0 n4 ns77 0 -0.00014925399047
Gc2_78 0 n4 ns78 0 -3.06939171396e-05
Gc2_79 0 n4 ns79 0 -1.19125203008e-05
Gc2_80 0 n4 ns80 0 0.000422538681942
Gc2_81 0 n4 ns81 0 -5.53225034253e-05
Gc2_82 0 n4 ns82 0 -0.000385684879645
Gc2_83 0 n4 ns83 0 0.000344359883332
Gc2_84 0 n4 ns84 0 -0.000176749415023
Gc2_85 0 n4 ns85 0 0.000562041457149
Gc2_86 0 n4 ns86 0 -0.00131350354435
Gc2_87 0 n4 ns87 0 -0.000796219243683
Gc2_88 0 n4 ns88 0 -0.000321382490749
Gc2_89 0 n4 ns89 0 0.000399781676424
Gc2_90 0 n4 ns90 0 -3.4021313659e-05
Gc2_91 0 n4 ns91 0 0.000463830099842
Gc2_92 0 n4 ns92 0 0.00129488559407
Gc2_93 0 n4 ns93 0 -0.000231779433246
Gc2_94 0 n4 ns94 0 -0.000219913038315
Gc2_95 0 n4 ns95 0 0.000897289563627
Gc2_96 0 n4 ns96 0 0.0013345225053
Gc2_97 0 n4 ns97 0 0.00102674028509
Gc2_98 0 n4 ns98 0 -0.00184799584112
Gc2_99 0 n4 ns99 0 0.000214243237835
Gc2_100 0 n4 ns100 0 -0.000410977314922
Gc2_101 0 n4 ns101 0 0.00152420556576
Gc2_102 0 n4 ns102 0 0.00384645749683
Gc2_103 0 n4 ns103 0 0.00587962269951
Gc2_104 0 n4 ns104 0 0.0100318830063
Gc2_105 0 n4 ns105 0 0.00164305854602
Gc2_106 0 n4 ns106 0 -0.00301798403914
Gc2_107 0 n4 ns107 0 0.00195452607041
Gc2_108 0 n4 ns108 0 -0.00185968777111
Gc2_109 0 n4 ns109 0 -0.0113527306012
Gc2_110 0 n4 ns110 0 0.00214933508651
Gc2_111 0 n4 ns111 0 4.3313987259e-06
Gc2_112 0 n4 ns112 0 0.00771492429977
Gc2_113 0 n4 ns113 0 -0.000608905294568
Gc2_114 0 n4 ns114 0 -0.000864652452881
Gc2_115 0 n4 ns115 0 -1.01158258342e-05
Gc2_116 0 n4 ns116 0 3.65373165151e-06
Gc2_117 0 n4 ns117 0 0.000334455175408
Gc2_118 0 n4 ns118 0 -7.0471818245e-05
Gc2_119 0 n4 ns119 0 -0.000327246029187
Gc2_120 0 n4 ns120 0 0.000416007120892
Gc2_121 0 n4 ns121 0 2.65089270702e-05
Gc2_122 0 n4 ns122 0 0.00027123273367
Gc2_123 0 n4 ns123 0 -0.00141125401102
Gc2_124 0 n4 ns124 0 2.27509306634e-05
Gc2_125 0 n4 ns125 0 -0.000382300506097
Gc2_126 0 n4 ns126 0 0.000444698959007
Gc2_127 0 n4 ns127 0 -0.000633141981862
Gc2_128 0 n4 ns128 0 -0.000107751946929
Gc2_129 0 n4 ns129 0 0.000703741795663
Gc2_130 0 n4 ns130 0 -0.000623052706137
Gc2_131 0 n4 ns131 0 -0.00031638797516
Gc2_132 0 n4 ns132 0 0.0010098994879
Gc2_133 0 n4 ns133 0 0.00104129553592
Gc2_134 0 n4 ns134 0 0.00234078420582
Gc2_135 0 n4 ns135 0 -0.000665229270145
Gc2_136 0 n4 ns136 0 0.000588408683983
Gc2_137 0 n4 ns137 0 -0.000535854142929
Gc2_138 0 n4 ns138 0 0.00193830648253
Gc2_139 0 n4 ns139 0 0.00278560191768
Gc2_140 0 n4 ns140 0 0.00555805763819
Gc2_141 0 n4 ns141 0 0.0054275930499
Gc2_142 0 n4 ns142 0 0.000520679228271
Gc2_143 0 n4 ns143 0 -0.00332866421578
Gc2_144 0 n4 ns144 0 0.00226496111304
Gc2_145 0 n4 ns145 0 -0.0136298509568
Gc2_146 0 n4 ns146 0 -0.00887386569867
Gc2_147 0 n4 ns147 0 0.00845547478319
Gc2_148 0 n4 ns148 0 3.66622502579e-06
Gc2_149 0 n4 ns149 0 0.00308942158893
Gc2_150 0 n4 ns150 0 -0.000982873366334
Gc2_151 0 n4 ns151 0 0.000689655568728
Gc2_152 0 n4 ns152 0 -2.13649950085e-05
Gc2_153 0 n4 ns153 0 -2.27333834822e-06
Gc2_154 0 n4 ns154 0 0.000436598930722
Gc2_155 0 n4 ns155 0 -0.00014237874172
Gc2_156 0 n4 ns156 0 -0.000646471536482
Gc2_157 0 n4 ns157 0 0.000755857007223
Gc2_158 0 n4 ns158 0 -0.000684144397633
Gc2_159 0 n4 ns159 0 0.000312916595143
Gc2_160 0 n4 ns160 0 0.00135321634677
Gc2_161 0 n4 ns161 0 0.000339576727642
Gc2_162 0 n4 ns162 0 0.000267441961464
Gc2_163 0 n4 ns163 0 -0.00038432006448
Gc2_164 0 n4 ns164 0 0.000449625704937
Gc2_165 0 n4 ns165 0 -0.000994870024813
Gc2_166 0 n4 ns166 0 -0.000723634521999
Gc2_167 0 n4 ns167 0 0.000937539568817
Gc2_168 0 n4 ns168 0 -0.000149037250512
Gc2_169 0 n4 ns169 0 0.000926859358588
Gc2_170 0 n4 ns170 0 0.0113005431745
Gc2_171 0 n4 ns171 0 -0.00591516905293
Gc2_172 0 n4 ns172 0 -0.00186948737682
Gc2_173 0 n4 ns173 0 -0.000109109469853
Gc2_174 0 n4 ns174 0 0.000361779953751
Gc2_175 0 n4 ns175 0 -0.00171196992656
Gc2_176 0 n4 ns176 0 -0.00252873385471
Gc2_177 0 n4 ns177 0 -0.0301088556674
Gc2_178 0 n4 ns178 0 -0.0043223351472
Gc2_179 0 n4 ns179 0 -0.010850272905
Gc2_180 0 n4 ns180 0 -0.00311111761003
Gc2_181 0 n4 ns181 0 0.00225380850348
Gc2_182 0 n4 ns182 0 -0.0150095753092
Gc2_183 0 n4 ns183 0 0.0126980662811
Gc2_184 0 n4 ns184 0 0.0181943532783
Gc2_185 0 n4 ns185 0 -1.23297933126e-05
Gc2_186 0 n4 ns186 0 -0.00032880076285
Gc2_187 0 n4 ns187 0 -5.05393171709e-05
Gc2_188 0 n4 ns188 0 -0.00104537507027
Gc2_189 0 n4 ns189 0 1.56091714114e-05
Gc2_190 0 n4 ns190 0 -1.21897220495e-06
Gc2_191 0 n4 ns191 0 3.06285681893e-05
Gc2_192 0 n4 ns192 0 0.000168642063364
Gc2_193 0 n4 ns193 0 -0.000162058425083
Gc2_194 0 n4 ns194 0 -0.000246470266581
Gc2_195 0 n4 ns195 0 0.000321736717792
Gc2_196 0 n4 ns196 0 -0.000176097839869
Gc2_197 0 n4 ns197 0 -0.00237938449303
Gc2_198 0 n4 ns198 0 0.000207305799182
Gc2_199 0 n4 ns199 0 0.000379690341758
Gc2_200 0 n4 ns200 0 -0.000480273718659
Gc2_201 0 n4 ns201 0 -0.000625153519831
Gc2_202 0 n4 ns202 0 0.00119403781396
Gc2_203 0 n4 ns203 0 -0.00171497652687
Gc2_204 0 n4 ns204 0 0.000207316666904
Gc2_205 0 n4 ns205 0 -0.000314316857991
Gc2_206 0 n4 ns206 0 0.00106355475875
Gc2_207 0 n4 ns207 0 -0.00857417663023
Gc2_208 0 n4 ns208 0 0.00821160625606
Gc2_209 0 n4 ns209 0 -0.00185942135432
Gc2_210 0 n4 ns210 0 0.000269882730209
Gc2_211 0 n4 ns211 0 0.000426762337341
Gc2_212 0 n4 ns212 0 -0.00198927506289
Gc2_213 0 n4 ns213 0 0.00880745864912
Gc2_214 0 n4 ns214 0 0.0288486658198
Gc2_215 0 n4 ns215 0 -0.00495336044776
Gc2_216 0 n4 ns216 0 0.00996243973267
Gc2_217 0 n4 ns217 0 -0.00288268758713
Gc2_218 0 n4 ns218 0 0.00128771200617
Gc2_219 0 n4 ns219 0 0.0606554498573
Gc2_220 0 n4 ns220 0 -0.00372057863517
Gc2_221 0 n4 ns221 0 -0.0393302563852
Gc2_222 0 n4 ns222 0 1.74002039589e-05
Gc2_223 0 n4 ns223 0 0.000899858151181
Gc2_224 0 n4 ns224 0 0.000384024672199
Gc2_225 0 n4 ns225 0 0.000348907039136
Gc2_226 0 n4 ns226 0 1.0574732298e-05
Gc2_227 0 n4 ns227 0 1.19296060708e-05
Gc2_228 0 n4 ns228 0 1.55695231305e-05
Gc2_229 0 n4 ns229 0 -0.000211320393897
Gc2_230 0 n4 ns230 0 7.58481522066e-05
Gc2_231 0 n4 ns231 0 0.000240381090282
Gc2_232 0 n4 ns232 0 0.000301315896535
Gc2_233 0 n4 ns233 0 -0.000185065256295
Gc2_234 0 n4 ns234 0 0.00135994501661
Gc2_235 0 n4 ns235 0 -0.000506797567599
Gc2_236 0 n4 ns236 0 0.000324046314996
Gc2_237 0 n4 ns237 0 -0.000369211828775
Gc2_238 0 n4 ns238 0 0.000381180280116
Gc2_239 0 n4 ns239 0 0.000797227025684
Gc2_240 0 n4 ns240 0 0.00172319104998
Gc2_241 0 n4 ns241 0 -0.000170912607698
Gc2_242 0 n4 ns242 0 -0.000173175545461
Gc2_243 0 n4 ns243 0 0.000867915337869
Gc2_244 0 n4 ns244 0 -0.00204894058134
Gc2_245 0 n4 ns245 0 -0.00316342923793
Gc2_246 0 n4 ns246 0 0.00172826299708
Gc2_247 0 n4 ns247 0 -0.000510009953924
Gc2_248 0 n4 ns248 0 0.000461669286731
Gc2_249 0 n4 ns249 0 -0.00155431399938
Gc2_250 0 n4 ns250 0 -0.00302899074664
Gc2_251 0 n4 ns251 0 -0.000174317133803
Gc2_252 0 n4 ns252 0 0.00555405350411
Gc2_253 0 n4 ns253 0 -0.000825870682892
Gc2_254 0 n4 ns254 0 -0.00270145374595
Gc2_255 0 n4 ns255 0 0.0021851494235
Gc2_256 0 n4 ns256 0 0.00238937492845
Gc2_257 0 n4 ns257 0 0.0109090947593
Gc2_258 0 n4 ns258 0 -0.00219023752386
Gc2_259 0 n4 ns259 0 -5.57496340916e-06
Gc2_260 0 n4 ns260 0 0.00160303134279
Gc2_261 0 n4 ns261 0 -8.87190071409e-05
Gc2_262 0 n4 ns262 0 0.000446673532483
Gc2_263 0 n4 ns263 0 -5.93886449069e-06
Gc2_264 0 n4 ns264 0 1.17695465201e-05
Gc2_265 0 n4 ns265 0 0.000268865141772
Gc2_266 0 n4 ns266 0 -0.00018910838287
Gc2_267 0 n4 ns267 0 -0.000511741880332
Gc2_268 0 n4 ns268 0 0.000301172814192
Gc2_269 0 n4 ns269 0 -1.21231108023e-05
Gc2_270 0 n4 ns270 0 -1.26900857737e-05
Gc2_271 0 n4 ns271 0 0.00136663339326
Gc2_272 0 n4 ns272 0 -0.000158071984263
Gc2_273 0 n4 ns273 0 0.000395288144106
Gc2_274 0 n4 ns274 0 -0.000447288815685
Gc2_275 0 n4 ns275 0 0.000949426519006
Gc2_276 0 n4 ns276 0 0.000806267452461
Gc2_277 0 n4 ns277 0 0.00143593245474
Gc2_278 0 n4 ns278 0 0.000424966831518
Gc2_279 0 n4 ns279 0 -0.000188100668422
Gc2_280 0 n4 ns280 0 0.00103719865474
Gc2_281 0 n4 ns281 0 0.00106781725372
Gc2_282 0 n4 ns282 0 -0.00329561839411
Gc2_283 0 n4 ns283 0 0.00106161984305
Gc2_284 0 n4 ns284 0 -0.000322928444737
Gc2_285 0 n4 ns285 0 0.000516438761738
Gc2_286 0 n4 ns286 0 -0.0018468414149
Gc2_287 0 n4 ns287 0 -0.00157129103196
Gc2_288 0 n4 ns288 0 -0.00704567112977
Gc2_289 0 n4 ns289 0 0.00450243552422
Gc2_290 0 n4 ns290 0 -0.0032208423854
Gc2_291 0 n4 ns291 0 -0.00327010797433
Gc2_292 0 n4 ns292 0 0.00253284165661
Gc2_293 0 n4 ns293 0 0.00164444276588
Gc2_294 0 n4 ns294 0 0.0128961983263
Gc2_295 0 n4 ns295 0 -0.000325435476627
Gc2_296 0 n4 ns296 0 -6.31233974844e-06
Gd2_1 0 n4 ni1 0 -0.00254088311604
Gd2_2 0 n4 ni2 0 -0.000206815792148
Gd2_3 0 n4 ni3 0 -0.00379334480167
Gd2_4 0 n4 ni4 0 -0.00241578476693
Gd2_5 0 n4 ni5 0 -0.000408981188342
Gd2_6 0 n4 ni6 0 -4.81368855684e-06
Gd2_7 0 n4 ni7 0 -0.000535648896981
Gd2_8 0 n4 ni8 0 -0.000366569186702
Gc3_1 0 n6 ns1 0 0.0021764697717
Gc3_2 0 n6 ns2 0 -0.000914690220157
Gc3_3 0 n6 ns3 0 -0.000452826466697
Gc3_4 0 n6 ns4 0 -1.15241562897e-05
Gc3_5 0 n6 ns5 0 -3.37032167754e-06
Gc3_6 0 n6 ns6 0 0.000193134011334
Gc3_7 0 n6 ns7 0 -9.50392088361e-05
Gc3_8 0 n6 ns8 0 -0.000134244060173
Gc3_9 0 n6 ns9 0 0.000587456744427
Gc3_10 0 n6 ns10 0 -0.000172263727756
Gc3_11 0 n6 ns11 0 0.000468050616305
Gc3_12 0 n6 ns12 0 -0.00207330505805
Gc3_13 0 n6 ns13 0 0.000356072848607
Gc3_14 0 n6 ns14 0 -0.000299620780766
Gc3_15 0 n6 ns15 0 0.00032488215024
Gc3_16 0 n6 ns16 0 -0.000810879536633
Gc3_17 0 n6 ns17 0 0.000686466032223
Gc3_18 0 n6 ns18 0 0.00143757838068
Gc3_19 0 n6 ns19 0 -0.0012809697627
Gc3_20 0 n6 ns20 0 -0.000268566658431
Gc3_21 0 n6 ns21 0 0.000753425763541
Gc3_22 0 n6 ns22 0 0.00358463192868
Gc3_23 0 n6 ns23 0 0.00269292094594
Gc3_24 0 n6 ns24 0 -0.00214069964629
Gc3_25 0 n6 ns25 0 0.00102590918972
Gc3_26 0 n6 ns26 0 -0.000401528383955
Gc3_27 0 n6 ns27 0 0.00141552100753
Gc3_28 0 n6 ns28 0 0.00495880235107
Gc3_29 0 n6 ns29 0 0.00981629835124
Gc3_30 0 n6 ns30 0 0.0111791778597
Gc3_31 0 n6 ns31 0 0.00163721890324
Gc3_32 0 n6 ns32 0 -0.00244648375392
Gc3_33 0 n6 ns33 0 0.00182177428084
Gc3_34 0 n6 ns34 0 -0.0123122075992
Gc3_35 0 n6 ns35 0 -0.0084266323155
Gc3_36 0 n6 ns36 0 0.0121258702435
Gc3_37 0 n6 ns37 0 1.10240867633e-06
Gc3_38 0 n6 ns38 0 0.00847331943228
Gc3_39 0 n6 ns39 0 -0.000936779209847
Gc3_40 0 n6 ns40 0 -0.000149253997209
Gc3_41 0 n6 ns41 0 -3.06939169754e-05
Gc3_42 0 n6 ns42 0 -1.19125202512e-05
Gc3_43 0 n6 ns43 0 0.000422538680229
Gc3_44 0 n6 ns44 0 -5.53225034405e-05
Gc3_45 0 n6 ns45 0 -0.000385684879751
Gc3_46 0 n6 ns46 0 0.000344359882959
Gc3_47 0 n6 ns47 0 -0.000176749415046
Gc3_48 0 n6 ns48 0 0.000562041455709
Gc3_49 0 n6 ns49 0 -0.00131350354323
Gc3_50 0 n6 ns50 0 -0.00079621924059
Gc3_51 0 n6 ns51 0 -0.000321382490486
Gc3_52 0 n6 ns52 0 0.000399781676591
Gc3_53 0 n6 ns53 0 -3.40213161019e-05
Gc3_54 0 n6 ns54 0 0.0004638300908
Gc3_55 0 n6 ns55 0 0.00129488559011
Gc3_56 0 n6 ns56 0 -0.000231779440647
Gc3_57 0 n6 ns57 0 -0.000219913039272
Gc3_58 0 n6 ns58 0 0.000897289564352
Gc3_59 0 n6 ns59 0 0.00133452250578
Gc3_60 0 n6 ns60 0 0.00102674030799
Gc3_61 0 n6 ns61 0 -0.0018479958367
Gc3_62 0 n6 ns62 0 0.000214243242791
Gc3_63 0 n6 ns63 0 -0.000410977315104
Gc3_64 0 n6 ns64 0 0.00152420556776
Gc3_65 0 n6 ns65 0 0.00384645746244
Gc3_66 0 n6 ns66 0 0.00587962282612
Gc3_67 0 n6 ns67 0 0.0100318830304
Gc3_68 0 n6 ns68 0 0.00164305862318
Gc3_69 0 n6 ns69 0 -0.00301798404943
Gc3_70 0 n6 ns70 0 0.00195452606329
Gc3_71 0 n6 ns71 0 -0.0018596882424
Gc3_72 0 n6 ns72 0 -0.0113527305715
Gc3_73 0 n6 ns73 0 0.00214933551585
Gc3_74 0 n6 ns74 0 4.33139917048e-06
Gc3_75 0 n6 ns75 0 0.01054503254
Gc3_76 0 n6 ns76 0 0.000728151524075
Gc3_77 0 n6 ns77 0 -0.00106628816248
Gc3_78 0 n6 ns78 0 2.43023929877e-06
Gc3_79 0 n6 ns79 0 6.10622961635e-06
Gc3_80 0 n6 ns80 0 0.000105651663365
Gc3_81 0 n6 ns81 0 3.00510467748e-05
Gc3_82 0 n6 ns82 0 -0.000410516207985
Gc3_83 0 n6 ns83 0 1.66441295249e-06
Gc3_84 0 n6 ns84 0 0.000533982829396
Gc3_85 0 n6 ns85 0 -0.000220309806234
Gc3_86 0 n6 ns86 0 0.000806327875658
Gc3_87 0 n6 ns87 0 -0.000282880320079
Gc3_88 0 n6 ns88 0 -0.00020365678918
Gc3_89 0 n6 ns89 0 0.000281565756996
Gc3_90 0 n6 ns90 0 0.000655491327606
Gc3_91 0 n6 ns91 0 -0.00148037901952
Gc3_92 0 n6 ns92 0 -0.0012665381565
Gc3_93 0 n6 ns93 0 0.000762620481537
Gc3_94 0 n6 ns94 0 -0.000142839815924
Gc3_95 0 n6 ns95 0 0.000704291082155
Gc3_96 0 n6 ns96 0 -0.00543284866473
Gc3_97 0 n6 ns97 0 -0.000295588096127
Gc3_98 0 n6 ns98 0 0.00304461694913
Gc3_99 0 n6 ns99 0 -0.00040569857881
Gc3_100 0 n6 ns100 0 -0.000235795556932
Gc3_101 0 n6 ns101 0 0.00158615746609
Gc3_102 0 n6 ns102 0 -0.00679801311559
Gc3_103 0 n6 ns103 0 -0.00804628452419
Gc3_104 0 n6 ns104 0 -0.0129129861926
Gc3_105 0 n6 ns105 0 -0.00154217230081
Gc3_106 0 n6 ns106 0 -0.00195885883245
Gc3_107 0 n6 ns107 0 0.00143684118009
Gc3_108 0 n6 ns108 0 -0.0147630592298
Gc3_109 0 n6 ns109 0 -0.00273195320372
Gc3_110 0 n6 ns110 0 0.00312966725115
Gc3_111 0 n6 ns111 0 9.51079468889e-06
Gc3_112 0 n6 ns112 0 0.0115985199936
Gc3_113 0 n6 ns113 0 -0.000514465093991
Gc3_114 0 n6 ns114 0 -0.00131513268045
Gc3_115 0 n6 ns115 0 -6.23289115284e-06
Gc3_116 0 n6 ns116 0 -6.33377265491e-06
Gc3_117 0 n6 ns117 0 0.000231626051009
Gc3_118 0 n6 ns118 0 -2.11134902687e-05
Gc3_119 0 n6 ns119 0 -0.000447847874328
Gc3_120 0 n6 ns120 0 -1.35109314013e-05
Gc3_121 0 n6 ns121 0 0.000307496720853
Gc3_122 0 n6 ns122 0 -7.77665241981e-05
Gc3_123 0 n6 ns123 0 0.000579620662486
Gc3_124 0 n6 ns124 0 -0.000128627230996
Gc3_125 0 n6 ns125 0 -0.000293271768096
Gc3_126 0 n6 ns126 0 0.000368772263399
Gc3_127 0 n6 ns127 0 9.63062697939e-05
Gc3_128 0 n6 ns128 0 -0.000851324418094
Gc3_129 0 n6 ns129 0 -0.00107558359444
Gc3_130 0 n6 ns130 0 0.000404443949942
Gc3_131 0 n6 ns131 0 -0.000196794191236
Gc3_132 0 n6 ns132 0 0.000876499288758
Gc3_133 0 n6 ns133 0 -0.00254383660475
Gc3_134 0 n6 ns134 0 0.000534949851881
Gc3_135 0 n6 ns135 0 0.0024092631166
Gc3_136 0 n6 ns136 0 -0.000237180973478
Gc3_137 0 n6 ns137 0 -0.00028388419867
Gc3_138 0 n6 ns138 0 0.00176471410236
Gc3_139 0 n6 ns139 0 -0.00286923727363
Gc3_140 0 n6 ns140 0 -0.00193752544796
Gc3_141 0 n6 ns141 0 -0.00771429834162
Gc3_142 0 n6 ns142 0 0.000202174495553
Gc3_143 0 n6 ns143 0 -0.00263727411913
Gc3_144 0 n6 ns144 0 0.00151510832881
Gc3_145 0 n6 ns145 0 -0.0187877349184
Gc3_146 0 n6 ns146 0 -0.00375997488174
Gc3_147 0 n6 ns147 0 0.00688057677642
Gc3_148 0 n6 ns148 0 5.2966239271e-06
Gc3_149 0 n6 ns149 0 -0.00221425834306
Gc3_150 0 n6 ns150 0 0.000905823012605
Gc3_151 0 n6 ns151 0 2.36904855797e-05
Gc3_152 0 n6 ns152 0 2.10359803631e-05
Gc3_153 0 n6 ns153 0 2.41612054159e-05
Gc3_154 0 n6 ns154 0 -0.000170990085873
Gc3_155 0 n6 ns155 0 -0.000155897853756
Gc3_156 0 n6 ns156 0 -6.5026371559e-06
Gc3_157 0 n6 ns157 0 -0.00012324463491
Gc3_158 0 n6 ns158 0 0.000506095175752
Gc3_159 0 n6 ns159 0 -0.000397134146507
Gc3_160 0 n6 ns160 0 0.000955078376965
Gc3_161 0 n6 ns161 0 -0.000661855466639
Gc3_162 0 n6 ns162 0 0.000323339363122
Gc3_163 0 n6 ns163 0 -0.000315534548186
Gc3_164 0 n6 ns164 0 0.000915990995669
Gc3_165 0 n6 ns165 0 0.00104757028767
Gc3_166 0 n6 ns166 0 0.00237914188625
Gc3_167 0 n6 ns167 0 -0.000917138952935
Gc3_168 0 n6 ns168 0 -0.000174579824859
Gc3_169 0 n6 ns169 0 0.000698517131638
Gc3_170 0 n6 ns170 0 -0.0062373839875
Gc3_171 0 n6 ns171 0 0.000335356754203
Gc3_172 0 n6 ns172 0 0.00273381559841
Gc3_173 0 n6 ns173 0 -0.000668702641802
Gc3_174 0 n6 ns174 0 0.000425221835187
Gc3_175 0 n6 ns175 0 -0.00126604052938
Gc3_176 0 n6 ns176 0 -0.00268355735558
Gc3_177 0 n6 ns177 0 0.0102837123663
Gc3_178 0 n6 ns178 0 0.00761074589181
Gc3_179 0 n6 ns179 0 0.00327320888927
Gc3_180 0 n6 ns180 0 -0.00214889089131
Gc3_181 0 n6 ns181 0 0.00174988889182
Gc3_182 0 n6 ns182 0 0.00230678325067
Gc3_183 0 n6 ns183 0 0.00874268305489
Gc3_184 0 n6 ns184 0 -0.00331689445735
Gc3_185 0 n6 ns185 0 -4.86389707058e-06
Gc3_186 0 n6 ns186 0 0.000905682078281
Gc3_187 0 n6 ns187 0 0.000379093839319
Gc3_188 0 n6 ns188 0 0.000343390700281
Gc3_189 0 n6 ns189 0 1.05182793328e-05
Gc3_190 0 n6 ns190 0 1.19235006255e-05
Gc3_191 0 n6 ns191 0 1.58275209972e-05
Gc3_192 0 n6 ns192 0 -0.000211116378257
Gc3_193 0 n6 ns193 0 7.75028663486e-05
Gc3_194 0 n6 ns194 0 0.00024063394599
Gc3_195 0 n6 ns195 0 0.00030291106423
Gc3_196 0 n6 ns196 0 -0.000187264814833
Gc3_197 0 n6 ns197 0 0.00136204509746
Gc3_198 0 n6 ns198 0 -0.000499873389697
Gc3_199 0 n6 ns199 0 0.000323604274111
Gc3_200 0 n6 ns200 0 -0.000369022089196
Gc3_201 0 n6 ns201 0 0.000377283602923
Gc3_202 0 n6 ns202 0 0.00080142672737
Gc3_203 0 n6 ns203 0 0.00172301423429
Gc3_204 0 n6 ns204 0 -0.000170187181398
Gc3_205 0 n6 ns205 0 -0.000173536527716
Gc3_206 0 n6 ns206 0 0.000868063737637
Gc3_207 0 n6 ns207 0 -0.00204356756211
Gc3_208 0 n6 ns208 0 -0.00315369487507
Gc3_209 0 n6 ns209 0 0.00173216358098
Gc3_210 0 n6 ns210 0 -0.00051109854389
Gc3_211 0 n6 ns211 0 0.000463032214832
Gc3_212 0 n6 ns212 0 -0.00155404922326
Gc3_213 0 n6 ns213 0 -0.00301822266666
Gc3_214 0 n6 ns214 0 -0.00012463896553
Gc3_215 0 n6 ns215 0 0.00557334346534
Gc3_216 0 n6 ns216 0 -0.000802966437319
Gc3_217 0 n6 ns217 0 -0.00270386162414
Gc3_218 0 n6 ns218 0 0.00218398693049
Gc3_219 0 n6 ns219 0 0.002304949487
Gc3_220 0 n6 ns220 0 0.0109193498218
Gc3_221 0 n6 ns221 0 -0.00211819832056
Gc3_222 0 n6 ns222 0 -5.61711356045e-06
Gc3_223 0 n6 ns223 0 -0.000168729706669
Gc3_224 0 n6 ns224 0 -0.00131117287392
Gc3_225 0 n6 ns225 0 -0.00103025462778
Gc3_226 0 n6 ns226 0 -3.60186643129e-06
Gc3_227 0 n6 ns227 0 -2.06145581856e-05
Gc3_228 0 n6 ns228 0 6.6502109123e-05
Gc3_229 0 n6 ns229 0 0.000263278158379
Gc3_230 0 n6 ns230 0 -0.00056545313395
Gc3_231 0 n6 ns231 0 -0.000213992039595
Gc3_232 0 n6 ns232 0 -0.000158432042984
Gc3_233 0 n6 ns233 0 0.00023253388788
Gc3_234 0 n6 ns234 0 -0.00282344387637
Gc3_235 0 n6 ns235 0 0.000637177068853
Gc3_236 0 n6 ns236 0 0.000253761585288
Gc3_237 0 n6 ns237 0 -0.000319909577047
Gc3_238 0 n6 ns238 0 -0.00075309825326
Gc3_239 0 n6 ns239 0 0.0006692752801
Gc3_240 0 n6 ns240 0 -0.00285371967956
Gc3_241 0 n6 ns241 0 0.00104238601274
Gc3_242 0 n6 ns242 0 -0.000243001594104
Gc3_243 0 n6 ns243 0 0.000799717798394
Gc3_244 0 n6 ns244 0 -0.00456487091617
Gc3_245 0 n6 ns245 0 0.00875766540616
Gc3_246 0 n6 ns246 0 -0.00313571584849
Gc3_247 0 n6 ns247 0 0.000914891880435
Gc3_248 0 n6 ns248 0 0.000198689328204
Gc3_249 0 n6 ns249 0 -0.00155528628521
Gc3_250 0 n6 ns250 0 0.0109722495229
Gc3_251 0 n6 ns251 0 0.024605271852
Gc3_252 0 n6 ns252 0 -0.0080843962465
Gc3_253 0 n6 ns253 0 0.00939471158656
Gc3_254 0 n6 ns254 0 -0.0021378001197
Gc3_255 0 n6 ns255 0 0.000688316941164
Gc3_256 0 n6 ns256 0 0.0574093948619
Gc3_257 0 n6 ns257 0 -0.00714700359866
Gc3_258 0 n6 ns258 0 -0.035508024946
Gc3_259 0 n6 ns259 0 2.10276864604e-05
Gc3_260 0 n6 ns260 0 0.00303855681907
Gc3_261 0 n6 ns261 0 -0.000983268823797
Gc3_262 0 n6 ns262 0 0.00068467243224
Gc3_263 0 n6 ns263 0 -2.12746305167e-05
Gc3_264 0 n6 ns264 0 -2.36731989038e-06
Gc3_265 0 n6 ns265 0 0.000433137852904
Gc3_266 0 n6 ns266 0 -0.000141332652281
Gc3_267 0 n6 ns267 0 -0.000643567406984
Gc3_268 0 n6 ns268 0 0.000754568520383
Gc3_269 0 n6 ns269 0 -0.000685288264493
Gc3_270 0 n6 ns270 0 0.000308917972015
Gc3_271 0 n6 ns271 0 0.00135627779759
Gc3_272 0 n6 ns272 0 0.000353934563579
Gc3_273 0 n6 ns273 0 0.000265682948426
Gc3_274 0 n6 ns274 0 -0.000379766799267
Gc3_275 0 n6 ns275 0 0.000439835611592
Gc3_276 0 n6 ns276 0 -0.000995177215422
Gc3_277 0 n6 ns277 0 -0.000733175090991
Gc3_278 0 n6 ns278 0 0.000943955602917
Gc3_279 0 n6 ns279 0 -0.000150302823961
Gc3_280 0 n6 ns280 0 0.000922028215722
Gc3_281 0 n6 ns281 0 0.0113027189114
Gc3_282 0 n6 ns282 0 -0.00591883395776
Gc3_283 0 n6 ns283 0 -0.00186547177872
Gc3_284 0 n6 ns284 0 -0.000100667006424
Gc3_285 0 n6 ns285 0 0.000367864536765
Gc3_286 0 n6 ns286 0 -0.00170214516583
Gc3_287 0 n6 ns287 0 -0.0025615881371
Gc3_288 0 n6 ns288 0 -0.0301002309576
Gc3_289 0 n6 ns289 0 -0.00433576365179
Gc3_290 0 n6 ns290 0 -0.010819133851
Gc3_291 0 n6 ns291 0 -0.0031149780577
Gc3_292 0 n6 ns292 0 0.0022383369035
Gc3_293 0 n6 ns293 0 -0.0150198138428
Gc3_294 0 n6 ns294 0 0.0127522892019
Gc3_295 0 n6 ns295 0 0.0181925103978
Gc3_296 0 n6 ns296 0 -1.23212392444e-05
Gd3_1 0 n6 ni1 0 -0.00085793373239
Gd3_2 0 n6 ni2 0 -0.00379334478599
Gd3_3 0 n6 ni3 0 -0.00264162384632
Gd3_4 0 n6 ni4 0 -0.00252227958497
Gd3_5 0 n6 ni5 0 0.00055145158742
Gd3_6 0 n6 ni6 0 -0.000536840959505
Gd3_7 0 n6 ni7 0 0.000563891773645
Gd3_8 0 n6 ni8 0 -0.000387208131844
Gc4_1 0 n8 ns1 0 0.00847015165182
Gc4_2 0 n8 ns2 0 -0.000945692160437
Gc4_3 0 n8 ns3 0 -0.000156415025753
Gc4_4 0 n8 ns4 0 -3.03632371845e-05
Gc4_5 0 n8 ns5 0 -1.19322879901e-05
Gc4_6 0 n8 ns6 0 0.000423610619785
Gc4_7 0 n8 ns7 0 -5.74635568409e-05
Gc4_8 0 n8 ns8 0 -0.000386445823419
Gc4_9 0 n8 ns9 0 0.00034356560092
Gc4_10 0 n8 ns10 0 -0.000178826535201
Gc4_11 0 n8 ns11 0 0.000564148281264
Gc4_12 0 n8 ns12 0 -0.00131703294615
Gc4_13 0 n8 ns13 0 -0.000788183493195
Gc4_14 0 n8 ns14 0 -0.000322514422006
Gc4_15 0 n8 ns15 0 0.000401992584672
Gc4_16 0 n8 ns16 0 -4.49266984551e-05
Gc4_17 0 n8 ns17 0 0.000471290765633
Gc4_18 0 n8 ns18 0 0.00129397130176
Gc4_19 0 n8 ns19 0 -0.000235411805685
Gc4_20 0 n8 ns20 0 -0.000219880819173
Gc4_21 0 n8 ns21 0 0.000900548524107
Gc4_22 0 n8 ns22 0 0.0013601923909
Gc4_23 0 n8 ns23 0 0.00103277775036
Gc4_24 0 n8 ns24 0 -0.00184579944344
Gc4_25 0 n8 ns25 0 0.000224234577564
Gc4_26 0 n8 ns26 0 -0.000407867869791
Gc4_27 0 n8 ns27 0 0.00153129149397
Gc4_28 0 n8 ns28 0 0.00387717706733
Gc4_29 0 n8 ns29 0 0.00593218908579
Gc4_30 0 n8 ns30 0 0.0100558491878
Gc4_31 0 n8 ns31 0 0.00164799855534
Gc4_32 0 n8 ns32 0 -0.00301940765426
Gc4_33 0 n8 ns33 0 0.00196009222188
Gc4_34 0 n8 ns34 0 -0.00197886593687
Gc4_35 0 n8 ns35 0 -0.0113338491922
Gc4_36 0 n8 ns36 0 0.00224891839654
Gc4_37 0 n8 ns37 0 4.36079607456e-06
Gc4_38 0 n8 ns38 0 0.00771492434885
Gc4_39 0 n8 ns39 0 -0.000608905282162
Gc4_40 0 n8 ns40 0 -0.000864652440546
Gc4_41 0 n8 ns41 0 -1.01158261112e-05
Gc4_42 0 n8 ns42 0 3.65373157579e-06
Gc4_43 0 n8 ns43 0 0.000334455178586
Gc4_44 0 n8 ns44 0 -7.04718180054e-05
Gc4_45 0 n8 ns45 0 -0.000327246029708
Gc4_46 0 n8 ns46 0 0.000416007121922
Gc4_47 0 n8 ns47 0 2.65089272376e-05
Gc4_48 0 n8 ns48 0 0.000271232737386
Gc4_49 0 n8 ns49 0 -0.00141125401438
Gc4_50 0 n8 ns50 0 2.27509224079e-05
Gc4_51 0 n8 ns51 0 -0.000382300506438
Gc4_52 0 n8 ns52 0 0.000444698958815
Gc4_53 0 n8 ns53 0 -0.000633141972289
Gc4_54 0 n8 ns54 0 -0.000107751930455
Gc4_55 0 n8 ns55 0 0.000703741806903
Gc4_56 0 n8 ns56 0 -0.000623052692199
Gc4_57 0 n8 ns57 0 -0.000316387973026
Gc4_58 0 n8 ns58 0 0.00100989948616
Gc4_59 0 n8 ns59 0 0.00104129550954
Gc4_60 0 n8 ns60 0 0.00234078416299
Gc4_61 0 n8 ns61 0 -0.000665229278378
Gc4_62 0 n8 ns62 0 0.000588408686307
Gc4_63 0 n8 ns63 0 -0.000535854146416
Gc4_64 0 n8 ns64 0 0.00193830648165
Gc4_65 0 n8 ns65 0 0.00278560195275
Gc4_66 0 n8 ns66 0 0.00555805749501
Gc4_67 0 n8 ns67 0 0.00542759302567
Gc4_68 0 n8 ns68 0 0.000520679132731
Gc4_69 0 n8 ns69 0 -0.00332866419986
Gc4_70 0 n8 ns70 0 0.00226496112377
Gc4_71 0 n8 ns71 0 -0.0136298502543
Gc4_72 0 n8 ns72 0 -0.0088738657283
Gc4_73 0 n8 ns73 0 0.00845547413975
Gc4_74 0 n8 ns74 0 3.66622370947e-06
Gc4_75 0 n8 ns75 0 0.0115985200059
Gc4_76 0 n8 ns76 0 -0.000514465096957
Gc4_77 0 n8 ns77 0 -0.00131513268143
Gc4_78 0 n8 ns78 0 -6.23289126914e-06
Gc4_79 0 n8 ns79 0 -6.33377274099e-06
Gc4_80 0 n8 ns80 0 0.000231626051467
Gc4_81 0 n8 ns81 0 -2.11134905379e-05
Gc4_82 0 n8 ns82 0 -0.000447847874508
Gc4_83 0 n8 ns83 0 -1.3510931791e-05
Gc4_84 0 n8 ns84 0 0.000307496720076
Gc4_85 0 n8 ns85 0 -7.77665239246e-05
Gc4_86 0 n8 ns86 0 0.000579620663901
Gc4_87 0 n8 ns87 0 -0.000128627232839
Gc4_88 0 n8 ns88 0 -0.000293271768156
Gc4_89 0 n8 ns89 0 0.000368772263516
Gc4_90 0 n8 ns90 0 9.63062725599e-05
Gc4_91 0 n8 ns91 0 -0.000851324413981
Gc4_92 0 n8 ns92 0 -0.00107558359101
Gc4_93 0 n8 ns93 0 0.000404443952956
Gc4_94 0 n8 ns94 0 -0.000196794190652
Gc4_95 0 n8 ns95 0 0.000876499288185
Gc4_96 0 n8 ns96 0 -0.00254383661785
Gc4_97 0 n8 ns97 0 0.000534949851281
Gc4_98 0 n8 ns98 0 0.00240926311875
Gc4_99 0 n8 ns99 0 -0.000237180970487
Gc4_100 0 n8 ns100 0 -0.000283884198527
Gc4_101 0 n8 ns101 0 0.00176471410329
Gc4_102 0 n8 ns102 0 -0.00286923731324
Gc4_103 0 n8 ns103 0 -0.00193752539855
Gc4_104 0 n8 ns104 0 -0.0077142983519
Gc4_105 0 n8 ns105 0 0.000202174546495
Gc4_106 0 n8 ns106 0 -0.00263727411666
Gc4_107 0 n8 ns107 0 0.00151510832131
Gc4_108 0 n8 ns108 0 -0.0187877350777
Gc4_109 0 n8 ns109 0 -0.00375997489481
Gc4_110 0 n8 ns110 0 0.00688057691749
Gc4_111 0 n8 ns111 0 5.2966230049e-06
Gc4_112 0 n8 ns112 0 0.00626729187278
Gc4_113 0 n8 ns113 0 0.000550062527733
Gc4_114 0 n8 ns114 0 -0.00123576642336
Gc4_115 0 n8 ns115 0 1.63960796966e-05
Gc4_116 0 n8 ns116 0 5.30454424871e-06
Gc4_117 0 n8 ns117 0 9.54952665481e-05
Gc4_118 0 n8 ns118 0 1.98833684096e-05
Gc4_119 0 n8 ns119 0 -0.000315933340673
Gc4_120 0 n8 ns120 0 0.000124896924126
Gc4_121 0 n8 ns121 0 0.000323665385875
Gc4_122 0 n8 ns122 0 -0.000160447418687
Gc4_123 0 n8 ns123 0 0.00015439198751
Gc4_124 0 n8 ns124 0 0.000505372911651
Gc4_125 0 n8 ns125 0 -0.000382817169018
Gc4_126 0 n8 ns126 0 0.000442738113626
Gc4_127 0 n8 ns127 0 -0.000145796456139
Gc4_128 0 n8 ns128 0 -0.000924349049638
Gc4_129 0 n8 ns129 0 -0.00080961772332
Gc4_130 0 n8 ns130 0 7.86109354346e-05
Gc4_131 0 n8 ns131 0 -0.000260636446395
Gc4_132 0 n8 ns132 0 0.00104382717953
Gc4_133 0 n8 ns133 0 -0.00261405391873
Gc4_134 0 n8 ns134 0 0.00102562170197
Gc4_135 0 n8 ns135 0 0.00170427290043
Gc4_136 0 n8 ns136 0 -0.000100271072489
Gc4_137 0 n8 ns137 0 -0.000396705091062
Gc4_138 0 n8 ns138 0 0.00196346199012
Gc4_139 0 n8 ns139 0 -0.00341714964157
Gc4_140 0 n8 ns140 0 -0.00354424065957
Gc4_141 0 n8 ns141 0 -0.00594496666546
Gc4_142 0 n8 ns142 0 -0.000898843655558
Gc4_143 0 n8 ns143 0 -0.00304640390693
Gc4_144 0 n8 ns144 0 0.00198219073321
Gc4_145 0 n8 ns145 0 -0.0143431114942
Gc4_146 0 n8 ns146 0 -0.00760555063245
Gc4_147 0 n8 ns147 0 0.00461369236465
Gc4_148 0 n8 ns148 0 1.06219180115e-05
Gc4_149 0 n8 ns149 0 0.000933487499133
Gc4_150 0 n8 ns150 0 0.00038937505109
Gc4_151 0 n8 ns151 0 0.000351882995622
Gc4_152 0 n8 ns152 0 1.04634986562e-05
Gc4_153 0 n8 ns153 0 1.20351097196e-05
Gc4_154 0 n8 ns154 0 1.72658692228e-05
Gc4_155 0 n8 ns155 0 -0.000211479338317
Gc4_156 0 n8 ns156 0 7.29462278743e-05
Gc4_157 0 n8 ns157 0 0.000241686096505
Gc4_158 0 n8 ns158 0 0.000303780122242
Gc4_159 0 n8 ns159 0 -0.000183800794875
Gc4_160 0 n8 ns160 0 0.00135689958194
Gc4_161 0 n8 ns161 0 -0.000519188513844
Gc4_162 0 n8 ns162 0 0.00032518694971
Gc4_163 0 n8 ns163 0 -0.00037236922922
Gc4_164 0 n8 ns164 0 0.000391805287513
Gc4_165 0 n8 ns165 0 0.00079340844986
Gc4_166 0 n8 ns166 0 0.00172930864818
Gc4_167 0 n8 ns167 0 -0.000184172982852
Gc4_168 0 n8 ns168 0 -0.000172591891936
Gc4_169 0 n8 ns169 0 0.000870976711613
Gc4_170 0 n8 ns170 0 -0.00204346984835
Gc4_171 0 n8 ns171 0 -0.00315591362412
Gc4_172 0 n8 ns172 0 0.00172345956781
Gc4_173 0 n8 ns173 0 -0.000521187813283
Gc4_174 0 n8 ns174 0 0.000458232717557
Gc4_175 0 n8 ns175 0 -0.00156025245671
Gc4_176 0 n8 ns176 0 -0.00302596904722
Gc4_177 0 n8 ns177 0 -0.000222189960796
Gc4_178 0 n8 ns178 0 0.00553342976554
Gc4_179 0 n8 ns179 0 -0.000864019358577
Gc4_180 0 n8 ns180 0 -0.00269632775276
Gc4_181 0 n8 ns181 0 0.00219445730496
Gc4_182 0 n8 ns182 0 0.00230619241874
Gc4_183 0 n8 ns183 0 0.0108965314128
Gc4_184 0 n8 ns184 0 -0.00210753972122
Gc4_185 0 n8 ns185 0 -5.63221940063e-06
Gc4_186 0 n8 ns186 0 0.00158428346909
Gc4_187 0 n8 ns187 0 -7.6849370123e-05
Gc4_188 0 n8 ns188 0 0.000451111171528
Gc4_189 0 n8 ns189 0 -5.92549503971e-06
Gc4_190 0 n8 ns190 0 1.18593865403e-05
Gc4_191 0 n8 ns191 0 0.000268202501949
Gc4_192 0 n8 ns192 0 -0.000187885552572
Gc4_193 0 n8 ns193 0 -0.000510091537752
Gc4_194 0 n8 ns194 0 0.000303461551089
Gc4_195 0 n8 ns195 0 -9.99379167571e-06
Gc4_196 0 n8 ns196 0 -1.16408850326e-05
Gc4_197 0 n8 ns197 0 0.00136081900411
Gc4_198 0 n8 ns198 0 -0.000155506684053
Gc4_199 0 n8 ns199 0 0.000395365509443
Gc4_200 0 n8 ns200 0 -0.000447125441786
Gc4_201 0 n8 ns201 0 0.000950133363232
Gc4_202 0 n8 ns202 0 0.000803075380803
Gc4_203 0 n8 ns203 0 0.00143918712765
Gc4_204 0 n8 ns204 0 0.000424903612536
Gc4_205 0 n8 ns205 0 -0.000188613639905
Gc4_206 0 n8 ns206 0 0.00103655721829
Gc4_207 0 n8 ns207 0 0.00105142419475
Gc4_208 0 n8 ns208 0 -0.00329539562019
Gc4_209 0 n8 ns209 0 0.001063468248
Gc4_210 0 n8 ns210 0 -0.000319900657459
Gc4_211 0 n8 ns211 0 0.000516853553019
Gc4_212 0 n8 ns212 0 -0.00184649841766
Gc4_213 0 n8 ns213 0 -0.00158201415644
Gc4_214 0 n8 ns214 0 -0.00706185853328
Gc4_215 0 n8 ns215 0 0.00450197454751
Gc4_216 0 n8 ns216 0 -0.00323119070504
Gc4_217 0 n8 ns217 0 -0.00327151989462
Gc4_218 0 n8 ns218 0 0.00253509644323
Gc4_219 0 n8 ns219 0 0.00173127457349
Gc4_220 0 n8 ns220 0 0.0128916648689
Gc4_221 0 n8 ns221 0 -0.000402179575642
Gc4_222 0 n8 ns222 0 -6.25908471199e-06
Gc4_223 0 n8 ns223 0 0.00303150678908
Gc4_224 0 n8 ns224 0 -0.000982506783468
Gc4_225 0 n8 ns225 0 0.000681028833823
Gc4_226 0 n8 ns226 0 -2.10745753434e-05
Gc4_227 0 n8 ns227 0 -2.41266559865e-06
Gc4_228 0 n8 ns228 0 0.000433821525707
Gc4_229 0 n8 ns229 0 -0.000142442011414
Gc4_230 0 n8 ns230 0 -0.000642636356262
Gc4_231 0 n8 ns231 0 0.000752675431397
Gc4_232 0 n8 ns232 0 -0.000686366971127
Gc4_233 0 n8 ns233 0 0.000308148061369
Gc4_234 0 n8 ns234 0 0.00135821544472
Gc4_235 0 n8 ns235 0 0.000356615637692
Gc4_236 0 n8 ns236 0 0.000265588709669
Gc4_237 0 n8 ns237 0 -0.000379873494989
Gc4_238 0 n8 ns238 0 0.000436163768826
Gc4_239 0 n8 ns239 0 -0.000993720651441
Gc4_240 0 n8 ns240 0 -0.000734531120852
Gc4_241 0 n8 ns241 0 0.000944599338052
Gc4_242 0 n8 ns242 0 -0.000150805263674
Gc4_243 0 n8 ns243 0 0.000922113956881
Gc4_244 0 n8 ns244 0 0.0113116494268
Gc4_245 0 n8 ns245 0 -0.00591799110289
Gc4_246 0 n8 ns246 0 -0.00186632389896
Gc4_247 0 n8 ns247 0 -0.000102376309593
Gc4_248 0 n8 ns248 0 0.000368425455578
Gc4_249 0 n8 ns249 0 -0.00170279517502
Gc4_250 0 n8 ns250 0 -0.00255149287899
Gc4_251 0 n8 ns251 0 -0.0301046056374
Gc4_252 0 n8 ns252 0 -0.00432755760469
Gc4_253 0 n8 ns253 0 -0.0108252547366
Gc4_254 0 n8 ns254 0 -0.00311677076708
Gc4_255 0 n8 ns255 0 0.00223942972342
Gc4_256 0 n8 ns256 0 -0.0149946460324
Gc4_257 0 n8 ns257 0 0.0127497465218
Gc4_258 0 n8 ns258 0 0.018170751951
Gc4_259 0 n8 ns259 0 -1.23142708465e-05
Gc4_260 0 n8 ns260 0 -0.0003377444936
Gc4_261 0 n8 ns261 0 -6.61515195215e-05
Gc4_262 0 n8 ns262 0 -0.00104924733972
Gc4_263 0 n8 ns263 0 1.54325057778e-05
Gc4_264 0 n8 ns264 0 -1.43124509986e-06
Gc4_265 0 n8 ns265 0 3.00868695131e-05
Gc4_266 0 n8 ns266 0 0.00016892428998
Gc4_267 0 n8 ns267 0 -0.000161604870288
Gc4_268 0 n8 ns268 0 -0.000247428999531
Gc4_269 0 n8 ns269 0 0.000318180371051
Gc4_270 0 n8 ns270 0 -0.000175621270885
Gc4_271 0 n8 ns271 0 -0.00237630508359
Gc4_272 0 n8 ns272 0 0.000214948690339
Gc4_273 0 n8 ns273 0 0.000378777455873
Gc4_274 0 n8 ns274 0 -0.000478760049267
Gc4_275 0 n8 ns275 0 -0.000625536664856
Gc4_276 0 n8 ns276 0 0.00120197469838
Gc4_277 0 n8 ns277 0 -0.00171385719168
Gc4_278 0 n8 ns278 0 0.000217393794517
Gc4_279 0 n8 ns279 0 -0.000314418047811
Gc4_280 0 n8 ns280 0 0.00106105059845
Gc4_281 0 n8 ns281 0 -0.00858039460359
Gc4_282 0 n8 ns282 0 0.00822723058237
Gc4_283 0 n8 ns283 0 -0.0018543263577
Gc4_284 0 n8 ns284 0 0.000279834640712
Gc4_285 0 n8 ns285 0 0.000427692592764
Gc4_286 0 n8 ns286 0 -0.00198435376631
Gc4_287 0 n8 ns287 0 0.00881730478052
Gc4_288 0 n8 ns288 0 0.0289700150658
Gc4_289 0 n8 ns289 0 -0.00491415028011
Gc4_290 0 n8 ns290 0 0.0100368764108
Gc4_291 0 n8 ns291 0 -0.00288762686827
Gc4_292 0 n8 ns292 0 0.00127809524102
Gc4_293 0 n8 ns293 0 0.0606085821254
Gc4_294 0 n8 ns294 0 -0.00370655028604
Gc4_295 0 n8 ns295 0 -0.0392998139483
Gc4_296 0 n8 ns296 0 1.74211205547e-05
Gd4_1 0 n8 ni1 0 -0.00378329761633
Gd4_2 0 n8 ni2 0 -0.00241578479749
Gd4_3 0 n8 ni3 0 -0.00252227959084
Gd4_4 0 n8 ni4 0 -0.000222291896074
Gd4_5 0 n8 ni5 0 -0.000550578024646
Gd4_6 0 n8 ni6 0 -0.000360951540129
Gd4_7 0 n8 ni7 0 -0.000383522687516
Gd4_8 0 n8 ni8 0 4.38357363666e-06
Gc5_1 0 n10 ns1 0 -0.000137579301957
Gc5_2 0 n10 ns2 0 -0.00131688852456
Gc5_3 0 n10 ns3 0 -0.00102576899885
Gc5_4 0 n10 ns4 0 -3.52957995164e-06
Gc5_5 0 n10 ns5 0 -2.05807589035e-05
Gc5_6 0 n10 ns6 0 6.89510110657e-05
Gc5_7 0 n10 ns7 0 0.000261083353452
Gc5_8 0 n10 ns8 0 -0.000570040339677
Gc5_9 0 n10 ns9 0 -0.0002123326455
Gc5_10 0 n10 ns10 0 -0.000160822558714
Gc5_11 0 n10 ns11 0 0.000237007525513
Gc5_12 0 n10 ns12 0 -0.00281942067931
Gc5_13 0 n10 ns13 0 0.000631987781029
Gc5_14 0 n10 ns14 0 0.000255810921456
Gc5_15 0 n10 ns15 0 -0.000324534255416
Gc5_16 0 n10 ns16 0 -0.000751490995487
Gc5_17 0 n10 ns17 0 0.00068189171364
Gc5_18 0 n10 ns18 0 -0.00284915402985
Gc5_19 0 n10 ns19 0 0.00105681770191
Gc5_20 0 n10 ns20 0 -0.000238168216064
Gc5_21 0 n10 ns21 0 0.00080914797865
Gc5_22 0 n10 ns22 0 -0.00459328755692
Gc5_23 0 n10 ns23 0 0.00873010482778
Gc5_24 0 n10 ns24 0 -0.0031354752304
Gc5_25 0 n10 ns25 0 0.000920313718897
Gc5_26 0 n10 ns26 0 0.000188696255545
Gc5_27 0 n10 ns27 0 -0.00156698126565
Gc5_28 0 n10 ns28 0 0.0109925809643
Gc5_29 0 n10 ns29 0 0.0246304680157
Gc5_30 0 n10 ns30 0 -0.00808679814023
Gc5_31 0 n10 ns31 0 0.00937920154365
Gc5_32 0 n10 ns32 0 -0.00212424101619
Gc5_33 0 n10 ns33 0 0.0007116423742
Gc5_34 0 n10 ns34 0 0.0575919942462
Gc5_35 0 n10 ns35 0 -0.00719689702972
Gc5_36 0 n10 ns36 0 -0.0356754949361
Gc5_37 0 n10 ns37 0 2.10961235033e-05
Gc5_38 0 n10 ns38 0 0.00308942158442
Gc5_39 0 n10 ns39 0 -0.000982873366439
Gc5_40 0 n10 ns40 0 0.000689655568556
Gc5_41 0 n10 ns41 0 -2.13649950333e-05
Gc5_42 0 n10 ns42 0 -2.2733383505e-06
Gc5_43 0 n10 ns43 0 0.000436598930485
Gc5_44 0 n10 ns44 0 -0.000142378741546
Gc5_45 0 n10 ns45 0 -0.000646471536518
Gc5_46 0 n10 ns46 0 0.000755857007439
Gc5_47 0 n10 ns47 0 -0.000684144397382
Gc5_48 0 n10 ns48 0 0.000312916595198
Gc5_49 0 n10 ns49 0 0.00135321634608
Gc5_50 0 n10 ns50 0 0.000339576728008
Gc5_51 0 n10 ns51 0 0.000267441961517
Gc5_52 0 n10 ns52 0 -0.000384320064494
Gc5_53 0 n10 ns53 0 0.000449625704327
Gc5_54 0 n10 ns54 0 -0.000994870026658
Gc5_55 0 n10 ns55 0 -0.000723634522879
Gc5_56 0 n10 ns56 0 0.000937539567461
Gc5_57 0 n10 ns57 0 -0.000149037250708
Gc5_58 0 n10 ns58 0 0.000926859358725
Gc5_59 0 n10 ns59 0 0.0113005431774
Gc5_60 0 n10 ns60 0 -0.00591516905025
Gc5_61 0 n10 ns61 0 -0.00186948737656
Gc5_62 0 n10 ns62 0 -0.000109109471316
Gc5_63 0 n10 ns63 0 0.000361779954454
Gc5_64 0 n10 ns64 0 -0.00171196992707
Gc5_65 0 n10 ns65 0 -0.00252873386382
Gc5_66 0 n10 ns66 0 -0.0301088556709
Gc5_67 0 n10 ns67 0 -0.00432233515521
Gc5_68 0 n10 ns68 0 -0.0108502729029
Gc5_69 0 n10 ns69 0 -0.00311111760993
Gc5_70 0 n10 ns70 0 0.00225380850319
Gc5_71 0 n10 ns71 0 -0.015009575386
Gc5_72 0 n10 ns72 0 0.0126980662783
Gc5_73 0 n10 ns73 0 0.0181943533505
Gc5_74 0 n10 ns74 0 -1.23297935014e-05
Gc5_75 0 n10 ns75 0 -0.00221425841049
Gc5_76 0 n10 ns76 0 0.000905823005616
Gc5_77 0 n10 ns77 0 2.36904682928e-05
Gc5_78 0 n10 ns78 0 2.10359807017e-05
Gc5_79 0 n10 ns79 0 2.41612055781e-05
Gc5_80 0 n10 ns80 0 -0.000170990089831
Gc5_81 0 n10 ns81 0 -0.00015589785327
Gc5_82 0 n10 ns82 0 -6.50263687262e-06
Gc5_83 0 n10 ns83 0 -0.000123244634917
Gc5_84 0 n10 ns84 0 0.000506095176696
Gc5_85 0 n10 ns85 0 -0.000397134148773
Gc5_86 0 n10 ns86 0 0.000955078373485
Gc5_87 0 n10 ns87 0 -0.000661855459688
Gc5_88 0 n10 ns88 0 0.000323339364132
Gc5_89 0 n10 ns89 0 -0.000315534548426
Gc5_90 0 n10 ns90 0 0.000915990989444
Gc5_91 0 n10 ns91 0 0.00104757025725
Gc5_92 0 n10 ns92 0 0.00237914187679
Gc5_93 0 n10 ns93 0 -0.00091713897636
Gc5_94 0 n10 ns94 0 -0.000174579827655
Gc5_95 0 n10 ns95 0 0.000698517133118
Gc5_96 0 n10 ns96 0 -0.00623738399264
Gc5_97 0 n10 ns97 0 0.000335356834862
Gc5_98 0 n10 ns98 0 0.00273381562019
Gc5_99 0 n10 ns99 0 -0.000668702630756
Gc5_100 0 n10 ns100 0 0.000425221838351
Gc5_101 0 n10 ns101 0 -0.00126604052208
Gc5_102 0 n10 ns102 0 -0.00268355743312
Gc5_103 0 n10 ns103 0 0.0102837126713
Gc5_104 0 n10 ns104 0 0.00761074592896
Gc5_105 0 n10 ns105 0 0.00327320907496
Gc5_106 0 n10 ns106 0 -0.00214889091126
Gc5_107 0 n10 ns107 0 0.0017498888734
Gc5_108 0 n10 ns108 0 0.00230678211658
Gc5_109 0 n10 ns109 0 0.00874268318039
Gc5_110 0 n10 ns110 0 -0.00331689342919
Gc5_111 0 n10 ns111 0 -4.86389493732e-06
Gc5_112 0 n10 ns112 0 0.000933487546695
Gc5_113 0 n10 ns113 0 0.000389375052394
Gc5_114 0 n10 ns114 0 0.000351883002892
Gc5_115 0 n10 ns115 0 1.04634983806e-05
Gc5_116 0 n10 ns116 0 1.20351096416e-05
Gc5_117 0 n10 ns117 0 1.72658720649e-05
Gc5_118 0 n10 ns118 0 -0.000211479338384
Gc5_119 0 n10 ns119 0 7.29462283333e-05
Gc5_120 0 n10 ns120 0 0.000241686096908
Gc5_121 0 n10 ns121 0 0.000303780122171
Gc5_122 0 n10 ns122 0 -0.000183800793545
Gc5_123 0 n10 ns123 0 0.0013568995819
Gc5_124 0 n10 ns124 0 -0.000519188517013
Gc5_125 0 n10 ns125 0 0.000325186949136
Gc5_126 0 n10 ns126 0 -0.000372369229437
Gc5_127 0 n10 ns127 0 0.000391805289638
Gc5_128 0 n10 ns128 0 0.00079340846526
Gc5_129 0 n10 ns129 0 0.00172930865395
Gc5_130 0 n10 ns130 0 -0.000184172970802
Gc5_131 0 n10 ns131 0 -0.000172591890426
Gc5_132 0 n10 ns132 0 0.000870976710371
Gc5_133 0 n10 ns133 0 -0.0020434698481
Gc5_134 0 n10 ns134 0 -0.00315591365162
Gc5_135 0 n10 ns135 0 0.00172345956409
Gc5_136 0 n10 ns136 0 -0.000521187819644
Gc5_137 0 n10 ns137 0 0.000458232718425
Gc5_138 0 n10 ns138 0 -0.0015602524586
Gc5_139 0 n10 ns139 0 -0.00302596898971
Gc5_140 0 n10 ns140 0 -0.00022219010454
Gc5_141 0 n10 ns141 0 0.00553342974287
Gc5_142 0 n10 ns142 0 -0.000864019460564
Gc5_143 0 n10 ns143 0 -0.00269632773729
Gc5_144 0 n10 ns144 0 0.00219445731743
Gc5_145 0 n10 ns145 0 0.00230619286802
Gc5_146 0 n10 ns146 0 0.0108965313453
Gc5_147 0 n10 ns147 0 -0.00210754012827
Gc5_148 0 n10 ns148 0 -5.63222034449e-06
Gc5_149 0 n10 ns149 0 0.0104639882963
Gc5_150 0 n10 ns150 0 0.000750601875772
Gc5_151 0 n10 ns151 0 -0.00106032082057
Gc5_152 0 n10 ns152 0 2.85124224113e-06
Gc5_153 0 n10 ns153 0 6.30163172807e-06
Gc5_154 0 n10 ns154 0 0.000104890291471
Gc5_155 0 n10 ns155 0 2.92820481523e-05
Gc5_156 0 n10 ns156 0 -0.000417303575204
Gc5_157 0 n10 ns157 0 2.99412818313e-06
Gc5_158 0 n10 ns158 0 0.000535921787356
Gc5_159 0 n10 ns159 0 -0.000217557488578
Gc5_160 0 n10 ns160 0 0.00078986163755
Gc5_161 0 n10 ns161 0 -0.000292941154481
Gc5_162 0 n10 ns162 0 -0.000205315941835
Gc5_163 0 n10 ns163 0 0.000285857293829
Gc5_164 0 n10 ns164 0 0.00065407214622
Gc5_165 0 n10 ns165 0 -0.00149503818957
Gc5_166 0 n10 ns166 0 -0.00124791748268
Gc5_167 0 n10 ns167 0 0.000757243986752
Gc5_168 0 n10 ns168 0 -0.000139118780804
Gc5_169 0 n10 ns169 0 0.000710814429537
Gc5_170 0 n10 ns170 0 -0.0054506837757
Gc5_171 0 n10 ns171 0 -0.000246464474034
Gc5_172 0 n10 ns172 0 0.00303264509624
Gc5_173 0 n10 ns173 0 -0.000398553824706
Gc5_174 0 n10 ns174 0 -0.000226591219995
Gc5_175 0 n10 ns175 0 0.00159581529386
Gc5_176 0 n10 ns176 0 -0.00678221002539
Gc5_177 0 n10 ns177 0 -0.00796292280967
Gc5_178 0 n10 ns178 0 -0.0128356443447
Gc5_179 0 n10 ns179 0 -0.00153827673759
Gc5_180 0 n10 ns180 0 -0.00195288599971
Gc5_181 0 n10 ns181 0 0.00145311565855
Gc5_182 0 n10 ns182 0 -0.0148016963023
Gc5_183 0 n10 ns183 0 -0.00268730427658
Gc5_184 0 n10 ns184 0 0.00319567496172
Gc5_185 0 n10 ns185 0 9.69851764178e-06
Gc5_186 0 n10 ns186 0 0.0115643732944
Gc5_187 0 n10 ns187 0 -0.000514011054883
Gc5_188 0 n10 ns188 0 -0.00133236209603
Gc5_189 0 n10 ns189 0 -5.74727699716e-06
Gc5_190 0 n10 ns190 0 -6.2793292342e-06
Gc5_191 0 n10 ns191 0 0.00023030961018
Gc5_192 0 n10 ns192 0 -2.46189845172e-05
Gc5_193 0 n10 ns193 0 -0.000439694347475
Gc5_194 0 n10 ns194 0 -1.00435801057e-05
Gc5_195 0 n10 ns195 0 0.000308448610536
Gc5_196 0 n10 ns196 0 -8.43204105671e-05
Gc5_197 0 n10 ns197 0 0.000580300215508
Gc5_198 0 n10 ns198 0 -9.15757119667e-05
Gc5_199 0 n10 ns199 0 -0.000293803088681
Gc5_200 0 n10 ns200 0 0.000371293553903
Gc5_201 0 n10 ns201 0 7.86296840041e-05
Gc5_202 0 n10 ns202 0 -0.000840566967134
Gc5_203 0 n10 ns203 0 -0.00108994602875
Gc5_204 0 n10 ns204 0 0.000396490740975
Gc5_205 0 n10 ns205 0 -0.000196046174616
Gc5_206 0 n10 ns206 0 0.000880449929454
Gc5_207 0 n10 ns207 0 -0.00252894565757
Gc5_208 0 n10 ns208 0 0.000543292411718
Gc5_209 0 n10 ns209 0 0.00243629458025
Gc5_210 0 n10 ns210 0 -0.000225870908038
Gc5_211 0 n10 ns211 0 -0.000274396580719
Gc5_212 0 n10 ns212 0 0.00177694321718
Gc5_213 0 n10 ns213 0 -0.00281395577547
Gc5_214 0 n10 ns214 0 -0.00196349808733
Gc5_215 0 n10 ns215 0 -0.00773815921036
Gc5_216 0 n10 ns216 0 0.000144538311903
Gc5_217 0 n10 ns217 0 -0.0026287894112
Gc5_218 0 n10 ns218 0 0.00153164925301
Gc5_219 0 n10 ns219 0 -0.0188195663565
Gc5_220 0 n10 ns220 0 -0.00373623749659
Gc5_221 0 n10 ns221 0 0.00689736006259
Gc5_222 0 n10 ns222 0 5.12767403887e-06
Gc5_223 0 n10 ns223 0 0.00222309576774
Gc5_224 0 n10 ns224 0 -0.000908844895864
Gc5_225 0 n10 ns225 0 -0.000432184367764
Gc5_226 0 n10 ns226 0 -1.22955657021e-05
Gc5_227 0 n10 ns227 0 -3.59374316374e-06
Gc5_228 0 n10 ns228 0 0.000196223428493
Gc5_229 0 n10 ns229 0 -9.30742508832e-05
Gc5_230 0 n10 ns230 0 -0.000135975399227
Gc5_231 0 n10 ns231 0 0.000585929496037
Gc5_232 0 n10 ns232 0 -0.000174103677463
Gc5_233 0 n10 ns233 0 0.0004693965434
Gc5_234 0 n10 ns234 0 -0.0020709806691
Gc5_235 0 n10 ns235 0 0.000335128817221
Gc5_236 0 n10 ns236 0 -0.000299256225282
Gc5_237 0 n10 ns237 0 0.000324821948714
Gc5_238 0 n10 ns238 0 -0.000796514527385
Gc5_239 0 n10 ns239 0 0.000684338865353
Gc5_240 0 n10 ns240 0 0.00144494997799
Gc5_241 0 n10 ns241 0 -0.00127266692473
Gc5_242 0 n10 ns242 0 -0.000267850476232
Gc5_243 0 n10 ns243 0 0.000752679346223
Gc5_244 0 n10 ns244 0 0.00356229759444
Gc5_245 0 n10 ns245 0 0.00266287568947
Gc5_246 0 n10 ns246 0 -0.00215123043264
Gc5_247 0 n10 ns247 0 0.00101799086567
Gc5_248 0 n10 ns248 0 -0.000405226778431
Gc5_249 0 n10 ns249 0 0.00141104479159
Gc5_250 0 n10 ns250 0 0.00496367708549
Gc5_251 0 n10 ns251 0 0.00968218889018
Gc5_252 0 n10 ns252 0 0.011160696832
Gc5_253 0 n10 ns253 0 0.00156743357591
Gc5_254 0 n10 ns254 0 -0.00244737451887
Gc5_255 0 n10 ns255 0 0.00182759168165
Gc5_256 0 n10 ns256 0 -0.0120004720911
Gc5_257 0 n10 ns257 0 -0.00846870645583
Gc5_258 0 n10 ns258 0 0.0118573374041
Gc5_259 0 n10 ns259 0 1.21167090674e-06
Gc5_260 0 n10 ns260 0 0.00852676892869
Gc5_261 0 n10 ns261 0 -0.000928228049606
Gc5_262 0 n10 ns262 0 -0.000139506469426
Gc5_263 0 n10 ns263 0 -3.11201037232e-05
Gc5_264 0 n10 ns264 0 -1.21075988414e-05
Gc5_265 0 n10 ns265 0 0.00042698115099
Gc5_266 0 n10 ns266 0 -5.50141331165e-05
Gc5_267 0 n10 ns267 0 -0.00038492558606
Gc5_268 0 n10 ns268 0 0.000345685513104
Gc5_269 0 n10 ns269 0 -0.000176254626833
Gc5_270 0 n10 ns270 0 0.000567016711224
Gc5_271 0 n10 ns271 0 -0.00132094625824
Gc5_272 0 n10 ns272 0 -0.000801205284274
Gc5_273 0 n10 ns273 0 -0.000321384898499
Gc5_274 0 n10 ns274 0 0.000400841302078
Gc5_275 0 n10 ns275 0 -2.95501934777e-05
Gc5_276 0 n10 ns276 0 0.000466137198319
Gc5_277 0 n10 ns277 0 0.00129895999476
Gc5_278 0 n10 ns278 0 -0.000228823874072
Gc5_279 0 n10 ns279 0 -0.000219517977456
Gc5_280 0 n10 ns280 0 0.000898798345041
Gc5_281 0 n10 ns281 0 0.00131931986583
Gc5_282 0 n10 ns282 0 0.00100473024368
Gc5_283 0 n10 ns283 0 -0.00184677050783
Gc5_284 0 n10 ns284 0 0.000222034416336
Gc5_285 0 n10 ns285 0 -0.000409236202225
Gc5_286 0 n10 ns286 0 0.00152844671467
Gc5_287 0 n10 ns287 0 0.00384986280559
Gc5_288 0 n10 ns288 0 0.00584019964521
Gc5_289 0 n10 ns289 0 0.0100307069332
Gc5_290 0 n10 ns290 0 0.00161681577175
Gc5_291 0 n10 ns291 0 -0.00302057749028
Gc5_292 0 n10 ns292 0 0.00196017501716
Gc5_293 0 n10 ns293 0 -0.00174893318784
Gc5_294 0 n10 ns294 0 -0.0113616010901
Gc5_295 0 n10 ns295 0 0.0020493166566
Gc5_296 0 n10 ns296 0 4.32728218551e-06
Gd5_1 0 n10 ni1 0 0.000552791703577
Gd5_2 0 n10 ni2 0 -0.000408981185784
Gd5_3 0 n10 ni3 0 0.000551451628771
Gd5_4 0 n10 ni4 0 -0.00055057805119
Gd5_5 0 n10 ni5 0 -0.00256983729392
Gd5_6 0 n10 ni6 0 -0.00252123010055
Gd5_7 0 n10 ni7 0 -0.00088416154234
Gd5_8 0 n10 ni8 0 -0.00381869966076
Gc6_1 0 n12 ns1 0 0.00307828984355
Gc6_2 0 n12 ns2 0 -0.00097863306228
Gc6_3 0 n12 ns3 0 0.000686667792336
Gc6_4 0 n12 ns4 0 -2.09924006919e-05
Gc6_5 0 n12 ns5 0 -2.16809900362e-06
Gc6_6 0 n12 ns6 0 0.000435801497886
Gc6_7 0 n12 ns7 0 -0.000143547058342
Gc6_8 0 n12 ns8 0 -0.000647475563171
Gc6_9 0 n12 ns9 0 0.000754299844093
Gc6_10 0 n12 ns10 0 -0.000683730866121
Gc6_11 0 n12 ns11 0 0.000313575463173
Gc6_12 0 n12 ns12 0 0.00135305506343
Gc6_13 0 n12 ns13 0 0.000342380563533
Gc6_14 0 n12 ns14 0 0.000267149396647
Gc6_15 0 n12 ns15 0 -0.000383475567639
Gc6_16 0 n12 ns16 0 0.000445476708839
Gc6_17 0 n12 ns17 0 -0.000996329304926
Gc6_18 0 n12 ns18 0 -0.000725658714299
Gc6_19 0 n12 ns19 0 0.000938988787008
Gc6_20 0 n12 ns20 0 -0.000149479519657
Gc6_21 0 n12 ns21 0 0.00092643667802
Gc6_22 0 n12 ns22 0 0.0112996385319
Gc6_23 0 n12 ns23 0 -0.00591408836641
Gc6_24 0 n12 ns24 0 -0.00186677247484
Gc6_25 0 n12 ns25 0 -0.00010972125936
Gc6_26 0 n12 ns26 0 0.000362921227606
Gc6_27 0 n12 ns27 0 -0.00171186339771
Gc6_28 0 n12 ns28 0 -0.00252591783869
Gc6_29 0 n12 ns29 0 -0.0301118096612
Gc6_30 0 n12 ns30 0 -0.00432126013705
Gc6_31 0 n12 ns31 0 -0.0108536224577
Gc6_32 0 n12 ns32 0 -0.00311158215992
Gc6_33 0 n12 ns33 0 0.00225422806517
Gc6_34 0 n12 ns34 0 -0.0149352910569
Gc6_35 0 n12 ns35 0 0.0127056777947
Gc6_36 0 n12 ns36 0 0.0181232301954
Gc6_37 0 n12 ns37 0 -1.22184931914e-05
Gc6_38 0 n12 ns38 0 -0.000328800773058
Gc6_39 0 n12 ns39 0 -5.05393124991e-05
Gc6_40 0 n12 ns40 0 -0.0010453750726
Gc6_41 0 n12 ns41 0 1.56091714957e-05
Gc6_42 0 n12 ns42 0 -1.21897217731e-06
Gc6_43 0 n12 ns43 0 3.06285679136e-05
Gc6_44 0 n12 ns44 0 0.000168642063633
Gc6_45 0 n12 ns45 0 -0.00016205842494
Gc6_46 0 n12 ns46 0 -0.000246470266013
Gc6_47 0 n12 ns47 0 0.000321736718856
Gc6_48 0 n12 ns48 0 -0.000176097839587
Gc6_49 0 n12 ns49 0 -0.00237938449622
Gc6_50 0 n12 ns50 0 0.000207305800511
Gc6_51 0 n12 ns51 0 0.000379690341881
Gc6_52 0 n12 ns52 0 -0.000480273718844
Gc6_53 0 n12 ns53 0 -0.00062515352053
Gc6_54 0 n12 ns54 0 0.00119403780825
Gc6_55 0 n12 ns55 0 -0.00171497652798
Gc6_56 0 n12 ns56 0 0.000207316662931
Gc6_57 0 n12 ns57 0 -0.000314316858445
Gc6_58 0 n12 ns58 0 0.00106355475892
Gc6_59 0 n12 ns59 0 -0.00857417663267
Gc6_60 0 n12 ns60 0 0.00821160626529
Gc6_61 0 n12 ns61 0 -0.00185942135409
Gc6_62 0 n12 ns62 0 0.000269882730741
Gc6_63 0 n12 ns63 0 0.000426762337141
Gc6_64 0 n12 ns64 0 -0.00198927506292
Gc6_65 0 n12 ns65 0 0.00880745859063
Gc6_66 0 n12 ns66 0 0.0288486658558
Gc6_67 0 n12 ns67 0 -0.00495336047657
Gc6_68 0 n12 ns68 0 0.00996243978884
Gc6_69 0 n12 ns69 0 -0.00288268758487
Gc6_70 0 n12 ns70 0 0.00128771199527
Gc6_71 0 n12 ns71 0 0.0606554496901
Gc6_72 0 n12 ns72 0 -0.00372057862382
Gc6_73 0 n12 ns73 0 -0.0393302562375
Gc6_74 0 n12 ns74 0 1.74002036435e-05
Gc6_75 0 n12 ns75 0 0.000905682087216
Gc6_76 0 n12 ns76 0 0.000379093840812
Gc6_77 0 n12 ns77 0 0.000343390703059
Gc6_78 0 n12 ns78 0 1.05182792646e-05
Gc6_79 0 n12 ns79 0 1.19235005643e-05
Gc6_80 0 n12 ns80 0 1.582752165e-05
Gc6_81 0 n12 ns81 0 -0.000211116378347
Gc6_82 0 n12 ns82 0 7.75028666603e-05
Gc6_83 0 n12 ns83 0 0.000240633946104
Gc6_84 0 n12 ns84 0 0.000302911064319
Gc6_85 0 n12 ns85 0 -0.00018726481503
Gc6_86 0 n12 ns86 0 0.00136204509813
Gc6_87 0 n12 ns87 0 -0.00049987338927
Gc6_88 0 n12 ns88 0 0.000323604273869
Gc6_89 0 n12 ns89 0 -0.000369022089274
Gc6_90 0 n12 ns90 0 0.000377283601059
Gc6_91 0 n12 ns91 0 0.000801426731897
Gc6_92 0 n12 ns92 0 0.00172301423338
Gc6_93 0 n12 ns93 0 -0.00017018717814
Gc6_94 0 n12 ns94 0 -0.000173536527521
Gc6_95 0 n12 ns95 0 0.000868063737717
Gc6_96 0 n12 ns96 0 -0.00204356754607
Gc6_97 0 n12 ns97 0 -0.00315369488886
Gc6_98 0 n12 ns98 0 0.00173216357716
Gc6_99 0 n12 ns99 0 -0.000511098552651
Gc6_100 0 n12 ns100 0 0.000463032216482
Gc6_101 0 n12 ns101 0 -0.00155404922612
Gc6_102 0 n12 ns102 0 -0.00301822264386
Gc6_103 0 n12 ns103 0 -0.000124639083651
Gc6_104 0 n12 ns104 0 0.0055733434367
Gc6_105 0 n12 ns105 0 -0.000802966498383
Gc6_106 0 n12 ns106 0 -0.00270386161897
Gc6_107 0 n12 ns107 0 0.00218398693379
Gc6_108 0 n12 ns108 0 0.00230494976472
Gc6_109 0 n12 ns109 0 0.0109193497889
Gc6_110 0 n12 ns110 0 -0.00211819857044
Gc6_111 0 n12 ns111 0 -5.61711393022e-06
Gc6_112 0 n12 ns112 0 0.00158428345394
Gc6_113 0 n12 ns113 0 -7.68493767954e-05
Gc6_114 0 n12 ns114 0 0.00045111116393
Gc6_115 0 n12 ns115 0 -5.92549492297e-06
Gc6_116 0 n12 ns116 0 1.18593865782e-05
Gc6_117 0 n12 ns117 0 0.000268202500844
Gc6_118 0 n12 ns118 0 -0.000187885552716
Gc6_119 0 n12 ns119 0 -0.00051009153763
Gc6_120 0 n12 ns120 0 0.000303461550558
Gc6_121 0 n12 ns121 0 -9.99379161299e-06
Gc6_122 0 n12 ns122 0 -1.16408859353e-05
Gc6_123 0 n12 ns123 0 0.00136081900407
Gc6_124 0 n12 ns124 0 -0.000155506680975
Gc6_125 0 n12 ns125 0 0.0003953655096
Gc6_126 0 n12 ns126 0 -0.000447125441829
Gc6_127 0 n12 ns127 0 0.000950133359856
Gc6_128 0 n12 ns128 0 0.000803075372746
Gc6_129 0 n12 ns129 0 0.00143918712419
Gc6_130 0 n12 ns130 0 0.000424903605972
Gc6_131 0 n12 ns131 0 -0.000188613640765
Gc6_132 0 n12 ns132 0 0.00103655721871
Gc6_133 0 n12 ns133 0 0.00105142419561
Gc6_134 0 n12 ns134 0 -0.0032953955938
Gc6_135 0 n12 ns135 0 0.00106346825255
Gc6_136 0 n12 ns136 0 -0.000319900653373
Gc6_137 0 n12 ns137 0 0.000516853552638
Gc6_138 0 n12 ns138 0 -0.00184649841582
Gc6_139 0 n12 ns139 0 -0.00158201419307
Gc6_140 0 n12 ns140 0 -0.00706185838031
Gc6_141 0 n12 ns141 0 0.0045019745791
Gc6_142 0 n12 ns142 0 -0.00323119060682
Gc6_143 0 n12 ns143 0 -0.00327151990457
Gc6_144 0 n12 ns144 0 0.00253509643354
Gc6_145 0 n12 ns145 0 0.00173127418121
Gc6_146 0 n12 ns146 0 0.0128916649184
Gc6_147 0 n12 ns147 0 -0.00040217922546
Gc6_148 0 n12 ns148 0 -6.25908414951e-06
Gc6_149 0 n12 ns149 0 0.0115643733094
Gc6_150 0 n12 ns150 0 -0.000514011053227
Gc6_151 0 n12 ns151 0 -0.00133236209386
Gc6_152 0 n12 ns152 0 -5.74727703462e-06
Gc6_153 0 n12 ns153 0 -6.27932927583e-06
Gc6_154 0 n12 ns154 0 0.000230309610839
Gc6_155 0 n12 ns155 0 -2.46189847756e-05
Gc6_156 0 n12 ns156 0 -0.000439694348022
Gc6_157 0 n12 ns157 0 -1.00435803397e-05
Gc6_158 0 n12 ns158 0 0.00030844860989
Gc6_159 0 n12 ns159 0 -8.43204095778e-05
Gc6_160 0 n12 ns160 0 0.0005803002161
Gc6_161 0 n12 ns161 0 -9.15757153772e-05
Gc6_162 0 n12 ns162 0 -0.000293803088715
Gc6_163 0 n12 ns163 0 0.000371293553984
Gc6_164 0 n12 ns164 0 7.86296886231e-05
Gc6_165 0 n12 ns165 0 -0.000840566961473
Gc6_166 0 n12 ns166 0 -0.00108994602396
Gc6_167 0 n12 ns167 0 0.000396490745544
Gc6_168 0 n12 ns168 0 -0.000196046173787
Gc6_169 0 n12 ns169 0 0.000880449928795
Gc6_170 0 n12 ns170 0 -0.00252894567568
Gc6_171 0 n12 ns171 0 0.000543292401038
Gc6_172 0 n12 ns172 0 0.00243629457934
Gc6_173 0 n12 ns173 0 -0.000225870902288
Gc6_174 0 n12 ns174 0 -0.000274396582793
Gc6_175 0 n12 ns175 0 0.00177694321855
Gc6_176 0 n12 ns176 0 -0.00281395578762
Gc6_177 0 n12 ns177 0 -0.00196349806864
Gc6_178 0 n12 ns178 0 -0.00773815920888
Gc6_179 0 n12 ns179 0 0.000144538328959
Gc6_180 0 n12 ns180 0 -0.00262878940857
Gc6_181 0 n12 ns181 0 0.00153164925042
Gc6_182 0 n12 ns182 0 -0.018819566234
Gc6_183 0 n12 ns183 0 -0.00373623748844
Gc6_184 0 n12 ns184 0 0.0068973599444
Gc6_185 0 n12 ns185 0 5.12767372812e-06
Gc6_186 0 n12 ns186 0 0.00623363575244
Gc6_187 0 n12 ns187 0 0.000544732406249
Gc6_188 0 n12 ns188 0 -0.00124176837539
Gc6_189 0 n12 ns189 0 1.6301586585e-05
Gc6_190 0 n12 ns190 0 5.10249984796e-06
Gc6_191 0 n12 ns191 0 9.66511975894e-05
Gc6_192 0 n12 ns192 0 1.87600524262e-05
Gc6_193 0 n12 ns193 0 -0.000314826339092
Gc6_194 0 n12 ns194 0 0.000122345059758
Gc6_195 0 n12 ns195 0 0.000324098126281
Gc6_196 0 n12 ns196 0 -0.000160183984106
Gc6_197 0 n12 ns197 0 0.00015196653225
Gc6_198 0 n12 ns198 0 0.000506133312062
Gc6_199 0 n12 ns199 0 -0.000383984781657
Gc6_200 0 n12 ns200 0 0.000442609217535
Gc6_201 0 n12 ns201 0 -0.000150080106882
Gc6_202 0 n12 ns202 0 -0.000923981162147
Gc6_203 0 n12 ns203 0 -0.00079851741137
Gc6_204 0 n12 ns204 0 7.74366738185e-05
Gc6_205 0 n12 ns205 0 -0.000260391554572
Gc6_206 0 n12 ns206 0 0.00104377093278
Gc6_207 0 n12 ns207 0 -0.0026138819893
Gc6_208 0 n12 ns208 0 0.00106930483237
Gc6_209 0 n12 ns209 0 0.00170172917935
Gc6_210 0 n12 ns210 0 -9.08228338604e-05
Gc6_211 0 n12 ns211 0 -0.000395613596796
Gc6_212 0 n12 ns212 0 0.00196552071347
Gc6_213 0 n12 ns213 0 -0.00343912048604
Gc6_214 0 n12 ns214 0 -0.00331200019597
Gc6_215 0 n12 ns215 0 -0.00588064691936
Gc6_216 0 n12 ns216 0 -0.000779208724213
Gc6_217 0 n12 ns217 0 -0.00305331632012
Gc6_218 0 n12 ns218 0 0.00197062039799
Gc6_219 0 n12 ns219 0 -0.0146478074327
Gc6_220 0 n12 ns220 0 -0.00749476974573
Gc6_221 0 n12 ns221 0 0.00485362326973
Gc6_222 0 n12 ns222 0 1.08795361578e-05
Gc6_223 0 n12 ns223 0 0.0085002042265
Gc6_224 0 n12 ns224 0 -0.000923039394763
Gc6_225 0 n12 ns225 0 -0.000142275732491
Gc6_226 0 n12 ns226 0 -3.09337040581e-05
Gc6_227 0 n12 ns227 0 -1.21788060156e-05
Gc6_228 0 n12 ns228 0 0.000426409625326
Gc6_229 0 n12 ns229 0 -5.52139534784e-05
Gc6_230 0 n12 ns230 0 -0.000384958020956
Gc6_231 0 n12 ns231 0 0.000341008198228
Gc6_232 0 n12 ns232 0 -0.000177089367643
Gc6_233 0 n12 ns233 0 0.000562304041026
Gc6_234 0 n12 ns234 0 -0.00130874933928
Gc6_235 0 n12 ns235 0 -0.000803030451308
Gc6_236 0 n12 ns236 0 -0.0003215081255
Gc6_237 0 n12 ns237 0 0.000398903179028
Gc6_238 0 n12 ns238 0 -2.63449109862e-05
Gc6_239 0 n12 ns239 0 0.000464598900806
Gc6_240 0 n12 ns240 0 0.00129596490321
Gc6_241 0 n12 ns241 0 -0.000225465479282
Gc6_242 0 n12 ns242 0 -0.000219942012841
Gc6_243 0 n12 ns243 0 0.000897121238496
Gc6_244 0 n12 ns244 0 0.00131774501399
Gc6_245 0 n12 ns245 0 0.0010064556209
Gc6_246 0 n12 ns246 0 -0.00185267175981
Gc6_247 0 n12 ns247 0 0.000208725251644
Gc6_248 0 n12 ns248 0 -0.000413636881133
Gc6_249 0 n12 ns249 0 0.00152093287402
Gc6_250 0 n12 ns250 0 0.00384455030667
Gc6_251 0 n12 ns251 0 0.00583030866028
Gc6_252 0 n12 ns252 0 0.010040748535
Gc6_253 0 n12 ns253 0 0.00163090263344
Gc6_254 0 n12 ns254 0 -0.00302428064398
Gc6_255 0 n12 ns255 0 0.00195196162825
Gc6_256 0 n12 ns256 0 -0.00163393752972
Gc6_257 0 n12 ns257 0 -0.0113898752061
Gc6_258 0 n12 ns258 0 0.00195369983917
Gc6_259 0 n12 ns259 0 4.2408698666e-06
Gc6_260 0 n12 ns260 0 0.00763103526118
Gc6_261 0 n12 ns261 0 -0.000573185943796
Gc6_262 0 n12 ns262 0 -0.000855495858013
Gc6_263 0 n12 ns263 0 -9.95962601353e-06
Gc6_264 0 n12 ns264 0 3.80612738148e-06
Gc6_265 0 n12 ns265 0 0.000331062299426
Gc6_266 0 n12 ns266 0 -7.03325565204e-05
Gc6_267 0 n12 ns267 0 -0.00032584670741
Gc6_268 0 n12 ns268 0 0.000417831692218
Gc6_269 0 n12 ns269 0 2.94155153516e-05
Gc6_270 0 n12 ns270 0 0.000270419712958
Gc6_271 0 n12 ns271 0 -0.00142356905501
Gc6_272 0 n12 ns272 0 2.70182179118e-05
Gc6_273 0 n12 ns273 0 -0.000381569897997
Gc6_274 0 n12 ns274 0 0.000443826035975
Gc6_275 0 n12 ns275 0 -0.00062874558386
Gc6_276 0 n12 ns276 0 -0.000123278965226
Gc6_277 0 n12 ns277 0 0.000703627729107
Gc6_278 0 n12 ns278 0 -0.000631581147589
Gc6_279 0 n12 ns279 0 -0.00031596247109
Gc6_280 0 n12 ns280 0 0.00100921080945
Gc6_281 0 n12 ns281 0 0.000994903893788
Gc6_282 0 n12 ns282 0 0.00234481518302
Gc6_283 0 n12 ns283 0 -0.000659995517015
Gc6_284 0 n12 ns284 0 0.000593730798392
Gc6_285 0 n12 ns285 0 -0.000538812219621
Gc6_286 0 n12 ns286 0 0.00193931290745
Gc6_287 0 n12 ns287 0 0.00274526275132
Gc6_288 0 n12 ns288 0 0.00545266882734
Gc6_289 0 n12 ns289 0 0.00537521539608
Gc6_290 0 n12 ns290 0 0.000465410141255
Gc6_291 0 n12 ns291 0 -0.00332333859353
Gc6_292 0 n12 ns292 0 0.00226922545529
Gc6_293 0 n12 ns293 0 -0.0134095472817
Gc6_294 0 n12 ns294 0 -0.00888982595943
Gc6_295 0 n12 ns295 0 0.00826425512021
Gc6_296 0 n12 ns296 0 3.93530928412e-06
Gd6_1 0 n12 ni1 0 -0.00040589925805
Gd6_2 0 n12 ni2 0 -4.81368386918e-06
Gd6_3 0 n12 ni3 0 -0.000536840965277
Gd6_4 0 n12 ni4 0 -0.000360951529315
Gd6_5 0 n12 ni5 0 -0.00252123010927
Gd6_6 0 n12 ni6 0 -0.000163493682934
Gd6_7 0 n12 ni7 0 -0.00380616257058
Gd6_8 0 n12 ni8 0 -0.00239559162195
Gc7_1 0 n14 ns1 0 -0.00219636682013
Gc7_2 0 n14 ns2 0 0.000886758456026
Gc7_3 0 n14 ns3 0 1.08742981357e-05
Gc7_4 0 n14 ns4 0 2.08387022317e-05
Gc7_5 0 n14 ns5 0 2.39386819527e-05
Gc7_6 0 n14 ns6 0 -0.000170759883627
Gc7_7 0 n14 ns7 0 -0.000156196909034
Gc7_8 0 n14 ns8 0 -3.56763594673e-06
Gc7_9 0 n14 ns9 0 -0.000122465961025
Gc7_10 0 n14 ns10 0 0.000508298305837
Gc7_11 0 n14 ns11 0 -0.000402918271409
Gc7_12 0 n14 ns12 0 0.000961538488497
Gc7_13 0 n14 ns13 0 -0.000648406302267
Gc7_14 0 n14 ns14 0 0.000322566049506
Gc7_15 0 n14 ns15 0 -0.000316233934317
Gc7_16 0 n14 ns16 0 0.00090081950713
Gc7_17 0 n14 ns17 0 0.00105568815351
Gc7_18 0 n14 ns18 0 0.002371598113
Gc7_19 0 n14 ns19 0 -0.000915009049568
Gc7_20 0 n14 ns20 0 -0.000175080523599
Gc7_21 0 n14 ns21 0 0.000700317444818
Gc7_22 0 n14 ns22 0 -0.00619986618675
Gc7_23 0 n14 ns23 0 0.000345448855405
Gc7_24 0 n14 ns24 0 0.00273647140486
Gc7_25 0 n14 ns25 0 -0.000677324707839
Gc7_26 0 n14 ns26 0 0.000427347190276
Gc7_27 0 n14 ns27 0 -0.00126808616981
Gc7_28 0 n14 ns28 0 -0.00262718067155
Gc7_29 0 n14 ns29 0 0.0103353074573
Gc7_30 0 n14 ns30 0 0.00765271997994
Gc7_31 0 n14 ns31 0 0.00328242414464
Gc7_32 0 n14 ns32 0 -0.00215360499624
Gc7_33 0 n14 ns33 0 0.00175095931212
Gc7_34 0 n14 ns34 0 0.00225573941108
Gc7_35 0 n14 ns35 0 0.00875848189526
Gc7_36 0 n14 ns36 0 -0.00327727895151
Gc7_37 0 n14 ns37 0 -4.89664041398e-06
Gc7_38 0 n14 ns38 0 0.000899858123978
Gc7_39 0 n14 ns39 0 0.000384024670034
Gc7_40 0 n14 ns40 0 0.000348907034368
Gc7_41 0 n14 ns41 0 1.05747324867e-05
Gc7_42 0 n14 ns42 0 1.19296061066e-05
Gc7_43 0 n14 ns43 0 1.55695213494e-05
Gc7_44 0 n14 ns44 0 -0.000211320393977
Gc7_45 0 n14 ns45 0 7.58481516433e-05
Gc7_46 0 n14 ns46 0 0.00024038108974
Gc7_47 0 n14 ns47 0 0.000301315896229
Gc7_48 0 n14 ns48 0 -0.000185065256652
Gc7_49 0 n14 ns49 0 0.00135994501656
Gc7_50 0 n14 ns50 0 -0.000506797566576
Gc7_51 0 n14 ns51 0 0.000324046315384
Gc7_52 0 n14 ns52 0 -0.000369211828655
Gc7_53 0 n14 ns53 0 0.000381180279099
Gc7_54 0 n14 ns54 0 0.000797227016045
Gc7_55 0 n14 ns55 0 0.00172319104659
Gc7_56 0 n14 ns56 0 -0.000170912615297
Gc7_57 0 n14 ns57 0 -0.000173175546441
Gc7_58 0 n14 ns58 0 0.000867915338587
Gc7_59 0 n14 ns59 0 -0.00204894058119
Gc7_60 0 n14 ns60 0 -0.00316342922119
Gc7_61 0 n14 ns61 0 0.00172826299739
Gc7_62 0 n14 ns62 0 -0.000510009950037
Gc7_63 0 n14 ns63 0 0.000461669285281
Gc7_64 0 n14 ns64 0 -0.00155431399879
Gc7_65 0 n14 ns65 0 -0.00302899080179
Gc7_66 0 n14 ns66 0 -0.000174317025398
Gc7_67 0 n14 ns67 0 0.0055540535134
Gc7_68 0 n14 ns68 0 -0.000825870597396
Gc7_69 0 n14 ns69 0 -0.00270145375484
Gc7_70 0 n14 ns70 0 0.00218514941239
Gc7_71 0 n14 ns71 0 0.00238937460089
Gc7_72 0 n14 ns72 0 0.0109090948003
Gc7_73 0 n14 ns73 0 -0.00219023722942
Gc7_74 0 n14 ns74 0 -5.57496306799e-06
Gc7_75 0 n14 ns75 0 -0.000168729708317
Gc7_76 0 n14 ns76 0 -0.00131117287151
Gc7_77 0 n14 ns77 0 -0.00103025462747
Gc7_78 0 n14 ns78 0 -3.60186641902e-06
Gc7_79 0 n14 ns79 0 -2.061455814e-05
Gc7_80 0 n14 ns80 0 6.65021090611e-05
Gc7_81 0 n14 ns81 0 0.000263278158779
Gc7_82 0 n14 ns82 0 -0.000565453134014
Gc7_83 0 n14 ns83 0 -0.000213992038909
Gc7_84 0 n14 ns84 0 -0.000158432042213
Gc7_85 0 n14 ns85 0 0.000232533888507
Gc7_86 0 n14 ns86 0 -0.00282344387899
Gc7_87 0 n14 ns87 0 0.000637177068853
Gc7_88 0 n14 ns88 0 0.00025376158536
Gc7_89 0 n14 ns89 0 -0.000319909577207
Gc7_90 0 n14 ns90 0 -0.000753098253167
Gc7_91 0 n14 ns91 0 0.000669275277292
Gc7_92 0 n14 ns92 0 -0.00285371967964
Gc7_93 0 n14 ns93 0 0.00104238601083
Gc7_94 0 n14 ns94 0 -0.000243001594353
Gc7_95 0 n14 ns95 0 0.000799717798355
Gc7_96 0 n14 ns96 0 -0.00456487091689
Gc7_97 0 n14 ns97 0 0.00875766540991
Gc7_98 0 n14 ns98 0 -0.00313571584941
Gc7_99 0 n14 ns99 0 0.000914891879865
Gc7_100 0 n14 ns100 0 0.000198689327874
Gc7_101 0 n14 ns101 0 -0.00155528628584
Gc7_102 0 n14 ns102 0 0.0109722494966
Gc7_103 0 n14 ns103 0 0.0246052718675
Gc7_104 0 n14 ns104 0 -0.00808439625713
Gc7_105 0 n14 ns105 0 0.00939471161311
Gc7_106 0 n14 ns106 0 -0.00213780011902
Gc7_107 0 n14 ns107 0 0.000688316935833
Gc7_108 0 n14 ns108 0 0.0574093948292
Gc7_109 0 n14 ns109 0 -0.00714700359066
Gc7_110 0 n14 ns110 0 -0.0355080249191
Gc7_111 0 n14 ns111 0 2.10276865379e-05
Gc7_112 0 n14 ns112 0 0.00303150677888
Gc7_113 0 n14 ns113 0 -0.00098250678289
Gc7_114 0 n14 ns114 0 0.000681028832938
Gc7_115 0 n14 ns115 0 -2.10745752185e-05
Gc7_116 0 n14 ns116 0 -2.41266558876e-06
Gc7_117 0 n14 ns117 0 0.000433821525049
Gc7_118 0 n14 ns118 0 -0.000142442011635
Gc7_119 0 n14 ns119 0 -0.000642636356395
Gc7_120 0 n14 ns120 0 0.00075267543097
Gc7_121 0 n14 ns121 0 -0.000686366971637
Gc7_122 0 n14 ns122 0 0.000308148060757
Gc7_123 0 n14 ns123 0 0.00135821544629
Gc7_124 0 n14 ns124 0 0.000356615637755
Gc7_125 0 n14 ns125 0 0.000265588709825
Gc7_126 0 n14 ns126 0 -0.000379873494816
Gc7_127 0 n14 ns127 0 0.0004361637696
Gc7_128 0 n14 ns128 0 -0.000993720653219
Gc7_129 0 n14 ns129 0 -0.000734531121224
Gc7_130 0 n14 ns130 0 0.000944599336551
Gc7_131 0 n14 ns131 0 -0.000150805263807
Gc7_132 0 n14 ns132 0 0.000922113957109
Gc7_133 0 n14 ns133 0 0.0113116494229
Gc7_134 0 n14 ns134 0 -0.00591799110031
Gc7_135 0 n14 ns135 0 -0.00186632389737
Gc7_136 0 n14 ns136 0 -0.0001023763059
Gc7_137 0 n14 ns137 0 0.000368425454942
Gc7_138 0 n14 ns138 0 -0.00170279517353
Gc7_139 0 n14 ns139 0 -0.002551492861
Gc7_140 0 n14 ns140 0 -0.0301046056133
Gc7_141 0 n14 ns141 0 -0.00432755757835
Gc7_142 0 n14 ns142 0 -0.0108252547348
Gc7_143 0 n14 ns143 0 -0.00311677077334
Gc7_144 0 n14 ns144 0 0.00223942972397
Gc7_145 0 n14 ns145 0 -0.0149946459664
Gc7_146 0 n14 ns146 0 0.0127497465448
Gc7_147 0 n14 ns147 0 0.0181707518895
Gc7_148 0 n14 ns148 0 -1.23142701838e-05
Gc7_149 0 n14 ns149 0 0.0022230959179
Gc7_150 0 n14 ns150 0 -0.000908844990211
Gc7_151 0 n14 ns151 0 -0.000432184389499
Gc7_152 0 n14 ns152 0 -1.22955663467e-05
Gc7_153 0 n14 ns153 0 -3.59374343604e-06
Gc7_154 0 n14 ns154 0 0.00019622343293
Gc7_155 0 n14 ns155 0 -9.30742524144e-05
Gc7_156 0 n14 ns156 0 -0.000135975398482
Gc7_157 0 n14 ns157 0 0.0005859294942
Gc7_158 0 n14 ns158 0 -0.000174103675682
Gc7_159 0 n14 ns159 0 0.000469396542748
Gc7_160 0 n14 ns160 0 -0.00207098066719
Gc7_161 0 n14 ns161 0 0.000335128832344
Gc7_162 0 n14 ns162 0 -0.000299256227639
Gc7_163 0 n14 ns163 0 0.000324821946671
Gc7_164 0 n14 ns164 0 -0.000796514568278
Gc7_165 0 n14 ns165 0 0.000684338871513
Gc7_166 0 n14 ns166 0 0.00144494995602
Gc7_167 0 n14 ns167 0 -0.00127266692837
Gc7_168 0 n14 ns168 0 -0.0002678504795
Gc7_169 0 n14 ns169 0 0.000752679345418
Gc7_170 0 n14 ns170 0 0.00356229778414
Gc7_171 0 n14 ns171 0 0.00266287581271
Gc7_172 0 n14 ns172 0 -0.00215123040086
Gc7_173 0 n14 ns173 0 0.00101799080831
Gc7_174 0 n14 ns174 0 -0.000405226762023
Gc7_175 0 n14 ns175 0 0.0014110447933
Gc7_176 0 n14 ns176 0 0.00496367795319
Gc7_177 0 n14 ns177 0 0.00968218893339
Gc7_178 0 n14 ns178 0 0.0111606973846
Gc7_179 0 n14 ns179 0 0.00156743328362
Gc7_180 0 n14 ns180 0 -0.00244737458325
Gc7_181 0 n14 ns181 0 0.00182759171567
Gc7_182 0 n14 ns182 0 -0.0120004698821
Gc7_183 0 n14 ns183 0 -0.00846870655704
Gc7_184 0 n14 ns184 0 0.011857335372
Gc7_185 0 n14 ns185 0 1.21166964815e-06
Gc7_186 0 n14 ns186 0 0.00850020421811
Gc7_187 0 n14 ns187 0 -0.00092303939743
Gc7_188 0 n14 ns188 0 -0.000142275736481
Gc7_189 0 n14 ns189 0 -3.09337039729e-05
Gc7_190 0 n14 ns190 0 -1.21788059997e-05
Gc7_191 0 n14 ns191 0 0.000426409624707
Gc7_192 0 n14 ns192 0 -5.52139536317e-05
Gc7_193 0 n14 ns193 0 -0.000384958021139
Gc7_194 0 n14 ns194 0 0.000341008197838
Gc7_195 0 n14 ns195 0 -0.000177089367648
Gc7_196 0 n14 ns196 0 0.000562304041052
Gc7_197 0 n14 ns197 0 -0.00130874933996
Gc7_198 0 n14 ns198 0 -0.000803030450326
Gc7_199 0 n14 ns199 0 -0.000321508125409
Gc7_200 0 n14 ns200 0 0.000398903178995
Gc7_201 0 n14 ns201 0 -2.63449121594e-05
Gc7_202 0 n14 ns202 0 0.000464598896124
Gc7_203 0 n14 ns203 0 0.00129596490161
Gc7_204 0 n14 ns204 0 -0.000225465482896
Gc7_205 0 n14 ns205 0 -0.000219942013288
Gc7_206 0 n14 ns206 0 0.000897121238754
Gc7_207 0 n14 ns207 0 0.00131774501103
Gc7_208 0 n14 ns208 0 0.00100645563281
Gc7_209 0 n14 ns209 0 -0.00185267175951
Gc7_210 0 n14 ns210 0 0.000208725256632
Gc7_211 0 n14 ns211 0 -0.000413636883364
Gc7_212 0 n14 ns212 0 0.00152093287526
Gc7_213 0 n14 ns213 0 0.00384455029836
Gc7_214 0 n14 ns214 0 0.00583030876273
Gc7_215 0 n14 ns215 0 0.0100407485741
Gc7_216 0 n14 ns216 0 0.00163090268655
Gc7_217 0 n14 ns217 0 -0.00302428065296
Gc7_218 0 n14 ns218 0 0.00195196162446
Gc7_219 0 n14 ns219 0 -0.00163393765964
Gc7_220 0 n14 ns220 0 -0.0113898751618
Gc7_221 0 n14 ns221 0 0.00195369995172
Gc7_222 0 n14 ns222 0 4.24087025185e-06
Gc7_223 0 n14 ns223 0 0.0103970141588
Gc7_224 0 n14 ns224 0 0.000741844796154
Gc7_225 0 n14 ns225 0 -0.00106891465459
Gc7_226 0 n14 ns226 0 2.77620846079e-06
Gc7_227 0 n14 ns227 0 6.1740700868e-06
Gc7_228 0 n14 ns228 0 9.9782006499e-05
Gc7_229 0 n14 ns229 0 2.93052175264e-05
Gc7_230 0 n14 ns230 0 -0.000410113030246
Gc7_231 0 n14 ns231 0 7.39237042993e-07
Gc7_232 0 n14 ns232 0 0.000535960312496
Gc7_233 0 n14 ns233 0 -0.000223505823124
Gc7_234 0 n14 ns234 0 0.000800057502822
Gc7_235 0 n14 ns235 0 -0.000277182503624
Gc7_236 0 n14 ns236 0 -0.000204306921815
Gc7_237 0 n14 ns237 0 0.00028102333442
Gc7_238 0 n14 ns238 0 0.000653501913605
Gc7_239 0 n14 ns239 0 -0.00149490698106
Gc7_240 0 n14 ns240 0 -0.00125593013954
Gc7_241 0 n14 ns241 0 0.000752599141812
Gc7_242 0 n14 ns242 0 -0.000142943670637
Gc7_243 0 n14 ns243 0 0.000702459454006
Gc7_244 0 n14 ns244 0 -0.00545756085394
Gc7_245 0 n14 ns245 0 -0.000233846434938
Gc7_246 0 n14 ns246 0 0.00304819988952
Gc7_247 0 n14 ns247 0 -0.000394440195401
Gc7_248 0 n14 ns248 0 -0.000234549462991
Gc7_249 0 n14 ns249 0 0.00158747793909
Gc7_250 0 n14 ns250 0 -0.00684348932632
Gc7_251 0 n14 ns251 0 -0.00788035001245
Gc7_252 0 n14 ns252 0 -0.0128876769236
Gc7_253 0 n14 ns253 0 -0.00146330649169
Gc7_254 0 n14 ns254 0 -0.00195696359962
Gc7_255 0 n14 ns255 0 0.00142694380519
Gc7_256 0 n14 ns256 0 -0.0150522613594
Gc7_257 0 n14 ns257 0 -0.00262992229316
Gc7_258 0 n14 ns258 0 0.00337212928281
Gc7_259 0 n14 ns259 0 1.00535890787e-05
Gc7_260 0 n14 ns260 0 0.0114843830833
Gc7_261 0 n14 ns261 0 -0.000501750774889
Gc7_262 0 n14 ns262 0 -0.00132653155178
Gc7_263 0 n14 ns263 0 -5.59152664542e-06
Gc7_264 0 n14 ns264 0 -6.28015906242e-06
Gc7_265 0 n14 ns265 0 0.000226583339109
Gc7_266 0 n14 ns266 0 -2.32705210968e-05
Gc7_267 0 n14 ns267 0 -0.000439356865105
Gc7_268 0 n14 ns268 0 -1.44104482693e-05
Gc7_269 0 n14 ns269 0 0.000307242783757
Gc7_270 0 n14 ns270 0 -8.66220619734e-05
Gc7_271 0 n14 ns271 0 0.000590136904339
Gc7_272 0 n14 ns272 0 -9.56270815015e-05
Gc7_273 0 n14 ns273 0 -0.000293251891728
Gc7_274 0 n14 ns274 0 0.000368991820263
Gc7_275 0 n14 ns275 0 8.74686169826e-05
Gc7_276 0 n14 ns276 0 -0.000847227184574
Gc7_277 0 n14 ns277 0 -0.001092230023
Gc7_278 0 n14 ns278 0 0.000398674300908
Gc7_279 0 n14 ns279 0 -0.000196247732983
Gc7_280 0 n14 ns280 0 0.000876795203903
Gc7_281 0 n14 ns281 0 -0.00255500326591
Gc7_282 0 n14 ns282 0 0.000537153270359
Gc7_283 0 n14 ns283 0 0.00243307502361
Gc7_284 0 n14 ns284 0 -0.00023311366631
Gc7_285 0 n14 ns285 0 -0.000280102524085
Gc7_286 0 n14 ns286 0 0.00176769511963
Gc7_287 0 n14 ns287 0 -0.00287687257172
Gc7_288 0 n14 ns288 0 -0.00198598981892
Gc7_289 0 n14 ns289 0 -0.00776556232531
Gc7_290 0 n14 ns290 0 0.000175062111214
Gc7_291 0 n14 ns291 0 -0.00262917927002
Gc7_292 0 n14 ns292 0 0.00151588576794
Gc7_293 0 n14 ns293 0 -0.018760805193
Gc7_294 0 n14 ns294 0 -0.00375332259728
Gc7_295 0 n14 ns295 0 0.00685298110249
Gc7_296 0 n14 ns296 0 5.30103495469e-06
Gd7_1 0 n14 ni1 0 0.000546119737459
Gd7_2 0 n14 ni2 0 -0.000535648881537
Gd7_3 0 n14 ni3 0 0.000563891774361
Gd7_4 0 n14 ni4 0 -0.000383522682271
Gd7_5 0 n14 ni5 0 -0.000884161597368
Gd7_6 0 n14 ni6 0 -0.00380616256527
Gd7_7 0 n14 ni7 0 -0.00253984626321
Gd7_8 0 n14 ni8 0 -0.00248151814875
Gc8_1 0 n16 ns1 0 0.000930893720336
Gc8_2 0 n16 ns2 0 0.000390272177904
Gc8_3 0 n16 ns3 0 0.000346896712812
Gc8_4 0 n16 ns4 0 1.05835887157e-05
Gc8_5 0 n16 ns5 0 1.21332860989e-05
Gc8_6 0 n16 ns6 0 1.80528916665e-05
Gc8_7 0 n16 ns7 0 -0.000211783085902
Gc8_8 0 n16 ns8 0 7.44025816358e-05
Gc8_9 0 n16 ns9 0 0.000241499089185
Gc8_10 0 n16 ns10 0 0.000305806802029
Gc8_11 0 n16 ns11 0 -0.000186410892682
Gc8_12 0 n16 ns12 0 0.00135886257832
Gc8_13 0 n16 ns13 0 -0.000512160286
Gc8_14 0 n16 ns14 0 0.000324970833894
Gc8_15 0 n16 ns15 0 -0.000372851039632
Gc8_16 0 n16 ns16 0 0.000388750962574
Gc8_17 0 n16 ns17 0 0.000799795652237
Gc8_18 0 n16 ns18 0 0.00173043508026
Gc8_19 0 n16 ns19 0 -0.000183480396525
Gc8_20 0 n16 ns20 0 -0.000172766503357
Gc8_21 0 n16 ns21 0 0.000871929273123
Gc8_22 0 n16 ns22 0 -0.00204443941884
Gc8_23 0 n16 ns23 0 -0.00315159747354
Gc8_24 0 n16 ns24 0 0.00172590811239
Gc8_25 0 n16 ns25 0 -0.000523118097111
Gc8_26 0 n16 ns26 0 0.000458699652015
Gc8_27 0 n16 ns27 0 -0.00156143590833
Gc8_28 0 n16 ns28 0 -0.00301622218186
Gc8_29 0 n16 ns29 0 -0.00019238419613
Gc8_30 0 n16 ns30 0 0.00555291000597
Gc8_31 0 n16 ns31 0 -0.000854843556866
Gc8_32 0 n16 ns32 0 -0.00269912152914
Gc8_33 0 n16 ns33 0 0.00219540696246
Gc8_34 0 n16 ns34 0 0.0023035347535
Gc8_35 0 n16 ns35 0 0.0109005214097
Gc8_36 0 n16 ns36 0 -0.00210730198768
Gc8_37 0 n16 ns37 0 -5.6575114074e-06
Gc8_38 0 n16 ns38 0 0.00160303136355
Gc8_39 0 n16 ns39 0 -8.87190023233e-05
Gc8_40 0 n16 ns40 0 0.000446673538466
Gc8_41 0 n16 ns41 0 -5.93886462342e-06
Gc8_42 0 n16 ns42 0 1.17695464915e-05
Gc8_43 0 n16 ns43 0 0.000268865143246
Gc8_44 0 n16 ns44 0 -0.000189108382669
Gc8_45 0 n16 ns45 0 -0.000511741880121
Gc8_46 0 n16 ns46 0 0.000301172814833
Gc8_47 0 n16 ns47 0 -1.21231104893e-05
Gc8_48 0 n16 ns48 0 -1.26900850107e-05
Gc8_49 0 n16 ns49 0 0.00136663339275
Gc8_50 0 n16 ns50 0 -0.000158071986288
Gc8_51 0 n16 ns51 0 0.000395288143854
Gc8_52 0 n16 ns52 0 -0.00044728881575
Gc8_53 0 n16 ns53 0 0.000949426521242
Gc8_54 0 n16 ns54 0 0.000806267460323
Gc8_55 0 n16 ns55 0 0.00143593245798
Gc8_56 0 n16 ns56 0 0.000424966837822
Gc8_57 0 n16 ns57 0 -0.000188100667626
Gc8_58 0 n16 ns58 0 0.00103719865419
Gc8_59 0 n16 ns59 0 0.00106781725385
Gc8_60 0 n16 ns60 0 -0.0032956184147
Gc8_61 0 n16 ns61 0 0.00106161983963
Gc8_62 0 n16 ns62 0 -0.000322928448765
Gc8_63 0 n16 ns63 0 0.000516438762053
Gc8_64 0 n16 ns64 0 -0.0018468414164
Gc8_65 0 n16 ns65 0 -0.00157129099471
Gc8_66 0 n16 ns66 0 -0.00704567125533
Gc8_67 0 n16 ns67 0 0.0045024354981
Gc8_68 0 n16 ns68 0 -0.00322084246982
Gc8_69 0 n16 ns69 0 -0.00327010796371
Gc8_70 0 n16 ns70 0 0.00253284166539
Gc8_71 0 n16 ns71 0 0.0016444430923
Gc8_72 0 n16 ns72 0 0.0128961982804
Gc8_73 0 n16 ns73 0 -0.00032543576877
Gc8_74 0 n16 ns74 0 -6.31234022275e-06
Gc8_75 0 n16 ns75 0 0.0030385568282
Gc8_76 0 n16 ns76 0 -0.000983268825471
Gc8_77 0 n16 ns77 0 0.000684672432746
Gc8_78 0 n16 ns78 0 -2.12746306183e-05
Gc8_79 0 n16 ns79 0 -2.36731993992e-06
Gc8_80 0 n16 ns80 0 0.00043313785348
Gc8_81 0 n16 ns81 0 -0.00014133265241
Gc8_82 0 n16 ns82 0 -0.000643567406704
Gc8_83 0 n16 ns83 0 0.000754568520243
Gc8_84 0 n16 ns84 0 -0.000685288264663
Gc8_85 0 n16 ns85 0 0.00030891797195
Gc8_86 0 n16 ns86 0 0.00135627779829
Gc8_87 0 n16 ns87 0 0.000353934563758
Gc8_88 0 n16 ns88 0 0.00026568294822
Gc8_89 0 n16 ns89 0 -0.000379766799295
Gc8_90 0 n16 ns90 0 0.000439835610556
Gc8_91 0 n16 ns91 0 -0.000995177211752
Gc8_92 0 n16 ns92 0 -0.000733175090967
Gc8_93 0 n16 ns93 0 0.000943955605679
Gc8_94 0 n16 ns94 0 -0.000150302823681
Gc8_95 0 n16 ns95 0 0.000922028215635
Gc8_96 0 n16 ns96 0 0.0113027189165
Gc8_97 0 n16 ns97 0 -0.00591883396504
Gc8_98 0 n16 ns98 0 -0.00186547178094
Gc8_99 0 n16 ns99 0 -0.000100667009643
Gc8_100 0 n16 ns100 0 0.000367864537348
Gc8_101 0 n16 ns101 0 -0.00170214516726
Gc8_102 0 n16 ns102 0 -0.00256158814838
Gc8_103 0 n16 ns103 0 -0.0301002309849
Gc8_104 0 n16 ns104 0 -0.00433576367038
Gc8_105 0 n16 ns105 0 -0.0108191338543
Gc8_106 0 n16 ns106 0 -0.00311497805359
Gc8_107 0 n16 ns107 0 0.00223833690252
Gc8_108 0 n16 ns108 0 -0.0150198138066
Gc8_109 0 n16 ns109 0 0.0127522891874
Gc8_110 0 n16 ns110 0 0.0181925103639
Gc8_111 0 n16 ns111 0 -1.23212397547e-05
Gc8_112 0 n16 ns112 0 -0.000337744486198
Gc8_113 0 n16 ns113 0 -6.61515243022e-05
Gc8_114 0 n16 ns114 0 -0.0010492473369
Gc8_115 0 n16 ns115 0 1.54325056937e-05
Gc8_116 0 n16 ns116 0 -1.43124514809e-06
Gc8_117 0 n16 ns117 0 3.00868695046e-05
Gc8_118 0 n16 ns118 0 0.000168924289619
Gc8_119 0 n16 ns119 0 -0.00016160487068
Gc8_120 0 n16 ns120 0 -0.000247429000244
Gc8_121 0 n16 ns121 0 0.000318180369639
Gc8_122 0 n16 ns122 0 -0.00017562127118
Gc8_123 0 n16 ns123 0 -0.00237630507965
Gc8_124 0 n16 ns124 0 0.000214948688347
Gc8_125 0 n16 ns125 0 0.000378777455809
Gc8_126 0 n16 ns126 0 -0.000478760048988
Gc8_127 0 n16 ns127 0 -0.000625536663358
Gc8_128 0 n16 ns128 0 0.00120197470437
Gc8_129 0 n16 ns129 0 -0.00171385719029
Gc8_130 0 n16 ns130 0 0.000217393798682
Gc8_131 0 n16 ns131 0 -0.000314418047298
Gc8_132 0 n16 ns132 0 0.00106105059833
Gc8_133 0 n16 ns133 0 -0.00858039460272
Gc8_134 0 n16 ns134 0 0.00822723057112
Gc8_135 0 n16 ns135 0 -0.00185432635789
Gc8_136 0 n16 ns136 0 0.000279834640773
Gc8_137 0 n16 ns137 0 0.000427692592964
Gc8_138 0 n16 ns138 0 -0.00198435376606
Gc8_139 0 n16 ns139 0 0.00881730483623
Gc8_140 0 n16 ns140 0 0.0289700150227
Gc8_141 0 n16 ns141 0 -0.00491415025558
Gc8_142 0 n16 ns142 0 0.0100368763518
Gc8_143 0 n16 ns143 0 -0.00288762687028
Gc8_144 0 n16 ns144 0 0.00127809525197
Gc8_145 0 n16 ns145 0 0.0606085822886
Gc8_146 0 n16 ns146 0 -0.00370655029884
Gc8_147 0 n16 ns147 0 -0.0392998140915
Gc8_148 0 n16 ns148 0 1.742112078e-05
Gc8_149 0 n16 ns149 0 0.00852676888861
Gc8_150 0 n16 ns150 0 -0.000928228056204
Gc8_151 0 n16 ns151 0 -0.000139506479497
Gc8_152 0 n16 ns152 0 -3.1120103486e-05
Gc8_153 0 n16 ns153 0 -1.21075987798e-05
Gc8_154 0 n16 ns154 0 0.000426981148591
Gc8_155 0 n16 ns155 0 -5.50141332484e-05
Gc8_156 0 n16 ns156 0 -0.000384925585593
Gc8_157 0 n16 ns157 0 0.000345685512429
Gc8_158 0 n16 ns158 0 -0.000176254626931
Gc8_159 0 n16 ns159 0 0.000567016708109
Gc8_160 0 n16 ns160 0 -0.00132094625523
Gc8_161 0 n16 ns161 0 -0.000801205278281
Gc8_162 0 n16 ns162 0 -0.000321384898202
Gc8_163 0 n16 ns163 0 0.000400841302388
Gc8_164 0 n16 ns164 0 -2.9550198043e-05
Gc8_165 0 n16 ns165 0 0.000466137186062
Gc8_166 0 n16 ns166 0 0.00129895998816
Gc8_167 0 n16 ns167 0 -0.000228823884327
Gc8_168 0 n16 ns168 0 -0.00021951797882
Gc8_169 0 n16 ns169 0 0.000898798346262
Gc8_170 0 n16 ns170 0 0.00131931987024
Gc8_171 0 n16 ns171 0 0.00100473027475
Gc8_172 0 n16 ns172 0 -0.00184677050125
Gc8_173 0 n16 ns173 0 0.000222034422596
Gc8_174 0 n16 ns174 0 -0.000409236202205
Gc8_175 0 n16 ns175 0 0.00152844671747
Gc8_176 0 n16 ns176 0 0.00384986278146
Gc8_177 0 n16 ns177 0 0.00584019980302
Gc8_178 0 n16 ns178 0 0.0100307069765
Gc8_179 0 n16 ns179 0 0.00161681585832
Gc8_180 0 n16 ns180 0 -0.00302057750664
Gc8_181 0 n16 ns181 0 0.00196017500986
Gc8_182 0 n16 ns182 0 -0.00174893369741
Gc8_183 0 n16 ns183 0 -0.0113616010269
Gc8_184 0 n16 ns184 0 0.00204931712026
Gc8_185 0 n16 ns185 0 4.32728344905e-06
Gc8_186 0 n16 ns186 0 0.00763103524367
Gc8_187 0 n16 ns187 0 -0.000573185939106
Gc8_188 0 n16 ns188 0 -0.000855495854126
Gc8_189 0 n16 ns189 0 -9.95962597473e-06
Gc8_190 0 n16 ns190 0 3.806127393e-06
Gc8_191 0 n16 ns191 0 0.000331062298821
Gc8_192 0 n16 ns192 0 -7.03325563636e-05
Gc8_193 0 n16 ns193 0 -0.000325846706908
Gc8_194 0 n16 ns194 0 0.000417831692434
Gc8_195 0 n16 ns195 0 2.94155151997e-05
Gc8_196 0 n16 ns196 0 0.000270419711241
Gc8_197 0 n16 ns197 0 -0.00142356905215
Gc8_198 0 n16 ns198 0 2.70182194954e-05
Gc8_199 0 n16 ns199 0 -0.000381569897987
Gc8_200 0 n16 ns200 0 0.000443826036255
Gc8_201 0 n16 ns201 0 -0.00062874558507
Gc8_202 0 n16 ns202 0 -0.000123278964322
Gc8_203 0 n16 ns203 0 0.000703627726472
Gc8_204 0 n16 ns204 0 -0.000631581147129
Gc8_205 0 n16 ns205 0 -0.000315962471246
Gc8_206 0 n16 ns206 0 0.00100921081011
Gc8_207 0 n16 ns207 0 0.000994903910945
Gc8_208 0 n16 ns208 0 0.00234481516784
Gc8_209 0 n16 ns209 0 -0.000659995519268
Gc8_210 0 n16 ns210 0 0.000593730789499
Gc8_211 0 n16 ns211 0 -0.000538812216078
Gc8_212 0 n16 ns212 0 0.00193931290453
Gc8_213 0 n16 ns213 0 0.00274526276172
Gc8_214 0 n16 ns214 0 0.0054526686525
Gc8_215 0 n16 ns215 0 0.00537521533104
Gc8_216 0 n16 ns216 0 0.000465410040155
Gc8_217 0 n16 ns217 0 -0.00332333858418
Gc8_218 0 n16 ns218 0 0.00226922546488
Gc8_219 0 n16 ns219 0 -0.0134095472782
Gc8_220 0 n16 ns220 0 -0.00888982602847
Gc8_221 0 n16 ns221 0 0.00826425513552
Gc8_222 0 n16 ns222 0 3.93530957485e-06
Gc8_223 0 n16 ns223 0 0.0114843830907
Gc8_224 0 n16 ns224 0 -0.000501750775001
Gc8_225 0 n16 ns225 0 -0.00132653155049
Gc8_226 0 n16 ns226 0 -5.59152675885e-06
Gc8_227 0 n16 ns227 0 -6.28015903689e-06
Gc8_228 0 n16 ns228 0 0.000226583339841
Gc8_229 0 n16 ns229 0 -2.32705207484e-05
Gc8_230 0 n16 ns230 0 -0.00043935686453
Gc8_231 0 n16 ns231 0 -1.44104476369e-05
Gc8_232 0 n16 ns232 0 0.000307242784768
Gc8_233 0 n16 ns233 0 -8.66220616273e-05
Gc8_234 0 n16 ns234 0 0.000590136901866
Gc8_235 0 n16 ns235 0 -9.56270798204e-05
Gc8_236 0 n16 ns236 0 -0.000293251891971
Gc8_237 0 n16 ns237 0 0.000368991819941
Gc8_238 0 n16 ns238 0 8.74686130754e-05
Gc8_239 0 n16 ns239 0 -0.000847227184211
Gc8_240 0 n16 ns240 0 -0.00109223002539
Gc8_241 0 n16 ns241 0 0.000398674301359
Gc8_242 0 n16 ns242 0 -0.000196247733196
Gc8_243 0 n16 ns243 0 0.000876795204022
Gc8_244 0 n16 ns244 0 -0.00255500324837
Gc8_245 0 n16 ns245 0 0.000537153267097
Gc8_246 0 n16 ns246 0 0.00243307501956
Gc8_247 0 n16 ns247 0 -0.000233113674029
Gc8_248 0 n16 ns248 0 -0.000280102523484
Gc8_249 0 n16 ns249 0 0.00176769511676
Gc8_250 0 n16 ns250 0 -0.00287687254749
Gc8_251 0 n16 ns251 0 -0.00198598987975
Gc8_252 0 n16 ns252 0 -0.00776556233175
Gc8_253 0 n16 ns253 0 0.000175062069051
Gc8_254 0 n16 ns254 0 -0.00262917926716
Gc8_255 0 n16 ns255 0 0.00151588577316
Gc8_256 0 n16 ns256 0 -0.0187608050656
Gc8_257 0 n16 ns257 0 -0.00375332261977
Gc8_258 0 n16 ns258 0 0.00685298098967
Gc8_259 0 n16 ns259 0 5.30103462349e-06
Gc8_260 0 n16 ns260 0 0.00620268758069
Gc8_261 0 n16 ns261 0 0.000553931235234
Gc8_262 0 n16 ns262 0 -0.00124194937361
Gc8_263 0 n16 ns263 0 1.64754923048e-05
Gc8_264 0 n16 ns264 0 5.1534011752e-06
Gc8_265 0 n16 ns265 0 9.44219081872e-05
Gc8_266 0 n16 ns266 0 1.8410436586e-05
Gc8_267 0 n16 ns267 0 -0.000315639648566
Gc8_268 0 n16 ns268 0 0.000122106841436
Gc8_269 0 n16 ns269 0 0.000325614747439
Gc8_270 0 n16 ns270 0 -0.000163975921284
Gc8_271 0 n16 ns271 0 0.000152866418697
Gc8_272 0 n16 ns272 0 0.000504591737053
Gc8_273 0 n16 ns273 0 -0.000383719156309
Gc8_274 0 n16 ns274 0 0.000441990732617
Gc8_275 0 n16 ns275 0 -0.00015419116068
Gc8_276 0 n16 ns276 0 -0.000935520068277
Gc8_277 0 n16 ns277 0 -0.000803008115418
Gc8_278 0 n16 ns278 0 7.84011759253e-05
Gc8_279 0 n16 ns279 0 -0.000260646049704
Gc8_280 0 n16 ns280 0 0.00104268062906
Gc8_281 0 n16 ns281 0 -0.00260597318282
Gc8_282 0 n16 ns282 0 0.00106692660862
Gc8_283 0 n16 ns283 0 0.00169458741006
Gc8_284 0 n16 ns284 0 -9.93537696486e-05
Gc8_285 0 n16 ns285 0 -0.000396440940555
Gc8_286 0 n16 ns286 0 0.00196057382845
Gc8_287 0 n16 ns287 0 -0.0034193241404
Gc8_288 0 n16 ns288 0 -0.00340929651061
Gc8_289 0 n16 ns289 0 -0.00588702510098
Gc8_290 0 n16 ns290 0 -0.000839610978743
Gc8_291 0 n16 ns291 0 -0.00305122021844
Gc8_292 0 n16 ns292 0 0.00197433777653
Gc8_293 0 n16 ns293 0 -0.0144920119661
Gc8_294 0 n16 ns294 0 -0.00753078298837
Gc8_295 0 n16 ns295 0 0.00473555232561
Gc8_296 0 n16 ns296 0 1.10212926114e-05
Gd8_1 0 n16 ni1 0 -0.00054918314948
Gd8_2 0 n16 ni2 0 -0.000366569199659
Gd8_3 0 n16 ni3 0 -0.000387208136655
Gd8_4 0 n16 ni4 0 4.38357026971e-06
Gd8_5 0 n16 ni5 0 -0.00381869963683
Gd8_6 0 n16 ni6 0 -0.0023955916148
Gd8_7 0 n16 ni7 0 -0.00248151815281
Gd8_8 0 n16 ni8 0 -0.000157856163283
.ends m4lines_HFSS_fws
